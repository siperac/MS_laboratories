
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file_NBIT64_NREG32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file_NBIT64_NREG32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file_NBIT64_NREG32.all;

entity register_file_NBIT64_NREG32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_NBIT64_NREG32;

architecture SYN_A of register_file_NBIT64_NREG32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal OUT1_63_port, OUT1_62_port, OUT1_61_port, OUT1_60_port, OUT1_59_port,
      OUT1_58_port, OUT1_57_port, OUT1_56_port, OUT1_55_port, OUT1_54_port, 
      OUT1_53_port, OUT1_52_port, OUT1_51_port, OUT1_50_port, OUT1_49_port, 
      OUT1_48_port, OUT1_47_port, OUT1_46_port, OUT1_45_port, OUT1_44_port, 
      OUT1_43_port, OUT1_42_port, OUT1_41_port, OUT1_40_port, OUT1_39_port, 
      OUT1_38_port, OUT1_37_port, OUT1_36_port, OUT1_35_port, OUT1_34_port, 
      OUT1_33_port, OUT1_32_port, OUT1_31_port, OUT1_30_port, OUT1_29_port, 
      OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, 
      OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, 
      OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, 
      OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, 
      OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, 
      OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port, OUT2_63_port, 
      OUT2_62_port, OUT2_61_port, OUT2_60_port, OUT2_59_port, OUT2_58_port, 
      OUT2_57_port, OUT2_56_port, OUT2_55_port, OUT2_54_port, OUT2_53_port, 
      OUT2_52_port, OUT2_51_port, OUT2_50_port, OUT2_49_port, OUT2_48_port, 
      OUT2_47_port, OUT2_46_port, OUT2_45_port, OUT2_44_port, OUT2_43_port, 
      OUT2_42_port, OUT2_41_port, OUT2_40_port, OUT2_39_port, OUT2_38_port, 
      OUT2_37_port, OUT2_36_port, OUT2_35_port, OUT2_34_port, OUT2_33_port, 
      OUT2_32_port, OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, 
      OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, 
      OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, 
      OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, 
      OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, 
      OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port, n5311, n5312, n5313, n5314, n5315,
      n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, 
      n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, 
      n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, 
      n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, 
      n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, 
      n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, 
      n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, 
      n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, 
      n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, 
      n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, 
      n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, 
      n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, 
      n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, 
      n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, 
      n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, 
      n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, 
      n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, 
      n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, 
      n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, 
      n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, 
      n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, 
      n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, 
      n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, 
      n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, 
      n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, 
      n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, 
      n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, 
      n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, 
      n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, 
      n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, 
      n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, 
      n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, 
      n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, 
      n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, 
      n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, 
      n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, 
      n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, 
      n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, 
      n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, 
      n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, 
      n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, 
      n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, 
      n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, 
      n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, 
      n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, 
      n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, 
      n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, 
      n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, 
      n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, 
      n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, 
      n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, 
      n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, 
      n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, 
      n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, 
      n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, 
      n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, 
      n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, 
      n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, 
      n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, 
      n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, 
      n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, 
      n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, 
      n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, 
      n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, 
      n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, 
      n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, 
      n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, 
      n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, 
      n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, 
      n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, 
      n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, 
      n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, 
      n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, 
      n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, 
      n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, 
      n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, 
      n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, 
      n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, 
      n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, 
      n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, 
      n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, 
      n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, 
      n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, 
      n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, 
      n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, 
      n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, 
      n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, 
      n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, 
      n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, 
      n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, 
      n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, 
      n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, 
      n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, 
      n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, 
      n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, 
      n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, 
      n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, 
      n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, 
      n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, 
      n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, 
      n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, 
      n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, 
      n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, 
      n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, 
      n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, 
      n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, 
      n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, 
      n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, 
      n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, 
      n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, 
      n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, 
      n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, 
      n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, 
      n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, 
      n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, 
      n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, 
      n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, 
      n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, 
      n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, 
      n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, 
      n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, 
      n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, 
      n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, 
      n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, 
      n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, 
      n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, 
      n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, 
      n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, 
      n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, 
      n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, 
      n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, 
      n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, 
      n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, 
      n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, 
      n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, 
      n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, 
      n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, 
      n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, 
      n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, 
      n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, 
      n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, 
      n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, 
      n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, 
      n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, 
      n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, 
      n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, 
      n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, 
      n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, 
      n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, 
      n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, 
      n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, 
      n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, 
      n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, 
      n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, 
      n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, 
      n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, 
      n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, 
      n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, 
      n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, 
      n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, 
      n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, 
      n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, 
      n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, 
      n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, 
      n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, 
      n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, 
      n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, 
      n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, 
      n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, 
      n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, 
      n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, 
      n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, 
      n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, 
      n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, 
      n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, 
      n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, 
      n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, 
      n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, 
      n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, 
      n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, 
      n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, 
      n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, 
      n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, 
      n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, 
      n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, 
      n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, 
      n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, 
      n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, 
      n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, 
      n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, 
      n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, 
      n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, 
      n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, 
      n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, 
      n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, 
      n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, 
      n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, 
      n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, 
      n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, 
      n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, 
      n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, 
      n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, 
      n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, 
      n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, 
      n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, 
      n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, 
      n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, 
      n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, 
      n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, 
      n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, 
      n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, 
      n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, 
      n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, 
      n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, 
      n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, 
      n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, 
      n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, 
      n7486, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, 
      n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, 
      n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, 
      n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, 
      n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, 
      n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, 
      n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, 
      n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, 
      n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, 
      n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, 
      n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, 
      n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, 
      n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9223, 
      n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, 
      n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, 
      n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, 
      n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, 
      n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, 
      n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, 
      n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, 
      n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, 
      n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, 
      n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, 
      n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, 
      n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, 
      n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9415, n9416, n9417, 
      n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, 
      n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, 
      n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, 
      n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, 
      n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, 
      n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, 
      n9478, n17148, n17149, n17156, n17157, n17161, n17163, n17169, n17170, 
      n17177, n17178, n17182, n17184, n17190, n17191, n17198, n17199, n17203, 
      n17205, n17211, n17212, n17219, n17220, n17224, n17226, n17232, n17233, 
      n17240, n17241, n17245, n17247, n17253, n17254, n17261, n17262, n17266, 
      n17268, n17274, n17275, n17282, n17283, n17287, n17289, n17295, n17296, 
      n17303, n17304, n17308, n17310, n17316, n17317, n17324, n17325, n17329, 
      n17331, n17337, n17338, n17345, n17346, n17350, n17352, n17358, n17359, 
      n17366, n17367, n17371, n17373, n17379, n17380, n17387, n17388, n17392, 
      n17394, n17400, n17401, n17408, n17409, n17413, n17415, n17421, n17422, 
      n17429, n17430, n17434, n17436, n17442, n17443, n17450, n17451, n17455, 
      n17457, n17463, n17464, n17471, n17472, n17476, n17478, n17484, n17485, 
      n17492, n17493, n17497, n17499, n17505, n17506, n17513, n17514, n17518, 
      n17520, n17526, n17527, n17534, n17535, n17539, n17541, n17547, n17548, 
      n17555, n17556, n17560, n17562, n17568, n17569, n17576, n17577, n17581, 
      n17583, n17589, n17590, n17597, n17598, n17602, n17604, n17610, n17611, 
      n17618, n17619, n17623, n17625, n17631, n17632, n17639, n17640, n17644, 
      n17646, n17652, n17653, n17660, n17661, n17665, n17667, n17673, n17674, 
      n17681, n17682, n17686, n17688, n17694, n17695, n17702, n17703, n17707, 
      n17709, n17715, n17716, n17723, n17724, n17728, n17730, n17736, n17737, 
      n17744, n17745, n17749, n17751, n17757, n17758, n17765, n17766, n17770, 
      n17772, n17778, n17779, n17786, n17787, n17791, n17793, n17799, n17800, 
      n17807, n17808, n17812, n17814, n17820, n17821, n17828, n17829, n17833, 
      n17835, n17841, n17842, n17849, n17850, n17854, n17856, n17862, n17863, 
      n17870, n17871, n17875, n17877, n17883, n17884, n17891, n17892, n17896, 
      n17898, n17904, n17905, n17912, n17913, n17917, n17919, n17925, n17926, 
      n17933, n17934, n17938, n17940, n17946, n17947, n17954, n17955, n17959, 
      n17961, n17967, n17968, n17975, n17976, n17980, n17982, n17988, n17989, 
      n17996, n17997, n18001, n18003, n18009, n18010, n18017, n18018, n18022, 
      n18024, n18030, n18031, n18038, n18039, n18043, n18045, n18051, n18052, 
      n18059, n18060, n18064, n18066, n18072, n18073, n18080, n18081, n18085, 
      n18087, n18093, n18094, n18101, n18102, n18106, n18108, n18114, n18115, 
      n18122, n18123, n18127, n18129, n18135, n18136, n18143, n18144, n18148, 
      n18150, n18156, n18157, n18164, n18165, n18169, n18171, n18177, n18178, 
      n18185, n18186, n18190, n18192, n18198, n18199, n18206, n18207, n18211, 
      n18213, n18219, n18220, n18227, n18228, n18232, n18234, n18240, n18241, 
      n18248, n18249, n18253, n18255, n18261, n18262, n18269, n18270, n18274, 
      n18276, n18282, n18283, n18290, n18291, n18295, n18297, n18303, n18304, 
      n18311, n18312, n18316, n18318, n18324, n18325, n18332, n18333, n18337, 
      n18339, n18345, n18346, n18353, n18354, n18358, n18360, n18366, n18367, 
      n18374, n18375, n18379, n18381, n18387, n18388, n18395, n18396, n18400, 
      n18402, n18408, n18409, n18416, n18417, n18421, n18423, n18429, n18430, 
      n18437, n18438, n18442, n18444, n18450, n18451, n18458, n18459, n18463, 
      n18465, n18471, n18472, n18479, n18480, n18484, n18486, n19478, n19479, 
      n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, 
      n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, 
      n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, 
      n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, 
      n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, 
      n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, 
      n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, 
      n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, 
      n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, 
      n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, 
      n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, 
      n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, 
      n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, 
      n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, 
      n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, 
      n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, 
      n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, 
      n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, 
      n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, 
      n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, 
      n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, 
      n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, 
      n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, 
      n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, 
      n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, 
      n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, 
      n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, 
      n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, 
      n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, 
      n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, 
      n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, 
      n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, 
      n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, 
      n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, 
      n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, 
      n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, 
      n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, 
      n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, 
      n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, 
      n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, 
      n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, 
      n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, 
      n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, 
      n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, 
      n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, 
      n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, 
      n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, 
      n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, 
      n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, 
      n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, 
      n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, 
      n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, 
      n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, 
      n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, 
      n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, 
      n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, 
      n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, 
      n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, 
      n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, 
      n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, 
      n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, 
      n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, 
      n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, 
      n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, 
      n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, 
      n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, 
      n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, 
      n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, 
      n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, 
      n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, 
      n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, 
      n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, 
      n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, 
      n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, 
      n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, 
      n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, 
      n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, 
      n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, 
      n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, 
      n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, 
      n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, 
      n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, 
      n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, 
      n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, 
      n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, 
      n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, 
      n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, 
      n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, 
      n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, 
      n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, 
      n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, 
      n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, 
      n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, 
      n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, 
      n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, 
      n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, 
      n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, 
      n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, 
      n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, 
      n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, 
      n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, 
      n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, 
      n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, 
      n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, 
      n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, 
      n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, 
      n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, 
      n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, 
      n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, 
      n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, 
      n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, 
      n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, 
      n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, 
      n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, 
      n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, 
      n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, 
      n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, 
      n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, 
      n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, 
      n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, 
      n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, 
      n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, 
      n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, 
      n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, 
      n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, 
      n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, 
      n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, 
      n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, 
      n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, 
      n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, 
      n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, 
      n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, 
      n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, 
      n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, 
      n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, 
      n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, 
      n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, 
      n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, 
      n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, 
      n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, 
      n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, 
      n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, 
      n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, 
      n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, 
      n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, 
      n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, 
      n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, 
      n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, 
      n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, 
      n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, 
      n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, 
      n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, 
      n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, 
      n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, 
      n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, 
      n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, 
      n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, 
      n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, 
      n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, 
      n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, 
      n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, 
      n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, 
      n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, 
      n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, 
      n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, 
      n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, 
      n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, 
      n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, 
      n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, 
      n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, 
      n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, 
      n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, 
      n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, 
      n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, 
      n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, 
      n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, 
      n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, 
      n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, 
      n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, 
      n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, 
      n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, 
      n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, 
      n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, 
      n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, 
      n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, 
      n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, 
      n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, 
      n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, 
      n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, 
      n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, 
      n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, 
      n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, 
      n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, 
      n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, 
      n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, 
      n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, 
      n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, 
      n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, 
      n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, 
      n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, 
      n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, 
      n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, 
      n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, 
      n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, 
      n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, 
      n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, 
      n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, 
      n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, 
      n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, 
      n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, 
      n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, 
      n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, 
      n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, 
      n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, 
      n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, 
      n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, 
      n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, 
      n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, 
      n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, 
      n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, 
      n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, 
      n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, 
      n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, 
      n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, 
      n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, 
      n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, 
      n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, 
      n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, 
      n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, 
      n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, 
      n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, 
      n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, 
      n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, 
      n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, 
      n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, 
      n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, 
      n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, 
      n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, 
      n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, 
      n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, 
      n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, 
      n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, 
      n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, 
      n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, 
      n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, 
      n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, 
      n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, 
      n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, 
      n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, 
      n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, 
      n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, 
      n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, 
      n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, 
      n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, 
      n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, 
      n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, 
      n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, 
      n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, 
      n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, 
      n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, 
      n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, 
      n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, 
      n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, 
      n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, 
      n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, 
      n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, 
      n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, 
      n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, 
      n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, 
      n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, 
      n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, 
      n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, 
      n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, 
      n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, 
      n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, 
      n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, 
      n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, 
      n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, 
      n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, 
      n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, 
      n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, 
      n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, 
      n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, 
      n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, 
      n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, 
      n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, 
      n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, 
      n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, 
      n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, 
      n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, 
      n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, 
      n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, 
      n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, 
      n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, 
      n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, 
      n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, 
      n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, 
      n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, 
      n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, 
      n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, 
      n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, 
      n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, 
      n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, 
      n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, 
      n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, 
      n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, 
      n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, 
      n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, 
      n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, 
      n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, 
      n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, 
      n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, 
      n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, 
      n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, 
      n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, 
      n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, 
      n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, 
      n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, 
      n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, 
      n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, 
      n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, 
      n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, 
      n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, 
      n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, 
      n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, 
      n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, 
      n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, 
      n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, 
      n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, 
      n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, 
      n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, 
      n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, 
      n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, 
      n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, 
      n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, 
      n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, 
      n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, 
      n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, 
      n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, 
      n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, 
      n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, 
      n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, 
      n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, 
      n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, 
      n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, 
      n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, 
      n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, 
      n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, 
      n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, 
      n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, 
      n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, 
      n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, 
      n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, 
      n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, 
      n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, 
      n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, 
      n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, 
      n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, 
      n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, 
      n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, 
      n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, 
      n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, 
      n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, 
      n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, 
      n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, 
      n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, 
      n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, 
      n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, 
      n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, 
      n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, 
      n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, 
      n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, 
      n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, 
      n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, 
      n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, 
      n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, 
      n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, 
      n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, 
      n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, 
      n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, 
      n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, 
      n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, 
      n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, 
      n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, 
      n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, 
      n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, 
      n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, 
      n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, 
      n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, 
      n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, 
      n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, 
      n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, 
      n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, 
      n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, 
      n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, 
      n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, 
      n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, 
      n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, 
      n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, 
      n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, 
      n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, 
      n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, 
      n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, 
      n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, 
      n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, 
      n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, 
      n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, 
      n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, 
      n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, 
      n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, 
      n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, 
      n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, 
      n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, 
      n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, 
      n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, 
      n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, 
      n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, 
      n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, 
      n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, 
      n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, 
      n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, 
      n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, 
      n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, 
      n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, 
      n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, 
      n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, 
      n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, 
      n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, 
      n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, 
      n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, 
      n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, 
      n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, 
      n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, 
      n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, 
      n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, 
      n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, 
      n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, 
      n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, 
      n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, 
      n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, 
      n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, 
      n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, 
      n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, 
      n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, 
      n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, 
      n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, 
      n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, 
      n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, 
      n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, 
      n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, 
      n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, 
      n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, 
      n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, 
      n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, 
      n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, 
      n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, 
      n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, 
      n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, 
      n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, 
      n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, 
      n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, 
      n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, 
      n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, 
      n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, 
      n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, 
      n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, 
      n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, 
      n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, 
      n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700, 
      n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, 
      n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, 
      n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, 
      n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, 
      n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, 
      n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754, 
      n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, 
      n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, 
      n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781, 
      n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, 
      n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, 
      n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, 
      n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, 
      n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, 
      n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, 
      n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, 
      n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, 
      n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, 
      n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, 
      n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, 
      n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, 
      n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, 
      n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, 
      n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, 
      n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, 
      n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, 
      n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, 
      n23944, n23945, n23946, n23947, n23948, n23949, n23954, n23955, n23956, 
      n23957, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025, 
      n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034, 
      n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043, 
      n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052, 
      n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061, 
      n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070, 
      n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24079, n24081, 
      n24083, n24085, n24087, n24089, n24091, n24093, n24095, n24097, n24099, 
      n24101, n24103, n24105, n24107, n24109, n24111, n24113, n24115, n24117, 
      n24119, n24121, n24123, n24125, n24127, n24129, n24131, n24133, n24135, 
      n24137, n24139, n24141, n24143, n24145, n24147, n24149, n24151, n24153, 
      n24155, n24157, n24159, n24161, n24163, n24165, n24167, n24169, n24171, 
      n24173, n24175, n24177, n24179, n24181, n24183, n24185, n24187, n24189, 
      n24191, n24193, n24195, n24197, n24199, n24201, n24203, n24205, n24206, 
      n24208, n24210, n24212, n24214, n24216, n24218, n24220, n24222, n24224, 
      n24226, n24228, n24230, n24232, n24234, n24236, n24238, n24240, n24242, 
      n24244, n24246, n24248, n24250, n24252, n24254, n24256, n24258, n24260, 
      n24262, n24264, n24266, n24268, n24270, n24272, n24274, n24276, n24278, 
      n24280, n24282, n24284, n24286, n24288, n24290, n24292, n24294, n24296, 
      n24298, n24300, n24302, n24305, n24308, n24311, n24314, n24316, n24318, 
      n24320, n24322, n24324, n24326, n24328, n24330, n24332, n24334, n24336, 
      n24339, n24341, n24343, n24345, n24347, n24349, n24351, n24353, n24355, 
      n24357, n24359, n24361, n24363, n24365, n24367, n24369, n24371, n24373, 
      n24375, n24377, n24379, n24381, n24383, n24385, n24387, n24389, n24391, 
      n24393, n24395, n24397, n24399, n24401, n24403, n24405, n24407, n24409, 
      n24411, n24413, n24415, n24417, n24419, n24421, n24423, n24425, n24427, 
      n24429, n24431, n24433, n24435, n24437, n24439, n24441, n24443, n24445, 
      n24447, n24449, n24451, n24453, n24455, n24457, n24459, n24461, n24463, 
      n24465, n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481, 
      n24607, n24609, n24611, n24613, n24614, n24615, n24616, n24617, n24618, 
      n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, 
      n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, 
      n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, 
      n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, 
      n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, 
      n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, 
      n24673, n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, 
      n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, 
      n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, 
      n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, 
      n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, 
      n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, 
      n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, 
      n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, 
      n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, 
      n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, 
      n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, 
      n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, 
      n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, 
      n24910, n24911, n24912, n24913, n24974, n24975, n24976, n24977, n24978, 
      n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, 
      n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, 
      n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005, 
      n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, 
      n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, 
      n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, 
      n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, 
      n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, 
      n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, 
      n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, 
      n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, 
      n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, 
      n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, 
      n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, 
      n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, 
      n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, 
      n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, 
      n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, 
      n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, 
      n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, 
      n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, 
      n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, 
      n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, 
      n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, 
      n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, 
      n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, 
      n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, 
      n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, 
      n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, 
      n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, 
      n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, 
      n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, 
      n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, 
      n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, 
      n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, 
      n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, 
      n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, 
      n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, 
      n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, 
      n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, 
      n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, 
      n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, 
      n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, 
      n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, 
      n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, 
      n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, 
      n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, 
      n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, 
      n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, 
      n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, 
      n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, 
      n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, 
      n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, 
      n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, 
      n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, 
      n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, 
      n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, 
      n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, 
      n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, 
      n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, 
      n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, 
      n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, 
      n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, 
      n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, 
      n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, 
      n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, 
      n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, 
      n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, 
      n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, 
      n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, 
      n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, 
      n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, 
      n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, 
      n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, 
      n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, 
      n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, 
      n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, 
      n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680, 
      n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689, 
      n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698, 
      n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707, 
      n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, 
      n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725, 
      n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734, 
      n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743, 
      n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752, 
      n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761, 
      n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, 
      n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779, 
      n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788, 
      n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797, 
      n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, 
      n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815, 
      n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824, 
      n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833, 
      n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842, 
      n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851, 
      n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860, 
      n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869, 
      n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, 
      n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, 
      n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, 
      n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, 
      n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, 
      n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923, 
      n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932, 
      n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941, 
      n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, 
      n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, 
      n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968, 
      n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977, 
      n25978, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, 
      n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, 
      n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, 
      n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, 
      n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, 
      n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, 
      n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, 
      n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, 
      n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, 
      n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, 
      n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, 
      n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, 
      n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, 
      n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, 
      n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, 
      n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, 
      n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, 
      n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, 
      n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, 
      n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, 
      n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, 
      n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, 
      n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, 
      n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, 
      n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, 
      n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, 
      n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, 
      n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, 
      n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, 
      n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, 
      n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, 
      n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, 
      n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, 
      n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, 
      n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, 
      n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, 
      n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, 
      n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, 
      n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, 
      n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, 
      n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, 
      n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, 
      n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, 
      n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, 
      n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, 
      n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, 
      n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, 
      n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, 
      n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, 
      n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, 
      n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, 
      n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, 
      n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, 
      n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, 
      n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, 
      n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, 
      n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, 
      n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, 
      n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, 
      n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, 
      n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, 
      n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, 
      n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, 
      n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, 
      n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, 
      n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, 
      n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, 
      n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, 
      n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, 
      n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, 
      n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, 
      n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, 
      n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, 
      n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, 
      n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, 
      n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, 
      n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, 
      n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, 
      n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, 
      n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, 
      n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, 
      n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, 
      n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, 
      n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, 
      n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, 
      n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, 
      n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, 
      n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, 
      n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, 
      n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, 
      n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, 
      n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, 
      n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, 
      n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, 
      n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, 
      n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, 
      n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, 
      n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, 
      n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, 
      n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, 
      n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, 
      n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, 
      n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, 
      n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, 
      n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, 
      n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, 
      n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, 
      n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, 
      n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, 
      n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, 
      n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, 
      n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, 
      n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, 
      n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, 
      n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, 
      n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, 
      n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, 
      n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, 
      n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, 
      n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, 
      n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, 
      n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, 
      n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, 
      n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, 
      n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, 
      n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, 
      n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, 
      n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, 
      n_2151 : std_logic;

begin
   OUT1 <= ( OUT1_63_port, OUT1_62_port, OUT1_61_port, OUT1_60_port, 
      OUT1_59_port, OUT1_58_port, OUT1_57_port, OUT1_56_port, OUT1_55_port, 
      OUT1_54_port, OUT1_53_port, OUT1_52_port, OUT1_51_port, OUT1_50_port, 
      OUT1_49_port, OUT1_48_port, OUT1_47_port, OUT1_46_port, OUT1_45_port, 
      OUT1_44_port, OUT1_43_port, OUT1_42_port, OUT1_41_port, OUT1_40_port, 
      OUT1_39_port, OUT1_38_port, OUT1_37_port, OUT1_36_port, OUT1_35_port, 
      OUT1_34_port, OUT1_33_port, OUT1_32_port, OUT1_31_port, OUT1_30_port, 
      OUT1_29_port, OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, 
      OUT1_24_port, OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, 
      OUT1_19_port, OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, 
      OUT1_14_port, OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, 
      OUT1_9_port, OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, 
      OUT1_4_port, OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_63_port, OUT2_62_port, OUT2_61_port, OUT2_60_port, 
      OUT2_59_port, OUT2_58_port, OUT2_57_port, OUT2_56_port, OUT2_55_port, 
      OUT2_54_port, OUT2_53_port, OUT2_52_port, OUT2_51_port, OUT2_50_port, 
      OUT2_49_port, OUT2_48_port, OUT2_47_port, OUT2_46_port, OUT2_45_port, 
      OUT2_44_port, OUT2_43_port, OUT2_42_port, OUT2_41_port, OUT2_40_port, 
      OUT2_39_port, OUT2_38_port, OUT2_37_port, OUT2_36_port, OUT2_35_port, 
      OUT2_34_port, OUT2_33_port, OUT2_32_port, OUT2_31_port, OUT2_30_port, 
      OUT2_29_port, OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, 
      OUT2_24_port, OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, 
      OUT2_19_port, OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, 
      OUT2_14_port, OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, 
      OUT2_9_port, OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, 
      OUT2_4_port, OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   OUT1_reg_63_inst : DFF_X1 port map( D => n5438, CK => CLK, Q => OUT1_63_port
                           , QN => n_1000);
   OUT1_reg_62_inst : DFF_X1 port map( D => n5437, CK => CLK, Q => OUT1_62_port
                           , QN => n_1001);
   OUT1_reg_61_inst : DFF_X1 port map( D => n5436, CK => CLK, Q => OUT1_61_port
                           , QN => n_1002);
   OUT1_reg_60_inst : DFF_X1 port map( D => n5435, CK => CLK, Q => OUT1_60_port
                           , QN => n_1003);
   OUT1_reg_59_inst : DFF_X1 port map( D => n5434, CK => CLK, Q => OUT1_59_port
                           , QN => n_1004);
   OUT1_reg_58_inst : DFF_X1 port map( D => n5433, CK => CLK, Q => OUT1_58_port
                           , QN => n_1005);
   OUT1_reg_57_inst : DFF_X1 port map( D => n5432, CK => CLK, Q => OUT1_57_port
                           , QN => n_1006);
   OUT1_reg_56_inst : DFF_X1 port map( D => n5431, CK => CLK, Q => OUT1_56_port
                           , QN => n_1007);
   OUT1_reg_55_inst : DFF_X1 port map( D => n5430, CK => CLK, Q => OUT1_55_port
                           , QN => n_1008);
   OUT1_reg_54_inst : DFF_X1 port map( D => n5429, CK => CLK, Q => OUT1_54_port
                           , QN => n_1009);
   OUT1_reg_53_inst : DFF_X1 port map( D => n5428, CK => CLK, Q => OUT1_53_port
                           , QN => n_1010);
   OUT1_reg_52_inst : DFF_X1 port map( D => n5427, CK => CLK, Q => OUT1_52_port
                           , QN => n_1011);
   OUT1_reg_51_inst : DFF_X1 port map( D => n5426, CK => CLK, Q => OUT1_51_port
                           , QN => n_1012);
   OUT1_reg_50_inst : DFF_X1 port map( D => n5425, CK => CLK, Q => OUT1_50_port
                           , QN => n_1013);
   OUT1_reg_49_inst : DFF_X1 port map( D => n5424, CK => CLK, Q => OUT1_49_port
                           , QN => n_1014);
   OUT1_reg_48_inst : DFF_X1 port map( D => n5423, CK => CLK, Q => OUT1_48_port
                           , QN => n_1015);
   OUT1_reg_47_inst : DFF_X1 port map( D => n5422, CK => CLK, Q => OUT1_47_port
                           , QN => n_1016);
   OUT1_reg_46_inst : DFF_X1 port map( D => n5421, CK => CLK, Q => OUT1_46_port
                           , QN => n_1017);
   OUT1_reg_45_inst : DFF_X1 port map( D => n5420, CK => CLK, Q => OUT1_45_port
                           , QN => n_1018);
   OUT1_reg_44_inst : DFF_X1 port map( D => n5419, CK => CLK, Q => OUT1_44_port
                           , QN => n_1019);
   OUT1_reg_43_inst : DFF_X1 port map( D => n5418, CK => CLK, Q => OUT1_43_port
                           , QN => n_1020);
   OUT1_reg_42_inst : DFF_X1 port map( D => n5417, CK => CLK, Q => OUT1_42_port
                           , QN => n_1021);
   OUT1_reg_41_inst : DFF_X1 port map( D => n5416, CK => CLK, Q => OUT1_41_port
                           , QN => n_1022);
   OUT1_reg_40_inst : DFF_X1 port map( D => n5415, CK => CLK, Q => OUT1_40_port
                           , QN => n_1023);
   OUT1_reg_39_inst : DFF_X1 port map( D => n5414, CK => CLK, Q => OUT1_39_port
                           , QN => n_1024);
   OUT1_reg_38_inst : DFF_X1 port map( D => n5413, CK => CLK, Q => OUT1_38_port
                           , QN => n_1025);
   OUT1_reg_37_inst : DFF_X1 port map( D => n5412, CK => CLK, Q => OUT1_37_port
                           , QN => n_1026);
   OUT1_reg_36_inst : DFF_X1 port map( D => n5411, CK => CLK, Q => OUT1_36_port
                           , QN => n_1027);
   OUT1_reg_35_inst : DFF_X1 port map( D => n5410, CK => CLK, Q => OUT1_35_port
                           , QN => n_1028);
   OUT1_reg_34_inst : DFF_X1 port map( D => n5409, CK => CLK, Q => OUT1_34_port
                           , QN => n_1029);
   OUT1_reg_33_inst : DFF_X1 port map( D => n5408, CK => CLK, Q => OUT1_33_port
                           , QN => n_1030);
   OUT1_reg_32_inst : DFF_X1 port map( D => n5407, CK => CLK, Q => OUT1_32_port
                           , QN => n_1031);
   OUT1_reg_31_inst : DFF_X1 port map( D => n5406, CK => CLK, Q => OUT1_31_port
                           , QN => n_1032);
   OUT1_reg_30_inst : DFF_X1 port map( D => n5405, CK => CLK, Q => OUT1_30_port
                           , QN => n_1033);
   OUT1_reg_29_inst : DFF_X1 port map( D => n5404, CK => CLK, Q => OUT1_29_port
                           , QN => n_1034);
   OUT1_reg_28_inst : DFF_X1 port map( D => n5403, CK => CLK, Q => OUT1_28_port
                           , QN => n_1035);
   OUT1_reg_27_inst : DFF_X1 port map( D => n5402, CK => CLK, Q => OUT1_27_port
                           , QN => n_1036);
   OUT1_reg_26_inst : DFF_X1 port map( D => n5401, CK => CLK, Q => OUT1_26_port
                           , QN => n_1037);
   OUT1_reg_25_inst : DFF_X1 port map( D => n5400, CK => CLK, Q => OUT1_25_port
                           , QN => n_1038);
   OUT1_reg_24_inst : DFF_X1 port map( D => n5399, CK => CLK, Q => OUT1_24_port
                           , QN => n_1039);
   OUT1_reg_23_inst : DFF_X1 port map( D => n5398, CK => CLK, Q => OUT1_23_port
                           , QN => n_1040);
   OUT1_reg_22_inst : DFF_X1 port map( D => n5397, CK => CLK, Q => OUT1_22_port
                           , QN => n_1041);
   OUT1_reg_21_inst : DFF_X1 port map( D => n5396, CK => CLK, Q => OUT1_21_port
                           , QN => n_1042);
   OUT1_reg_20_inst : DFF_X1 port map( D => n5395, CK => CLK, Q => OUT1_20_port
                           , QN => n_1043);
   OUT1_reg_19_inst : DFF_X1 port map( D => n5394, CK => CLK, Q => OUT1_19_port
                           , QN => n_1044);
   OUT1_reg_18_inst : DFF_X1 port map( D => n5393, CK => CLK, Q => OUT1_18_port
                           , QN => n_1045);
   OUT1_reg_17_inst : DFF_X1 port map( D => n5392, CK => CLK, Q => OUT1_17_port
                           , QN => n_1046);
   OUT1_reg_16_inst : DFF_X1 port map( D => n5391, CK => CLK, Q => OUT1_16_port
                           , QN => n_1047);
   OUT1_reg_15_inst : DFF_X1 port map( D => n5390, CK => CLK, Q => OUT1_15_port
                           , QN => n_1048);
   OUT1_reg_14_inst : DFF_X1 port map( D => n5389, CK => CLK, Q => OUT1_14_port
                           , QN => n_1049);
   OUT1_reg_13_inst : DFF_X1 port map( D => n5388, CK => CLK, Q => OUT1_13_port
                           , QN => n_1050);
   OUT1_reg_12_inst : DFF_X1 port map( D => n5387, CK => CLK, Q => OUT1_12_port
                           , QN => n_1051);
   OUT1_reg_11_inst : DFF_X1 port map( D => n5386, CK => CLK, Q => OUT1_11_port
                           , QN => n_1052);
   OUT1_reg_10_inst : DFF_X1 port map( D => n5385, CK => CLK, Q => OUT1_10_port
                           , QN => n_1053);
   OUT1_reg_9_inst : DFF_X1 port map( D => n5384, CK => CLK, Q => OUT1_9_port, 
                           QN => n_1054);
   OUT1_reg_8_inst : DFF_X1 port map( D => n5383, CK => CLK, Q => OUT1_8_port, 
                           QN => n_1055);
   OUT1_reg_7_inst : DFF_X1 port map( D => n5382, CK => CLK, Q => OUT1_7_port, 
                           QN => n_1056);
   OUT1_reg_6_inst : DFF_X1 port map( D => n5381, CK => CLK, Q => OUT1_6_port, 
                           QN => n_1057);
   OUT1_reg_5_inst : DFF_X1 port map( D => n5380, CK => CLK, Q => OUT1_5_port, 
                           QN => n_1058);
   OUT1_reg_4_inst : DFF_X1 port map( D => n5379, CK => CLK, Q => OUT1_4_port, 
                           QN => n_1059);
   OUT1_reg_3_inst : DFF_X1 port map( D => n5378, CK => CLK, Q => OUT1_3_port, 
                           QN => n_1060);
   OUT1_reg_2_inst : DFF_X1 port map( D => n5377, CK => CLK, Q => OUT1_2_port, 
                           QN => n_1061);
   OUT1_reg_1_inst : DFF_X1 port map( D => n5376, CK => CLK, Q => OUT1_1_port, 
                           QN => n_1062);
   OUT1_reg_0_inst : DFF_X1 port map( D => n5375, CK => CLK, Q => OUT1_0_port, 
                           QN => n_1063);
   OUT2_reg_62_inst : DFF_X1 port map( D => n5373, CK => CLK, Q => OUT2_62_port
                           , QN => n_1064);
   OUT2_reg_61_inst : DFF_X1 port map( D => n5372, CK => CLK, Q => OUT2_61_port
                           , QN => n_1065);
   OUT2_reg_60_inst : DFF_X1 port map( D => n5371, CK => CLK, Q => OUT2_60_port
                           , QN => n_1066);
   OUT2_reg_59_inst : DFF_X1 port map( D => n5370, CK => CLK, Q => OUT2_59_port
                           , QN => n_1067);
   OUT2_reg_58_inst : DFF_X1 port map( D => n5369, CK => CLK, Q => OUT2_58_port
                           , QN => n_1068);
   OUT2_reg_57_inst : DFF_X1 port map( D => n5368, CK => CLK, Q => OUT2_57_port
                           , QN => n_1069);
   OUT2_reg_56_inst : DFF_X1 port map( D => n5367, CK => CLK, Q => OUT2_56_port
                           , QN => n_1070);
   OUT2_reg_55_inst : DFF_X1 port map( D => n5366, CK => CLK, Q => OUT2_55_port
                           , QN => n_1071);
   OUT2_reg_54_inst : DFF_X1 port map( D => n5365, CK => CLK, Q => OUT2_54_port
                           , QN => n_1072);
   OUT2_reg_53_inst : DFF_X1 port map( D => n5364, CK => CLK, Q => OUT2_53_port
                           , QN => n_1073);
   OUT2_reg_52_inst : DFF_X1 port map( D => n5363, CK => CLK, Q => OUT2_52_port
                           , QN => n_1074);
   OUT2_reg_51_inst : DFF_X1 port map( D => n5362, CK => CLK, Q => OUT2_51_port
                           , QN => n_1075);
   OUT2_reg_50_inst : DFF_X1 port map( D => n5361, CK => CLK, Q => OUT2_50_port
                           , QN => n_1076);
   OUT2_reg_49_inst : DFF_X1 port map( D => n5360, CK => CLK, Q => OUT2_49_port
                           , QN => n_1077);
   OUT2_reg_48_inst : DFF_X1 port map( D => n5359, CK => CLK, Q => OUT2_48_port
                           , QN => n_1078);
   OUT2_reg_47_inst : DFF_X1 port map( D => n5358, CK => CLK, Q => OUT2_47_port
                           , QN => n_1079);
   OUT2_reg_46_inst : DFF_X1 port map( D => n5357, CK => CLK, Q => OUT2_46_port
                           , QN => n_1080);
   OUT2_reg_45_inst : DFF_X1 port map( D => n5356, CK => CLK, Q => OUT2_45_port
                           , QN => n_1081);
   OUT2_reg_44_inst : DFF_X1 port map( D => n5355, CK => CLK, Q => OUT2_44_port
                           , QN => n_1082);
   OUT2_reg_43_inst : DFF_X1 port map( D => n5354, CK => CLK, Q => OUT2_43_port
                           , QN => n_1083);
   OUT2_reg_42_inst : DFF_X1 port map( D => n5353, CK => CLK, Q => OUT2_42_port
                           , QN => n_1084);
   OUT2_reg_41_inst : DFF_X1 port map( D => n5352, CK => CLK, Q => OUT2_41_port
                           , QN => n_1085);
   OUT2_reg_40_inst : DFF_X1 port map( D => n5351, CK => CLK, Q => OUT2_40_port
                           , QN => n_1086);
   OUT2_reg_39_inst : DFF_X1 port map( D => n5350, CK => CLK, Q => OUT2_39_port
                           , QN => n_1087);
   OUT2_reg_38_inst : DFF_X1 port map( D => n5349, CK => CLK, Q => OUT2_38_port
                           , QN => n_1088);
   OUT2_reg_37_inst : DFF_X1 port map( D => n5348, CK => CLK, Q => OUT2_37_port
                           , QN => n_1089);
   OUT2_reg_36_inst : DFF_X1 port map( D => n5347, CK => CLK, Q => OUT2_36_port
                           , QN => n_1090);
   OUT2_reg_35_inst : DFF_X1 port map( D => n5346, CK => CLK, Q => OUT2_35_port
                           , QN => n_1091);
   OUT2_reg_34_inst : DFF_X1 port map( D => n5345, CK => CLK, Q => OUT2_34_port
                           , QN => n_1092);
   OUT2_reg_33_inst : DFF_X1 port map( D => n5344, CK => CLK, Q => OUT2_33_port
                           , QN => n_1093);
   OUT2_reg_32_inst : DFF_X1 port map( D => n5343, CK => CLK, Q => OUT2_32_port
                           , QN => n_1094);
   OUT2_reg_31_inst : DFF_X1 port map( D => n5342, CK => CLK, Q => OUT2_31_port
                           , QN => n_1095);
   OUT2_reg_30_inst : DFF_X1 port map( D => n5341, CK => CLK, Q => OUT2_30_port
                           , QN => n_1096);
   OUT2_reg_29_inst : DFF_X1 port map( D => n5340, CK => CLK, Q => OUT2_29_port
                           , QN => n_1097);
   OUT2_reg_28_inst : DFF_X1 port map( D => n5339, CK => CLK, Q => OUT2_28_port
                           , QN => n_1098);
   OUT2_reg_27_inst : DFF_X1 port map( D => n5338, CK => CLK, Q => OUT2_27_port
                           , QN => n_1099);
   OUT2_reg_26_inst : DFF_X1 port map( D => n5337, CK => CLK, Q => OUT2_26_port
                           , QN => n_1100);
   OUT2_reg_25_inst : DFF_X1 port map( D => n5336, CK => CLK, Q => OUT2_25_port
                           , QN => n_1101);
   OUT2_reg_24_inst : DFF_X1 port map( D => n5335, CK => CLK, Q => OUT2_24_port
                           , QN => n_1102);
   OUT2_reg_23_inst : DFF_X1 port map( D => n5334, CK => CLK, Q => OUT2_23_port
                           , QN => n_1103);
   OUT2_reg_22_inst : DFF_X1 port map( D => n5333, CK => CLK, Q => OUT2_22_port
                           , QN => n_1104);
   OUT2_reg_21_inst : DFF_X1 port map( D => n5332, CK => CLK, Q => OUT2_21_port
                           , QN => n_1105);
   OUT2_reg_20_inst : DFF_X1 port map( D => n5331, CK => CLK, Q => OUT2_20_port
                           , QN => n_1106);
   OUT2_reg_19_inst : DFF_X1 port map( D => n5330, CK => CLK, Q => OUT2_19_port
                           , QN => n_1107);
   OUT2_reg_18_inst : DFF_X1 port map( D => n5329, CK => CLK, Q => OUT2_18_port
                           , QN => n_1108);
   OUT2_reg_17_inst : DFF_X1 port map( D => n5328, CK => CLK, Q => OUT2_17_port
                           , QN => n_1109);
   OUT2_reg_16_inst : DFF_X1 port map( D => n5327, CK => CLK, Q => OUT2_16_port
                           , QN => n_1110);
   OUT2_reg_15_inst : DFF_X1 port map( D => n5326, CK => CLK, Q => OUT2_15_port
                           , QN => n_1111);
   OUT2_reg_14_inst : DFF_X1 port map( D => n5325, CK => CLK, Q => OUT2_14_port
                           , QN => n_1112);
   OUT2_reg_13_inst : DFF_X1 port map( D => n5324, CK => CLK, Q => OUT2_13_port
                           , QN => n_1113);
   OUT2_reg_12_inst : DFF_X1 port map( D => n5323, CK => CLK, Q => OUT2_12_port
                           , QN => n_1114);
   OUT2_reg_11_inst : DFF_X1 port map( D => n5322, CK => CLK, Q => OUT2_11_port
                           , QN => n_1115);
   OUT2_reg_10_inst : DFF_X1 port map( D => n5321, CK => CLK, Q => OUT2_10_port
                           , QN => n_1116);
   OUT2_reg_9_inst : DFF_X1 port map( D => n5320, CK => CLK, Q => OUT2_9_port, 
                           QN => n_1117);
   OUT2_reg_8_inst : DFF_X1 port map( D => n5319, CK => CLK, Q => OUT2_8_port, 
                           QN => n_1118);
   OUT2_reg_7_inst : DFF_X1 port map( D => n5318, CK => CLK, Q => OUT2_7_port, 
                           QN => n_1119);
   OUT2_reg_6_inst : DFF_X1 port map( D => n5317, CK => CLK, Q => OUT2_6_port, 
                           QN => n_1120);
   OUT2_reg_5_inst : DFF_X1 port map( D => n5316, CK => CLK, Q => OUT2_5_port, 
                           QN => n_1121);
   OUT2_reg_4_inst : DFF_X1 port map( D => n5315, CK => CLK, Q => OUT2_4_port, 
                           QN => n_1122);
   OUT2_reg_3_inst : DFF_X1 port map( D => n5314, CK => CLK, Q => OUT2_3_port, 
                           QN => n_1123);
   OUT2_reg_2_inst : DFF_X1 port map( D => n5313, CK => CLK, Q => OUT2_2_port, 
                           QN => n_1124);
   OUT2_reg_1_inst : DFF_X1 port map( D => n5312, CK => CLK, Q => OUT2_1_port, 
                           QN => n_1125);
   OUT2_reg_0_inst : DFF_X1 port map( D => n5311, CK => CLK, Q => OUT2_0_port, 
                           QN => n_1126);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n7486, CK => CLK, Q => 
                           n_1127, QN => n9415);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n7485, CK => CLK, Q => 
                           n_1128, QN => n9416);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n7484, CK => CLK, Q => 
                           n_1129, QN => n9417);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n7483, CK => CLK, Q => 
                           n_1130, QN => n9418);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n7482, CK => CLK, Q => 
                           n_1131, QN => n9419);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n7481, CK => CLK, Q => 
                           n_1132, QN => n9420);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n7480, CK => CLK, Q => 
                           n_1133, QN => n9421);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n7479, CK => CLK, Q => 
                           n_1134, QN => n9422);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n7478, CK => CLK, Q => 
                           n_1135, QN => n9423);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n7477, CK => CLK, Q => 
                           n_1136, QN => n9424);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n7476, CK => CLK, Q => 
                           n_1137, QN => n9425);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n7475, CK => CLK, Q => 
                           n_1138, QN => n9426);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n7474, CK => CLK, Q => 
                           n_1139, QN => n9427);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n7473, CK => CLK, Q => 
                           n_1140, QN => n9428);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n7472, CK => CLK, Q => 
                           n_1141, QN => n9429);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n7471, CK => CLK, Q => 
                           n_1142, QN => n9430);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n7470, CK => CLK, Q => 
                           n_1143, QN => n9431);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n7469, CK => CLK, Q => 
                           n_1144, QN => n9432);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n7468, CK => CLK, Q => 
                           n_1145, QN => n9433);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n7467, CK => CLK, Q => 
                           n_1146, QN => n9434);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n7466, CK => CLK, Q => 
                           n_1147, QN => n9435);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n7465, CK => CLK, Q => 
                           n_1148, QN => n9436);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n7464, CK => CLK, Q => 
                           n_1149, QN => n9437);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n7463, CK => CLK, Q => 
                           n_1150, QN => n9438);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n7462, CK => CLK, Q => 
                           n_1151, QN => n9439);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n7461, CK => CLK, Q => 
                           n_1152, QN => n9440);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n7460, CK => CLK, Q => 
                           n_1153, QN => n9441);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n7459, CK => CLK, Q => 
                           n_1154, QN => n9442);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n7458, CK => CLK, Q => 
                           n_1155, QN => n9443);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n7457, CK => CLK, Q => 
                           n_1156, QN => n9444);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n7456, CK => CLK, Q => 
                           n_1157, QN => n9445);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n7455, CK => CLK, Q => 
                           n_1158, QN => n9446);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n7454, CK => CLK, Q => 
                           n_1159, QN => n9447);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n7453, CK => CLK, Q => 
                           n_1160, QN => n9448);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n7452, CK => CLK, Q => 
                           n_1161, QN => n9449);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n7451, CK => CLK, Q => 
                           n_1162, QN => n9450);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n7450, CK => CLK, Q => 
                           n_1163, QN => n9451);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n7449, CK => CLK, Q => 
                           n_1164, QN => n9452);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n7448, CK => CLK, Q => 
                           n_1165, QN => n9453);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n7447, CK => CLK, Q => 
                           n_1166, QN => n9454);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n7446, CK => CLK, Q => 
                           n_1167, QN => n9455);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n7445, CK => CLK, Q => 
                           n_1168, QN => n9456);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n7444, CK => CLK, Q => 
                           n_1169, QN => n9457);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n7443, CK => CLK, Q => 
                           n_1170, QN => n9458);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n7442, CK => CLK, Q => 
                           n_1171, QN => n9459);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n7441, CK => CLK, Q => 
                           n_1172, QN => n9460);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n7440, CK => CLK, Q => 
                           n_1173, QN => n9461);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n7439, CK => CLK, Q => 
                           n_1174, QN => n9462);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n7438, CK => CLK, Q => 
                           n_1175, QN => n9463);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n7437, CK => CLK, Q => 
                           n_1176, QN => n9464);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n7436, CK => CLK, Q => 
                           n_1177, QN => n9465);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n7435, CK => CLK, Q => 
                           n_1178, QN => n9466);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n7434, CK => CLK, Q => 
                           n_1179, QN => n9467);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n7433, CK => CLK, Q => 
                           n_1180, QN => n9468);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n7432, CK => CLK, Q => n_1181
                           , QN => n9469);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n7431, CK => CLK, Q => n_1182
                           , QN => n9470);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n7430, CK => CLK, Q => n_1183
                           , QN => n9471);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n7429, CK => CLK, Q => n_1184
                           , QN => n9472);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n7428, CK => CLK, Q => n_1185
                           , QN => n9473);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n7427, CK => CLK, Q => n_1186
                           , QN => n9474);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n7426, CK => CLK, Q => n_1187
                           , QN => n9475);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n7425, CK => CLK, Q => n_1188
                           , QN => n9476);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n7424, CK => CLK, Q => n_1189
                           , QN => n9477);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n7423, CK => CLK, Q => n_1190
                           , QN => n9478);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => n6141, CK => CLK, Q => 
                           n_1191, QN => n8968);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => n6140, CK => CLK, Q => 
                           n_1192, QN => n8969);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => n6139, CK => CLK, Q => 
                           n_1193, QN => n8970);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => n6138, CK => CLK, Q => 
                           n_1194, QN => n8971);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => n6137, CK => CLK, Q => 
                           n_1195, QN => n8972);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => n6136, CK => CLK, Q => 
                           n_1196, QN => n8973);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => n6135, CK => CLK, Q => 
                           n_1197, QN => n8974);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => n6134, CK => CLK, Q => 
                           n_1198, QN => n8975);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => n6133, CK => CLK, Q => 
                           n_1199, QN => n8976);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => n6132, CK => CLK, Q => 
                           n_1200, QN => n8977);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => n6131, CK => CLK, Q => 
                           n_1201, QN => n8978);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => n6130, CK => CLK, Q => 
                           n_1202, QN => n8979);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => n6129, CK => CLK, Q => 
                           n_1203, QN => n8980);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => n6128, CK => CLK, Q => 
                           n_1204, QN => n8981);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => n6127, CK => CLK, Q => 
                           n_1205, QN => n8982);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => n6126, CK => CLK, Q => 
                           n_1206, QN => n8983);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => n6125, CK => CLK, Q => 
                           n_1207, QN => n8984);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => n6124, CK => CLK, Q => 
                           n_1208, QN => n8985);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => n6123, CK => CLK, Q => 
                           n_1209, QN => n8986);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => n6122, CK => CLK, Q => 
                           n_1210, QN => n8987);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => n6121, CK => CLK, Q => 
                           n_1211, QN => n8988);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => n6120, CK => CLK, Q => 
                           n_1212, QN => n8989);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => n6119, CK => CLK, Q => 
                           n_1213, QN => n8990);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => n6118, CK => CLK, Q => 
                           n_1214, QN => n8991);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => n6117, CK => CLK, Q => 
                           n_1215, QN => n8992);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => n6116, CK => CLK, Q => 
                           n_1216, QN => n8993);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => n6115, CK => CLK, Q => 
                           n_1217, QN => n8994);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => n6114, CK => CLK, Q => 
                           n_1218, QN => n8995);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => n6113, CK => CLK, Q => 
                           n_1219, QN => n8996);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => n6112, CK => CLK, Q => 
                           n_1220, QN => n8997);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => n6111, CK => CLK, Q => 
                           n_1221, QN => n8998);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n6110, CK => CLK, Q => 
                           n_1222, QN => n8999);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n6109, CK => CLK, Q => 
                           n_1223, QN => n9000);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n6108, CK => CLK, Q => 
                           n_1224, QN => n9001);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n6107, CK => CLK, Q => 
                           n_1225, QN => n9002);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n6106, CK => CLK, Q => 
                           n_1226, QN => n9003);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n6105, CK => CLK, Q => 
                           n_1227, QN => n9004);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n6104, CK => CLK, Q => 
                           n_1228, QN => n9005);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n6103, CK => CLK, Q => 
                           n_1229, QN => n9006);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n6102, CK => CLK, Q => 
                           n_1230, QN => n9007);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n6101, CK => CLK, Q => 
                           n_1231, QN => n9008);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n6100, CK => CLK, Q => 
                           n_1232, QN => n9009);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n6099, CK => CLK, Q => 
                           n_1233, QN => n9010);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n6098, CK => CLK, Q => 
                           n_1234, QN => n9011);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n6097, CK => CLK, Q => 
                           n_1235, QN => n9012);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n6096, CK => CLK, Q => 
                           n_1236, QN => n9013);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n6095, CK => CLK, Q => 
                           n_1237, QN => n9014);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n6094, CK => CLK, Q => 
                           n_1238, QN => n9015);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n6093, CK => CLK, Q => 
                           n_1239, QN => n9016);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n6092, CK => CLK, Q => 
                           n_1240, QN => n9017);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n6091, CK => CLK, Q => 
                           n_1241, QN => n9018);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n6090, CK => CLK, Q => 
                           n_1242, QN => n9019);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n6089, CK => CLK, Q => 
                           n_1243, QN => n9020);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n6088, CK => CLK, Q => 
                           n_1244, QN => n9021);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n6087, CK => CLK, Q => 
                           n_1245, QN => n9022);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n6086, CK => CLK, Q => 
                           n_1246, QN => n9023);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n6085, CK => CLK, Q => 
                           n_1247, QN => n9024);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n6084, CK => CLK, Q => 
                           n_1248, QN => n9025);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n6083, CK => CLK, Q => 
                           n_1249, QN => n9026);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n6082, CK => CLK, Q => 
                           n_1250, QN => n9027);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n6081, CK => CLK, Q => 
                           n_1251, QN => n9028);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n6080, CK => CLK, Q => 
                           n_1252, QN => n9029);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n6079, CK => CLK, Q => 
                           n_1253, QN => n9030);
   U15207 : NOR3_X2 port map( A1 => n25244, A2 => ADD_RD1(1), A3 => n19486, ZN 
                           => n22733);
   U16467 : NOR3_X2 port map( A1 => n25046, A2 => ADD_RD2(1), A3 => n19491, ZN 
                           => n23930);
   U18471 : NAND3_X1 port map( A1 => n19481, A2 => n19480, A3 => n21491, ZN => 
                           n21480);
   U18472 : NAND3_X1 port map( A1 => n21491, A2 => n19480, A3 => ADD_WR(2), ZN 
                           => n21494);
   U18473 : NAND3_X1 port map( A1 => n21491, A2 => n19481, A3 => ADD_WR(3), ZN 
                           => n21503);
   U18474 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n21491, A3 => ADD_WR(3), 
                           ZN => n21512);
   U18475 : NAND3_X1 port map( A1 => n19481, A2 => n19480, A3 => n21528, ZN => 
                           n21521);
   U18476 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n19480, A3 => n21528, ZN 
                           => n21531);
   U18477 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n19481, A3 => n21528, ZN 
                           => n21540);
   U18478 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), A3 => n21528, 
                           ZN => n21549);
   U18479 : NAND3_X1 port map( A1 => ENABLE, A2 => n25978, A3 => RD1, ZN => 
                           n21591);
   U18480 : NAND3_X1 port map( A1 => ENABLE, A2 => n25978, A3 => RD2, ZN => 
                           n22788);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => n7038, CK => CLK, Q => 
                           n19941, QN => n9287);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => n7037, CK => CLK, Q => 
                           n19942, QN => n9288);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => n7036, CK => CLK, Q => 
                           n19943, QN => n9289);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => n7035, CK => CLK, Q => 
                           n19944, QN => n9290);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => n7034, CK => CLK, Q => 
                           n19945, QN => n9291);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => n7033, CK => CLK, Q => 
                           n19946, QN => n9292);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => n7032, CK => CLK, Q => 
                           n19947, QN => n9293);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => n7031, CK => CLK, Q => 
                           n19948, QN => n9294);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => n7030, CK => CLK, Q => 
                           n19949, QN => n9295);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => n7029, CK => CLK, Q => 
                           n19950, QN => n9296);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => n7028, CK => CLK, Q => 
                           n19951, QN => n9297);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => n7027, CK => CLK, Q => 
                           n19952, QN => n9298);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => n7026, CK => CLK, Q => 
                           n19953, QN => n9299);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => n7025, CK => CLK, Q => 
                           n19954, QN => n9300);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => n7024, CK => CLK, Q => 
                           n19955, QN => n9301);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => n7023, CK => CLK, Q => 
                           n19956, QN => n9302);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => n7022, CK => CLK, Q => 
                           n19957, QN => n9303);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => n7021, CK => CLK, Q => 
                           n19958, QN => n9304);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => n7020, CK => CLK, Q => 
                           n19959, QN => n9305);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => n7019, CK => CLK, Q => 
                           n19960, QN => n9306);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => n7018, CK => CLK, Q => 
                           n19961, QN => n9307);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => n7017, CK => CLK, Q => 
                           n19962, QN => n9308);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => n7016, CK => CLK, Q => 
                           n19963, QN => n9309);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => n7015, CK => CLK, Q => 
                           n19964, QN => n9310);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => n7014, CK => CLK, Q => 
                           n19965, QN => n9311);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => n7013, CK => CLK, Q => 
                           n19966, QN => n9312);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => n7012, CK => CLK, Q => 
                           n19967, QN => n9313);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => n7011, CK => CLK, Q => 
                           n19968, QN => n9314);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => n7010, CK => CLK, Q => 
                           n19969, QN => n9315);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => n7009, CK => CLK, Q => 
                           n19970, QN => n9316);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => n7008, CK => CLK, Q => 
                           n19971, QN => n9317);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => n7007, CK => CLK, Q => 
                           n19972, QN => n9318);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n7006, CK => CLK, Q => 
                           n19973, QN => n9319);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n7005, CK => CLK, Q => 
                           n19974, QN => n9320);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n7004, CK => CLK, Q => 
                           n19975, QN => n9321);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n7003, CK => CLK, Q => 
                           n19976, QN => n9322);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n7002, CK => CLK, Q => 
                           n19977, QN => n9323);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n7001, CK => CLK, Q => 
                           n19978, QN => n9324);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n7000, CK => CLK, Q => 
                           n19979, QN => n9325);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n6999, CK => CLK, Q => 
                           n19980, QN => n9326);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n6998, CK => CLK, Q => 
                           n19981, QN => n9327);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n6997, CK => CLK, Q => 
                           n19982, QN => n9328);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n6996, CK => CLK, Q => 
                           n19983, QN => n9329);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n6995, CK => CLK, Q => 
                           n19984, QN => n9330);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n6994, CK => CLK, Q => 
                           n19985, QN => n9331);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n6993, CK => CLK, Q => 
                           n19986, QN => n9332);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n6992, CK => CLK, Q => 
                           n19987, QN => n9333);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n6991, CK => CLK, Q => 
                           n19988, QN => n9334);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n6990, CK => CLK, Q => 
                           n19989, QN => n9335);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n6989, CK => CLK, Q => 
                           n19990, QN => n9336);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n6988, CK => CLK, Q => 
                           n19991, QN => n9337);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n6987, CK => CLK, Q => 
                           n19992, QN => n9338);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n6986, CK => CLK, Q => 
                           n19993, QN => n9339);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n6985, CK => CLK, Q => 
                           n19994, QN => n9340);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n6984, CK => CLK, Q => n19995
                           , QN => n9341);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n6983, CK => CLK, Q => n19996
                           , QN => n9342);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n6982, CK => CLK, Q => n19997
                           , QN => n9343);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n6981, CK => CLK, Q => n19998
                           , QN => n9344);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n6980, CK => CLK, Q => n19999
                           , QN => n9345);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n6979, CK => CLK, Q => n20000
                           , QN => n9346);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n6978, CK => CLK, Q => n20001
                           , QN => n9347);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n6977, CK => CLK, Q => n20002
                           , QN => n9348);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n6976, CK => CLK, Q => n20003
                           , QN => n9349);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n6975, CK => CLK, Q => n20004
                           , QN => n9350);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n7358, CK => CLK, Q => 
                           n20005, QN => n9031);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n7357, CK => CLK, Q => 
                           n20006, QN => n9032);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n7356, CK => CLK, Q => 
                           n20007, QN => n9033);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n7355, CK => CLK, Q => 
                           n20008, QN => n9034);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n7354, CK => CLK, Q => 
                           n20009, QN => n9035);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n7353, CK => CLK, Q => 
                           n20010, QN => n9036);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n7352, CK => CLK, Q => 
                           n20011, QN => n9037);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n7351, CK => CLK, Q => 
                           n20012, QN => n9038);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n7350, CK => CLK, Q => 
                           n20013, QN => n9039);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n7349, CK => CLK, Q => 
                           n20014, QN => n9040);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n7348, CK => CLK, Q => 
                           n20015, QN => n9041);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n7347, CK => CLK, Q => 
                           n20016, QN => n9042);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n7346, CK => CLK, Q => 
                           n20017, QN => n9043);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n7345, CK => CLK, Q => 
                           n20018, QN => n9044);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n7344, CK => CLK, Q => 
                           n20019, QN => n9045);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n7343, CK => CLK, Q => 
                           n20020, QN => n9046);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n7342, CK => CLK, Q => 
                           n20021, QN => n9047);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n7341, CK => CLK, Q => 
                           n20022, QN => n9048);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n7340, CK => CLK, Q => 
                           n20023, QN => n9049);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n7339, CK => CLK, Q => 
                           n20024, QN => n9050);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n7338, CK => CLK, Q => 
                           n20025, QN => n9051);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n7337, CK => CLK, Q => 
                           n20026, QN => n9052);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n7336, CK => CLK, Q => 
                           n20027, QN => n9053);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n7335, CK => CLK, Q => 
                           n20028, QN => n9054);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n7334, CK => CLK, Q => 
                           n20029, QN => n9055);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n7333, CK => CLK, Q => 
                           n20030, QN => n9056);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n7332, CK => CLK, Q => 
                           n20031, QN => n9057);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n7331, CK => CLK, Q => 
                           n20032, QN => n9058);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n7330, CK => CLK, Q => 
                           n20033, QN => n9059);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n7329, CK => CLK, Q => 
                           n20034, QN => n9060);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n7328, CK => CLK, Q => 
                           n20035, QN => n9061);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n7327, CK => CLK, Q => 
                           n20036, QN => n9062);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n7326, CK => CLK, Q => 
                           n20037, QN => n9063);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n7325, CK => CLK, Q => 
                           n20038, QN => n9064);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n7324, CK => CLK, Q => 
                           n20039, QN => n9065);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n7323, CK => CLK, Q => 
                           n20040, QN => n9066);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n7322, CK => CLK, Q => 
                           n20041, QN => n9067);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n7321, CK => CLK, Q => 
                           n20042, QN => n9068);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n7320, CK => CLK, Q => 
                           n20043, QN => n9069);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n7319, CK => CLK, Q => 
                           n20044, QN => n9070);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n7318, CK => CLK, Q => 
                           n20045, QN => n9071);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n7317, CK => CLK, Q => 
                           n20046, QN => n9072);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n7316, CK => CLK, Q => 
                           n20047, QN => n9073);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n7315, CK => CLK, Q => 
                           n20048, QN => n9074);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n7314, CK => CLK, Q => 
                           n20049, QN => n9075);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n7313, CK => CLK, Q => 
                           n20050, QN => n9076);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n7312, CK => CLK, Q => 
                           n20051, QN => n9077);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n7311, CK => CLK, Q => 
                           n20052, QN => n9078);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n7310, CK => CLK, Q => 
                           n20053, QN => n9079);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n7309, CK => CLK, Q => 
                           n20054, QN => n9080);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n7308, CK => CLK, Q => 
                           n20055, QN => n9081);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n7307, CK => CLK, Q => 
                           n20056, QN => n9082);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n7306, CK => CLK, Q => 
                           n20057, QN => n9083);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n7305, CK => CLK, Q => 
                           n20058, QN => n9084);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n7304, CK => CLK, Q => n20059
                           , QN => n9085);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n7303, CK => CLK, Q => n20060
                           , QN => n9086);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n7302, CK => CLK, Q => n20061
                           , QN => n9087);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n7301, CK => CLK, Q => n20062
                           , QN => n9088);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n7300, CK => CLK, Q => n20063
                           , QN => n9089);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n7299, CK => CLK, Q => n20064
                           , QN => n9090);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n7298, CK => CLK, Q => n20065
                           , QN => n9091);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n7297, CK => CLK, Q => n20066
                           , QN => n9092);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n7296, CK => CLK, Q => n20067
                           , QN => n9093);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n7295, CK => CLK, Q => n20068
                           , QN => n9094);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => n6526, CK => CLK, Q => 
                           n20069, QN => n9223);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => n6525, CK => CLK, Q => 
                           n20070, QN => n9224);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => n6524, CK => CLK, Q => 
                           n20071, QN => n9225);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => n6523, CK => CLK, Q => 
                           n20072, QN => n9226);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => n6522, CK => CLK, Q => 
                           n20073, QN => n9227);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => n6521, CK => CLK, Q => 
                           n20074, QN => n9228);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => n6520, CK => CLK, Q => 
                           n20075, QN => n9229);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => n6519, CK => CLK, Q => 
                           n20076, QN => n9230);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => n6518, CK => CLK, Q => 
                           n20077, QN => n9231);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => n6517, CK => CLK, Q => 
                           n20078, QN => n9232);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => n6516, CK => CLK, Q => 
                           n20079, QN => n9233);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => n6515, CK => CLK, Q => 
                           n20080, QN => n9234);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => n6514, CK => CLK, Q => 
                           n20081, QN => n9235);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => n6513, CK => CLK, Q => 
                           n20082, QN => n9236);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => n6512, CK => CLK, Q => 
                           n20083, QN => n9237);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => n6511, CK => CLK, Q => 
                           n20084, QN => n9238);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => n6510, CK => CLK, Q => 
                           n20085, QN => n9239);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => n6509, CK => CLK, Q => 
                           n20086, QN => n9240);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => n6508, CK => CLK, Q => 
                           n20087, QN => n9241);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => n6507, CK => CLK, Q => 
                           n20088, QN => n9242);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => n6506, CK => CLK, Q => 
                           n20089, QN => n9243);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => n6505, CK => CLK, Q => 
                           n20090, QN => n9244);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => n6504, CK => CLK, Q => 
                           n20091, QN => n9245);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => n6503, CK => CLK, Q => 
                           n20092, QN => n9246);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => n6502, CK => CLK, Q => 
                           n20093, QN => n9247);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => n6501, CK => CLK, Q => 
                           n20094, QN => n9248);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => n6500, CK => CLK, Q => 
                           n20095, QN => n9249);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => n6499, CK => CLK, Q => 
                           n20096, QN => n9250);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => n6498, CK => CLK, Q => 
                           n20097, QN => n9251);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => n6497, CK => CLK, Q => 
                           n20098, QN => n9252);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => n6496, CK => CLK, Q => 
                           n20099, QN => n9253);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => n6495, CK => CLK, Q => 
                           n20100, QN => n9254);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n6494, CK => CLK, Q => 
                           n20101, QN => n9255);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n6493, CK => CLK, Q => 
                           n20102, QN => n9256);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n6492, CK => CLK, Q => 
                           n20103, QN => n9257);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n6491, CK => CLK, Q => 
                           n20104, QN => n9258);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n6490, CK => CLK, Q => 
                           n20105, QN => n9259);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n6489, CK => CLK, Q => 
                           n20106, QN => n9260);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n6488, CK => CLK, Q => 
                           n20107, QN => n9261);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n6487, CK => CLK, Q => 
                           n20108, QN => n9262);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n6486, CK => CLK, Q => 
                           n20109, QN => n9263);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n6485, CK => CLK, Q => 
                           n20110, QN => n9264);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n6484, CK => CLK, Q => 
                           n20111, QN => n9265);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n6483, CK => CLK, Q => 
                           n20112, QN => n9266);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n6482, CK => CLK, Q => 
                           n20113, QN => n9267);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n6481, CK => CLK, Q => 
                           n20114, QN => n9268);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n6480, CK => CLK, Q => 
                           n20115, QN => n9269);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n6479, CK => CLK, Q => 
                           n20116, QN => n9270);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n6478, CK => CLK, Q => 
                           n20117, QN => n9271);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n6477, CK => CLK, Q => 
                           n20118, QN => n9272);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n6476, CK => CLK, Q => 
                           n20119, QN => n9273);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n6475, CK => CLK, Q => 
                           n20120, QN => n9274);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n6474, CK => CLK, Q => 
                           n20121, QN => n9275);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n6473, CK => CLK, Q => 
                           n20122, QN => n9276);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n6472, CK => CLK, Q => 
                           n20123, QN => n9277);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n6471, CK => CLK, Q => 
                           n20124, QN => n9278);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n6470, CK => CLK, Q => 
                           n20125, QN => n9279);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n6469, CK => CLK, Q => 
                           n20126, QN => n9280);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n6468, CK => CLK, Q => 
                           n20127, QN => n9281);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n6467, CK => CLK, Q => 
                           n20128, QN => n9282);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n6466, CK => CLK, Q => 
                           n20129, QN => n9283);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n6465, CK => CLK, Q => 
                           n20130, QN => n9284);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n6464, CK => CLK, Q => 
                           n20131, QN => n9285);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n6463, CK => CLK, Q => 
                           n20132, QN => n9286);
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => n6142, CK => CLK, Q => 
                           n_1254, QN => n8967);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => n5758, CK => CLK, Q => 
                           n_1255, QN => n20134);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => n5757, CK => CLK, Q => 
                           n_1256, QN => n20135);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => n5756, CK => CLK, Q => 
                           n_1257, QN => n20136);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => n5755, CK => CLK, Q => 
                           n_1258, QN => n20137);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => n5754, CK => CLK, Q => 
                           n_1259, QN => n20138);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => n5753, CK => CLK, Q => 
                           n_1260, QN => n20139);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => n5752, CK => CLK, Q => 
                           n_1261, QN => n20140);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => n5751, CK => CLK, Q => 
                           n_1262, QN => n20141);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => n5750, CK => CLK, Q => 
                           n_1263, QN => n20142);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => n5749, CK => CLK, Q => 
                           n_1264, QN => n20143);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => n5748, CK => CLK, Q => 
                           n_1265, QN => n20144);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => n5747, CK => CLK, Q => 
                           n_1266, QN => n20145);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => n5746, CK => CLK, Q => 
                           n_1267, QN => n20146);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => n5745, CK => CLK, Q => 
                           n_1268, QN => n20147);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => n5744, CK => CLK, Q => 
                           n_1269, QN => n20148);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => n5743, CK => CLK, Q => 
                           n_1270, QN => n20149);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => n5742, CK => CLK, Q => 
                           n_1271, QN => n20150);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => n5741, CK => CLK, Q => 
                           n_1272, QN => n20151);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => n5740, CK => CLK, Q => 
                           n_1273, QN => n20152);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => n5739, CK => CLK, Q => 
                           n_1274, QN => n20153);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => n5738, CK => CLK, Q => 
                           n_1275, QN => n20154);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => n5737, CK => CLK, Q => 
                           n_1276, QN => n20155);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => n5736, CK => CLK, Q => 
                           n_1277, QN => n20156);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => n5735, CK => CLK, Q => 
                           n_1278, QN => n20157);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => n5734, CK => CLK, Q => 
                           n_1279, QN => n20158);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => n5733, CK => CLK, Q => 
                           n_1280, QN => n20159);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => n5732, CK => CLK, Q => 
                           n_1281, QN => n20160);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => n5731, CK => CLK, Q => 
                           n_1282, QN => n20161);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => n5730, CK => CLK, Q => 
                           n_1283, QN => n20162);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => n5729, CK => CLK, Q => 
                           n_1284, QN => n20163);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => n5728, CK => CLK, Q => 
                           n_1285, QN => n20164);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => n5727, CK => CLK, Q => 
                           n_1286, QN => n20165);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n5726, CK => CLK, Q => 
                           n_1287, QN => n20166);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n5725, CK => CLK, Q => 
                           n_1288, QN => n20167);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n5724, CK => CLK, Q => 
                           n_1289, QN => n20168);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n5723, CK => CLK, Q => 
                           n_1290, QN => n20169);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n5722, CK => CLK, Q => 
                           n_1291, QN => n20170);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n5721, CK => CLK, Q => 
                           n_1292, QN => n20171);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n5720, CK => CLK, Q => 
                           n_1293, QN => n20172);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n5719, CK => CLK, Q => 
                           n_1294, QN => n20173);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n5718, CK => CLK, Q => 
                           n_1295, QN => n20174);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n5717, CK => CLK, Q => 
                           n_1296, QN => n20175);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n5716, CK => CLK, Q => 
                           n_1297, QN => n20176);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n5715, CK => CLK, Q => 
                           n_1298, QN => n20177);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n5714, CK => CLK, Q => 
                           n_1299, QN => n20178);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n5713, CK => CLK, Q => 
                           n_1300, QN => n20179);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n5712, CK => CLK, Q => 
                           n_1301, QN => n20180);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n5711, CK => CLK, Q => 
                           n_1302, QN => n20181);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n5710, CK => CLK, Q => 
                           n_1303, QN => n20182);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n5709, CK => CLK, Q => 
                           n_1304, QN => n20183);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n5708, CK => CLK, Q => 
                           n_1305, QN => n20184);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n5707, CK => CLK, Q => 
                           n_1306, QN => n20185);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n5706, CK => CLK, Q => 
                           n_1307, QN => n20186);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n5705, CK => CLK, Q => 
                           n_1308, QN => n20187);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n5704, CK => CLK, Q => 
                           n_1309, QN => n20188);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n5703, CK => CLK, Q => 
                           n_1310, QN => n20189);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n5702, CK => CLK, Q => 
                           n_1311, QN => n20190);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n5701, CK => CLK, Q => 
                           n_1312, QN => n20191);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n5700, CK => CLK, Q => 
                           n_1313, QN => n20192);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n5699, CK => CLK, Q => 
                           n_1314, QN => n20193);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n5698, CK => CLK, Q => 
                           n_1315, QN => n20194);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n5697, CK => CLK, Q => 
                           n_1316, QN => n20195);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n5696, CK => CLK, Q => 
                           n_1317, QN => n20196);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n5695, CK => CLK, Q => 
                           n_1318, QN => n20197);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => n7166, CK => CLK, Q => 
                           n_1319, QN => n19558);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => n7165, CK => CLK, Q => 
                           n_1320, QN => n19559);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => n7164, CK => CLK, Q => 
                           n_1321, QN => n19560);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => n7163, CK => CLK, Q => 
                           n_1322, QN => n19561);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => n7162, CK => CLK, Q => 
                           n_1323, QN => n19562);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => n7161, CK => CLK, Q => 
                           n_1324, QN => n19563);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => n7160, CK => CLK, Q => 
                           n_1325, QN => n19564);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => n7159, CK => CLK, Q => 
                           n_1326, QN => n19565);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => n7158, CK => CLK, Q => 
                           n_1327, QN => n19566);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => n7157, CK => CLK, Q => 
                           n_1328, QN => n19567);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => n7156, CK => CLK, Q => 
                           n_1329, QN => n19568);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => n7155, CK => CLK, Q => 
                           n_1330, QN => n19569);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => n7154, CK => CLK, Q => 
                           n_1331, QN => n19570);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => n7153, CK => CLK, Q => 
                           n_1332, QN => n19571);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => n7152, CK => CLK, Q => 
                           n_1333, QN => n19572);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => n7151, CK => CLK, Q => 
                           n_1334, QN => n19573);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => n7150, CK => CLK, Q => 
                           n_1335, QN => n19574);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => n7149, CK => CLK, Q => 
                           n_1336, QN => n19575);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => n7148, CK => CLK, Q => 
                           n_1337, QN => n19576);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => n7147, CK => CLK, Q => 
                           n_1338, QN => n19577);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => n7146, CK => CLK, Q => 
                           n_1339, QN => n19578);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => n7145, CK => CLK, Q => 
                           n_1340, QN => n19579);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => n7144, CK => CLK, Q => 
                           n_1341, QN => n19580);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => n7143, CK => CLK, Q => 
                           n_1342, QN => n19581);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => n7142, CK => CLK, Q => 
                           n_1343, QN => n19582);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => n7141, CK => CLK, Q => 
                           n_1344, QN => n19583);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => n7140, CK => CLK, Q => 
                           n_1345, QN => n19584);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => n7139, CK => CLK, Q => 
                           n_1346, QN => n19585);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => n7138, CK => CLK, Q => 
                           n_1347, QN => n19586);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => n7137, CK => CLK, Q => 
                           n_1348, QN => n19587);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => n7136, CK => CLK, Q => 
                           n_1349, QN => n19588);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => n7135, CK => CLK, Q => 
                           n_1350, QN => n19589);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n7134, CK => CLK, Q => 
                           n_1351, QN => n19590);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n7133, CK => CLK, Q => 
                           n_1352, QN => n19591);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n7132, CK => CLK, Q => 
                           n_1353, QN => n19592);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n7131, CK => CLK, Q => 
                           n_1354, QN => n19593);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n7130, CK => CLK, Q => 
                           n_1355, QN => n19594);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n7129, CK => CLK, Q => 
                           n_1356, QN => n19595);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n7128, CK => CLK, Q => 
                           n_1357, QN => n19596);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n7127, CK => CLK, Q => 
                           n_1358, QN => n19597);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n7126, CK => CLK, Q => 
                           n_1359, QN => n19598);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n7125, CK => CLK, Q => 
                           n_1360, QN => n19599);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n7124, CK => CLK, Q => 
                           n_1361, QN => n19600);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n7123, CK => CLK, Q => 
                           n_1362, QN => n19601);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n7122, CK => CLK, Q => 
                           n_1363, QN => n19602);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n7121, CK => CLK, Q => 
                           n_1364, QN => n19603);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n7120, CK => CLK, Q => 
                           n_1365, QN => n19604);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n7119, CK => CLK, Q => 
                           n_1366, QN => n19605);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n7118, CK => CLK, Q => 
                           n_1367, QN => n19606);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n7117, CK => CLK, Q => 
                           n_1368, QN => n19607);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n7116, CK => CLK, Q => 
                           n_1369, QN => n19608);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n7115, CK => CLK, Q => 
                           n_1370, QN => n19609);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n7114, CK => CLK, Q => 
                           n_1371, QN => n19610);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n7113, CK => CLK, Q => 
                           n_1372, QN => n19611);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n7112, CK => CLK, Q => n_1373
                           , QN => n19612);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n7111, CK => CLK, Q => n_1374
                           , QN => n19613);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n7110, CK => CLK, Q => n_1375
                           , QN => n19614);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n7109, CK => CLK, Q => n_1376
                           , QN => n19615);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n7108, CK => CLK, Q => n_1377
                           , QN => n19616);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n7107, CK => CLK, Q => n_1378
                           , QN => n19617);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n7106, CK => CLK, Q => n_1379
                           , QN => n19618);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n7105, CK => CLK, Q => n_1380
                           , QN => n19619);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n7104, CK => CLK, Q => n_1381
                           , QN => n19620);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n7103, CK => CLK, Q => n_1382
                           , QN => n19621);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n7422, CK => CLK, Q => 
                           n_1383, QN => n20966);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n7421, CK => CLK, Q => 
                           n_1384, QN => n20967);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n7420, CK => CLK, Q => 
                           n_1385, QN => n20968);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n7419, CK => CLK, Q => 
                           n_1386, QN => n20969);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n7418, CK => CLK, Q => 
                           n_1387, QN => n20970);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n7417, CK => CLK, Q => 
                           n_1388, QN => n20971);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n7416, CK => CLK, Q => 
                           n_1389, QN => n20972);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n7415, CK => CLK, Q => 
                           n_1390, QN => n20973);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n7414, CK => CLK, Q => 
                           n_1391, QN => n20974);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n7413, CK => CLK, Q => 
                           n_1392, QN => n20975);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n7412, CK => CLK, Q => 
                           n_1393, QN => n20976);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n7411, CK => CLK, Q => 
                           n_1394, QN => n20977);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n7410, CK => CLK, Q => 
                           n_1395, QN => n20978);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n7409, CK => CLK, Q => 
                           n_1396, QN => n20979);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n7408, CK => CLK, Q => 
                           n_1397, QN => n20980);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n7407, CK => CLK, Q => 
                           n_1398, QN => n20981);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n7406, CK => CLK, Q => 
                           n_1399, QN => n20982);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n7405, CK => CLK, Q => 
                           n_1400, QN => n20983);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n7404, CK => CLK, Q => 
                           n_1401, QN => n20984);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n7403, CK => CLK, Q => 
                           n_1402, QN => n20985);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n7402, CK => CLK, Q => 
                           n_1403, QN => n20986);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n7401, CK => CLK, Q => 
                           n_1404, QN => n20987);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n7400, CK => CLK, Q => 
                           n_1405, QN => n20988);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n7399, CK => CLK, Q => 
                           n_1406, QN => n20989);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n7398, CK => CLK, Q => 
                           n_1407, QN => n20990);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n7397, CK => CLK, Q => 
                           n_1408, QN => n20991);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n7396, CK => CLK, Q => 
                           n_1409, QN => n20992);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n7395, CK => CLK, Q => 
                           n_1410, QN => n20993);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n7394, CK => CLK, Q => 
                           n_1411, QN => n20994);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n7393, CK => CLK, Q => 
                           n_1412, QN => n20995);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n7392, CK => CLK, Q => 
                           n_1413, QN => n20996);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n7391, CK => CLK, Q => 
                           n_1414, QN => n20997);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n7390, CK => CLK, Q => 
                           n_1415, QN => n20998);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n7389, CK => CLK, Q => 
                           n_1416, QN => n20999);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n7388, CK => CLK, Q => 
                           n_1417, QN => n21000);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n7387, CK => CLK, Q => 
                           n_1418, QN => n21001);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n7386, CK => CLK, Q => 
                           n_1419, QN => n21002);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n7385, CK => CLK, Q => 
                           n_1420, QN => n21003);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n7384, CK => CLK, Q => 
                           n_1421, QN => n21004);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n7383, CK => CLK, Q => 
                           n_1422, QN => n21005);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n7382, CK => CLK, Q => 
                           n_1423, QN => n21006);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n7381, CK => CLK, Q => 
                           n_1424, QN => n21007);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n7380, CK => CLK, Q => 
                           n_1425, QN => n21008);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n7379, CK => CLK, Q => 
                           n_1426, QN => n21009);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n7378, CK => CLK, Q => 
                           n_1427, QN => n21010);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n7377, CK => CLK, Q => 
                           n_1428, QN => n21011);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n7376, CK => CLK, Q => 
                           n_1429, QN => n21012);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n7375, CK => CLK, Q => 
                           n_1430, QN => n21013);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n7374, CK => CLK, Q => 
                           n_1431, QN => n21014);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n7373, CK => CLK, Q => 
                           n_1432, QN => n21015);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n7372, CK => CLK, Q => 
                           n_1433, QN => n21016);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n7371, CK => CLK, Q => 
                           n_1434, QN => n21017);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n7370, CK => CLK, Q => 
                           n_1435, QN => n21018);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n7369, CK => CLK, Q => 
                           n_1436, QN => n21019);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n7368, CK => CLK, Q => n_1437
                           , QN => n21020);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n7367, CK => CLK, Q => n_1438
                           , QN => n21021);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n7366, CK => CLK, Q => n_1439
                           , QN => n21022);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n7365, CK => CLK, Q => n_1440
                           , QN => n21023);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n7364, CK => CLK, Q => n_1441
                           , QN => n21024);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n7363, CK => CLK, Q => n_1442
                           , QN => n21025);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n7362, CK => CLK, Q => n_1443
                           , QN => n21026);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n7361, CK => CLK, Q => n_1444
                           , QN => n21027);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n7360, CK => CLK, Q => n_1445
                           , QN => n21028);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n7359, CK => CLK, Q => n_1446
                           , QN => n21029);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => n6206, CK => CLK, Q => 
                           n_1447, QN => n20270);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => n6205, CK => CLK, Q => 
                           n_1448, QN => n20271);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => n6204, CK => CLK, Q => 
                           n_1449, QN => n20272);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => n6203, CK => CLK, Q => 
                           n_1450, QN => n20273);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => n6202, CK => CLK, Q => 
                           n_1451, QN => n20274);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => n6201, CK => CLK, Q => 
                           n_1452, QN => n20275);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => n6200, CK => CLK, Q => 
                           n_1453, QN => n20276);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => n6199, CK => CLK, Q => 
                           n_1454, QN => n20277);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => n6198, CK => CLK, Q => 
                           n_1455, QN => n20278);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => n6197, CK => CLK, Q => 
                           n_1456, QN => n20279);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => n6196, CK => CLK, Q => 
                           n_1457, QN => n20280);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => n6195, CK => CLK, Q => 
                           n_1458, QN => n20281);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => n6194, CK => CLK, Q => 
                           n_1459, QN => n20282);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => n6193, CK => CLK, Q => 
                           n_1460, QN => n20283);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => n6192, CK => CLK, Q => 
                           n_1461, QN => n20284);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => n6191, CK => CLK, Q => 
                           n_1462, QN => n20285);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => n6190, CK => CLK, Q => 
                           n_1463, QN => n20286);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => n6189, CK => CLK, Q => 
                           n_1464, QN => n20287);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => n6188, CK => CLK, Q => 
                           n_1465, QN => n20288);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => n6187, CK => CLK, Q => 
                           n_1466, QN => n20289);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => n6186, CK => CLK, Q => 
                           n_1467, QN => n20290);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => n6185, CK => CLK, Q => 
                           n_1468, QN => n20291);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => n6184, CK => CLK, Q => 
                           n_1469, QN => n20292);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => n6183, CK => CLK, Q => 
                           n_1470, QN => n20293);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => n6182, CK => CLK, Q => 
                           n_1471, QN => n20294);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => n6181, CK => CLK, Q => 
                           n_1472, QN => n20295);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => n6180, CK => CLK, Q => 
                           n_1473, QN => n20296);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => n6179, CK => CLK, Q => 
                           n_1474, QN => n20297);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => n6178, CK => CLK, Q => 
                           n_1475, QN => n20298);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => n6177, CK => CLK, Q => 
                           n_1476, QN => n20299);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => n6176, CK => CLK, Q => 
                           n_1477, QN => n20300);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => n6175, CK => CLK, Q => 
                           n_1478, QN => n20301);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n6174, CK => CLK, Q => 
                           n_1479, QN => n20302);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n6173, CK => CLK, Q => 
                           n_1480, QN => n20303);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n6172, CK => CLK, Q => 
                           n_1481, QN => n20304);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n6171, CK => CLK, Q => 
                           n_1482, QN => n20305);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n6170, CK => CLK, Q => 
                           n_1483, QN => n20306);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n6169, CK => CLK, Q => 
                           n_1484, QN => n20307);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n6168, CK => CLK, Q => 
                           n_1485, QN => n20308);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n6167, CK => CLK, Q => 
                           n_1486, QN => n20309);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n6166, CK => CLK, Q => 
                           n_1487, QN => n20310);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n6165, CK => CLK, Q => 
                           n_1488, QN => n20311);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n6164, CK => CLK, Q => 
                           n_1489, QN => n20312);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n6163, CK => CLK, Q => 
                           n_1490, QN => n20313);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n6162, CK => CLK, Q => 
                           n_1491, QN => n20314);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n6161, CK => CLK, Q => 
                           n_1492, QN => n20315);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n6160, CK => CLK, Q => 
                           n_1493, QN => n20316);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n6159, CK => CLK, Q => 
                           n_1494, QN => n20317);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n6158, CK => CLK, Q => 
                           n_1495, QN => n20318);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n6157, CK => CLK, Q => 
                           n_1496, QN => n20319);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n6156, CK => CLK, Q => 
                           n_1497, QN => n20320);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n6155, CK => CLK, Q => 
                           n_1498, QN => n20321);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n6154, CK => CLK, Q => 
                           n_1499, QN => n20322);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n6153, CK => CLK, Q => 
                           n_1500, QN => n20323);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n6152, CK => CLK, Q => 
                           n_1501, QN => n20324);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n6151, CK => CLK, Q => 
                           n_1502, QN => n20325);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n6150, CK => CLK, Q => 
                           n_1503, QN => n20326);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n6149, CK => CLK, Q => 
                           n_1504, QN => n20327);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n6148, CK => CLK, Q => 
                           n_1505, QN => n20328);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n6147, CK => CLK, Q => 
                           n_1506, QN => n20329);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n6146, CK => CLK, Q => 
                           n_1507, QN => n20330);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n6145, CK => CLK, Q => 
                           n_1508, QN => n20331);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n6144, CK => CLK, Q => 
                           n_1509, QN => n20332);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n6143, CK => CLK, Q => 
                           n_1510, QN => n20333);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => n6334, CK => CLK, Q => 
                           n_1511, QN => n20334);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => n6333, CK => CLK, Q => 
                           n_1512, QN => n20335);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => n6332, CK => CLK, Q => 
                           n_1513, QN => n20336);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => n6331, CK => CLK, Q => 
                           n_1514, QN => n20337);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => n6330, CK => CLK, Q => 
                           n_1515, QN => n20338);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => n6329, CK => CLK, Q => 
                           n_1516, QN => n20339);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => n6328, CK => CLK, Q => 
                           n_1517, QN => n20340);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => n6327, CK => CLK, Q => 
                           n_1518, QN => n20341);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => n6326, CK => CLK, Q => 
                           n_1519, QN => n20342);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => n6325, CK => CLK, Q => 
                           n_1520, QN => n20343);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => n6324, CK => CLK, Q => 
                           n_1521, QN => n20344);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => n6323, CK => CLK, Q => 
                           n_1522, QN => n20345);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => n6322, CK => CLK, Q => 
                           n_1523, QN => n20346);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => n6321, CK => CLK, Q => 
                           n_1524, QN => n20347);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => n6320, CK => CLK, Q => 
                           n_1525, QN => n20348);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => n6319, CK => CLK, Q => 
                           n_1526, QN => n20349);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => n6318, CK => CLK, Q => 
                           n_1527, QN => n20350);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => n6317, CK => CLK, Q => 
                           n_1528, QN => n20351);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => n6316, CK => CLK, Q => 
                           n_1529, QN => n20352);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => n6315, CK => CLK, Q => 
                           n_1530, QN => n20353);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => n6314, CK => CLK, Q => 
                           n_1531, QN => n20354);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => n6313, CK => CLK, Q => 
                           n_1532, QN => n20355);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => n6312, CK => CLK, Q => 
                           n_1533, QN => n20356);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => n6311, CK => CLK, Q => 
                           n_1534, QN => n20357);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => n6310, CK => CLK, Q => 
                           n_1535, QN => n20358);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => n6309, CK => CLK, Q => 
                           n_1536, QN => n20359);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => n6308, CK => CLK, Q => 
                           n_1537, QN => n20360);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => n6307, CK => CLK, Q => 
                           n_1538, QN => n20361);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => n6306, CK => CLK, Q => 
                           n_1539, QN => n20362);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => n6305, CK => CLK, Q => 
                           n_1540, QN => n20363);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => n6304, CK => CLK, Q => 
                           n_1541, QN => n20364);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => n6303, CK => CLK, Q => 
                           n_1542, QN => n20365);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n6302, CK => CLK, Q => 
                           n_1543, QN => n20366);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n6301, CK => CLK, Q => 
                           n_1544, QN => n20367);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n6300, CK => CLK, Q => 
                           n_1545, QN => n20368);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n6299, CK => CLK, Q => 
                           n_1546, QN => n20369);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n6298, CK => CLK, Q => 
                           n_1547, QN => n20370);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n6297, CK => CLK, Q => 
                           n_1548, QN => n20371);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n6296, CK => CLK, Q => 
                           n_1549, QN => n20372);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n6295, CK => CLK, Q => 
                           n_1550, QN => n20373);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n6294, CK => CLK, Q => 
                           n_1551, QN => n20374);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n6293, CK => CLK, Q => 
                           n_1552, QN => n20375);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n6292, CK => CLK, Q => 
                           n_1553, QN => n20376);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n6291, CK => CLK, Q => 
                           n_1554, QN => n20377);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n6290, CK => CLK, Q => 
                           n_1555, QN => n20378);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n6289, CK => CLK, Q => 
                           n_1556, QN => n20379);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n6288, CK => CLK, Q => 
                           n_1557, QN => n20380);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n6287, CK => CLK, Q => 
                           n_1558, QN => n20381);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n6286, CK => CLK, Q => 
                           n_1559, QN => n20382);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n6285, CK => CLK, Q => 
                           n_1560, QN => n20383);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n6284, CK => CLK, Q => 
                           n_1561, QN => n20384);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n6283, CK => CLK, Q => 
                           n_1562, QN => n20385);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n6282, CK => CLK, Q => 
                           n_1563, QN => n20386);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n6281, CK => CLK, Q => 
                           n_1564, QN => n20387);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n6280, CK => CLK, Q => 
                           n_1565, QN => n20388);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n6279, CK => CLK, Q => 
                           n_1566, QN => n20389);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n6278, CK => CLK, Q => 
                           n_1567, QN => n20390);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n6277, CK => CLK, Q => 
                           n_1568, QN => n20391);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n6276, CK => CLK, Q => 
                           n_1569, QN => n20392);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n6275, CK => CLK, Q => 
                           n_1570, QN => n20393);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n6274, CK => CLK, Q => 
                           n_1571, QN => n20394);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n6273, CK => CLK, Q => 
                           n_1572, QN => n20395);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n6272, CK => CLK, Q => 
                           n_1573, QN => n20396);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n6271, CK => CLK, Q => 
                           n_1574, QN => n20397);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => n6654, CK => CLK, Q => 
                           n_1575, QN => n19813);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => n6653, CK => CLK, Q => 
                           n_1576, QN => n19814);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => n6652, CK => CLK, Q => 
                           n_1577, QN => n19815);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => n6651, CK => CLK, Q => 
                           n_1578, QN => n19816);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => n6650, CK => CLK, Q => 
                           n_1579, QN => n19817);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => n6649, CK => CLK, Q => 
                           n_1580, QN => n19818);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => n6648, CK => CLK, Q => 
                           n_1581, QN => n19819);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => n6647, CK => CLK, Q => 
                           n_1582, QN => n19820);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => n6646, CK => CLK, Q => 
                           n_1583, QN => n19821);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => n6645, CK => CLK, Q => 
                           n_1584, QN => n19822);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => n6644, CK => CLK, Q => 
                           n_1585, QN => n19823);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => n6643, CK => CLK, Q => 
                           n_1586, QN => n19824);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => n6642, CK => CLK, Q => 
                           n_1587, QN => n19825);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => n6641, CK => CLK, Q => 
                           n_1588, QN => n19826);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => n6640, CK => CLK, Q => 
                           n_1589, QN => n19827);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => n6639, CK => CLK, Q => 
                           n_1590, QN => n19828);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => n6638, CK => CLK, Q => 
                           n_1591, QN => n19829);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => n6637, CK => CLK, Q => 
                           n_1592, QN => n19830);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => n6636, CK => CLK, Q => 
                           n_1593, QN => n19831);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => n6635, CK => CLK, Q => 
                           n_1594, QN => n19832);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => n6634, CK => CLK, Q => 
                           n_1595, QN => n19833);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => n6633, CK => CLK, Q => 
                           n_1596, QN => n19834);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => n6632, CK => CLK, Q => 
                           n_1597, QN => n19835);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => n6631, CK => CLK, Q => 
                           n_1598, QN => n19836);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => n6630, CK => CLK, Q => 
                           n_1599, QN => n19837);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => n6629, CK => CLK, Q => 
                           n_1600, QN => n19838);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => n6628, CK => CLK, Q => 
                           n_1601, QN => n19839);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => n6627, CK => CLK, Q => 
                           n_1602, QN => n19840);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => n6626, CK => CLK, Q => 
                           n_1603, QN => n19841);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => n6625, CK => CLK, Q => 
                           n_1604, QN => n19842);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => n6624, CK => CLK, Q => 
                           n_1605, QN => n19843);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => n6623, CK => CLK, Q => 
                           n_1606, QN => n19844);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n6622, CK => CLK, Q => 
                           n_1607, QN => n19845);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n6621, CK => CLK, Q => 
                           n_1608, QN => n19846);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n6620, CK => CLK, Q => 
                           n_1609, QN => n19847);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n6619, CK => CLK, Q => 
                           n_1610, QN => n19848);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n6618, CK => CLK, Q => 
                           n_1611, QN => n19849);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n6617, CK => CLK, Q => 
                           n_1612, QN => n19850);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n6616, CK => CLK, Q => 
                           n_1613, QN => n19851);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n6615, CK => CLK, Q => 
                           n_1614, QN => n19852);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n6614, CK => CLK, Q => 
                           n_1615, QN => n19853);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n6613, CK => CLK, Q => 
                           n_1616, QN => n19854);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n6612, CK => CLK, Q => 
                           n_1617, QN => n19855);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n6611, CK => CLK, Q => 
                           n_1618, QN => n19856);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n6610, CK => CLK, Q => 
                           n_1619, QN => n19857);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n6609, CK => CLK, Q => 
                           n_1620, QN => n19858);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n6608, CK => CLK, Q => 
                           n_1621, QN => n19859);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n6607, CK => CLK, Q => 
                           n_1622, QN => n19860);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n6606, CK => CLK, Q => 
                           n_1623, QN => n19861);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n6605, CK => CLK, Q => 
                           n_1624, QN => n19862);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n6604, CK => CLK, Q => 
                           n_1625, QN => n19863);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n6603, CK => CLK, Q => 
                           n_1626, QN => n19864);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n6602, CK => CLK, Q => 
                           n_1627, QN => n19865);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n6601, CK => CLK, Q => 
                           n_1628, QN => n19866);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n6600, CK => CLK, Q => 
                           n_1629, QN => n19867);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n6599, CK => CLK, Q => 
                           n_1630, QN => n19868);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n6598, CK => CLK, Q => 
                           n_1631, QN => n19869);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n6597, CK => CLK, Q => 
                           n_1632, QN => n19870);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n6596, CK => CLK, Q => 
                           n_1633, QN => n19871);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n6595, CK => CLK, Q => 
                           n_1634, QN => n19872);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n6594, CK => CLK, Q => 
                           n_1635, QN => n19873);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n6593, CK => CLK, Q => 
                           n_1636, QN => n19874);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n6592, CK => CLK, Q => 
                           n_1637, QN => n19875);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n6591, CK => CLK, Q => 
                           n_1638, QN => n19876);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => n6718, CK => CLK, Q => 
                           n_1639, QN => n20398);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => n6717, CK => CLK, Q => 
                           n_1640, QN => n20399);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => n6716, CK => CLK, Q => 
                           n_1641, QN => n20400);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => n6715, CK => CLK, Q => 
                           n_1642, QN => n20401);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => n6714, CK => CLK, Q => 
                           n_1643, QN => n20402);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => n6713, CK => CLK, Q => 
                           n_1644, QN => n20403);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => n6712, CK => CLK, Q => 
                           n_1645, QN => n20404);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => n6711, CK => CLK, Q => 
                           n_1646, QN => n20405);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => n6710, CK => CLK, Q => 
                           n_1647, QN => n20406);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => n6709, CK => CLK, Q => 
                           n_1648, QN => n20407);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => n6708, CK => CLK, Q => 
                           n_1649, QN => n20408);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => n6707, CK => CLK, Q => 
                           n_1650, QN => n20409);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => n6706, CK => CLK, Q => 
                           n_1651, QN => n20410);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => n6705, CK => CLK, Q => 
                           n_1652, QN => n20411);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => n6704, CK => CLK, Q => 
                           n_1653, QN => n20412);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => n6703, CK => CLK, Q => 
                           n_1654, QN => n20413);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => n6702, CK => CLK, Q => 
                           n_1655, QN => n20414);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => n6701, CK => CLK, Q => 
                           n_1656, QN => n20415);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => n6700, CK => CLK, Q => 
                           n_1657, QN => n20416);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => n6699, CK => CLK, Q => 
                           n_1658, QN => n20417);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => n6698, CK => CLK, Q => 
                           n_1659, QN => n20418);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => n6697, CK => CLK, Q => 
                           n_1660, QN => n20419);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => n6696, CK => CLK, Q => 
                           n_1661, QN => n20420);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => n6695, CK => CLK, Q => 
                           n_1662, QN => n20421);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => n6694, CK => CLK, Q => 
                           n_1663, QN => n20422);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => n6693, CK => CLK, Q => 
                           n_1664, QN => n20423);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => n6692, CK => CLK, Q => 
                           n_1665, QN => n20424);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => n6691, CK => CLK, Q => 
                           n_1666, QN => n20425);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => n6690, CK => CLK, Q => 
                           n_1667, QN => n20426);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => n6689, CK => CLK, Q => 
                           n_1668, QN => n20427);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => n6688, CK => CLK, Q => 
                           n_1669, QN => n20428);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => n6687, CK => CLK, Q => 
                           n_1670, QN => n20429);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n6686, CK => CLK, Q => 
                           n_1671, QN => n20430);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n6685, CK => CLK, Q => 
                           n_1672, QN => n20431);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n6684, CK => CLK, Q => 
                           n_1673, QN => n20432);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n6683, CK => CLK, Q => 
                           n_1674, QN => n20433);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n6682, CK => CLK, Q => 
                           n_1675, QN => n20434);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n6681, CK => CLK, Q => 
                           n_1676, QN => n20435);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n6680, CK => CLK, Q => 
                           n_1677, QN => n20436);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n6679, CK => CLK, Q => 
                           n_1678, QN => n20437);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n6678, CK => CLK, Q => 
                           n_1679, QN => n20438);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n6677, CK => CLK, Q => 
                           n_1680, QN => n20439);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n6676, CK => CLK, Q => 
                           n_1681, QN => n20440);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n6675, CK => CLK, Q => 
                           n_1682, QN => n20441);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n6674, CK => CLK, Q => 
                           n_1683, QN => n20442);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n6673, CK => CLK, Q => 
                           n_1684, QN => n20443);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n6672, CK => CLK, Q => 
                           n_1685, QN => n20444);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n6671, CK => CLK, Q => 
                           n_1686, QN => n20445);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n6670, CK => CLK, Q => 
                           n_1687, QN => n20446);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n6669, CK => CLK, Q => 
                           n_1688, QN => n20447);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n6668, CK => CLK, Q => 
                           n_1689, QN => n20448);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n6667, CK => CLK, Q => 
                           n_1690, QN => n20449);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n6666, CK => CLK, Q => 
                           n_1691, QN => n20450);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n6665, CK => CLK, Q => 
                           n_1692, QN => n20451);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n6664, CK => CLK, Q => 
                           n_1693, QN => n20452);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n6663, CK => CLK, Q => 
                           n_1694, QN => n20453);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n6662, CK => CLK, Q => 
                           n_1695, QN => n20454);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n6661, CK => CLK, Q => 
                           n_1696, QN => n20455);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n6660, CK => CLK, Q => 
                           n_1697, QN => n20456);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n6659, CK => CLK, Q => 
                           n_1698, QN => n20457);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n6658, CK => CLK, Q => 
                           n_1699, QN => n20458);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n6657, CK => CLK, Q => 
                           n_1700, QN => n20459);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n6656, CK => CLK, Q => 
                           n_1701, QN => n20460);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n6655, CK => CLK, Q => 
                           n_1702, QN => n20461);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => n5630, CK => CLK, Q => 
                           n_1703, QN => n21094);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => n5629, CK => CLK, Q => 
                           n_1704, QN => n21095);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => n5628, CK => CLK, Q => 
                           n_1705, QN => n21096);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => n5627, CK => CLK, Q => 
                           n_1706, QN => n21097);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => n5822, CK => CLK, Q => 
                           n_1707, QN => n21098);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => n5821, CK => CLK, Q => 
                           n_1708, QN => n21099);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => n5820, CK => CLK, Q => 
                           n_1709, QN => n21100);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => n5819, CK => CLK, Q => 
                           n_1710, QN => n21101);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => n5626, CK => CLK, Q => 
                           n_1711, QN => n21102);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => n5625, CK => CLK, Q => 
                           n_1712, QN => n21103);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => n5624, CK => CLK, Q => 
                           n_1713, QN => n21104);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => n5623, CK => CLK, Q => 
                           n_1714, QN => n21105);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => n5622, CK => CLK, Q => 
                           n_1715, QN => n21106);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => n5621, CK => CLK, Q => 
                           n_1716, QN => n21107);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => n5620, CK => CLK, Q => 
                           n_1717, QN => n21108);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => n5619, CK => CLK, Q => 
                           n_1718, QN => n21109);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => n5618, CK => CLK, Q => 
                           n_1719, QN => n21110);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => n5617, CK => CLK, Q => 
                           n_1720, QN => n21111);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => n5616, CK => CLK, Q => 
                           n_1721, QN => n21112);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => n5615, CK => CLK, Q => 
                           n_1722, QN => n21113);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => n5614, CK => CLK, Q => 
                           n_1723, QN => n21114);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => n5613, CK => CLK, Q => 
                           n_1724, QN => n21115);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => n5612, CK => CLK, Q => 
                           n_1725, QN => n21116);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => n5611, CK => CLK, Q => 
                           n_1726, QN => n21117);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => n5610, CK => CLK, Q => 
                           n_1727, QN => n21118);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => n5609, CK => CLK, Q => 
                           n_1728, QN => n21119);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => n5608, CK => CLK, Q => 
                           n_1729, QN => n21120);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => n5607, CK => CLK, Q => 
                           n_1730, QN => n21121);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => n5606, CK => CLK, Q => 
                           n_1731, QN => n21122);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => n5605, CK => CLK, Q => 
                           n_1732, QN => n21123);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => n5604, CK => CLK, Q => 
                           n_1733, QN => n21124);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => n5603, CK => CLK, Q => 
                           n_1734, QN => n21125);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => n5602, CK => CLK, Q => 
                           n_1735, QN => n21126);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => n5601, CK => CLK, Q => 
                           n_1736, QN => n21127);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => n5600, CK => CLK, Q => 
                           n_1737, QN => n21128);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => n5599, CK => CLK, Q => 
                           n_1738, QN => n21129);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n5598, CK => CLK, Q => 
                           n_1739, QN => n21130);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n5597, CK => CLK, Q => 
                           n_1740, QN => n21131);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n5596, CK => CLK, Q => 
                           n_1741, QN => n21132);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n5595, CK => CLK, Q => 
                           n_1742, QN => n21133);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n5594, CK => CLK, Q => 
                           n_1743, QN => n21134);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n5593, CK => CLK, Q => 
                           n_1744, QN => n21135);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n5592, CK => CLK, Q => 
                           n_1745, QN => n21136);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n5591, CK => CLK, Q => 
                           n_1746, QN => n21137);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n5590, CK => CLK, Q => 
                           n_1747, QN => n21138);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n5589, CK => CLK, Q => 
                           n_1748, QN => n21139);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n5588, CK => CLK, Q => 
                           n_1749, QN => n21140);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n5587, CK => CLK, Q => 
                           n_1750, QN => n21141);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n5586, CK => CLK, Q => 
                           n_1751, QN => n21142);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n5585, CK => CLK, Q => 
                           n_1752, QN => n21143);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n5584, CK => CLK, Q => 
                           n_1753, QN => n21144);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n5583, CK => CLK, Q => 
                           n_1754, QN => n21145);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n5582, CK => CLK, Q => 
                           n_1755, QN => n21146);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n5581, CK => CLK, Q => 
                           n_1756, QN => n21147);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n5580, CK => CLK, Q => 
                           n_1757, QN => n21148);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n5579, CK => CLK, Q => 
                           n_1758, QN => n21149);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n5578, CK => CLK, Q => 
                           n_1759, QN => n21150);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n5577, CK => CLK, Q => 
                           n_1760, QN => n21151);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n5576, CK => CLK, Q => 
                           n_1761, QN => n21152);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n5575, CK => CLK, Q => 
                           n_1762, QN => n21153);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n5574, CK => CLK, Q => 
                           n_1763, QN => n21154);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n5573, CK => CLK, Q => 
                           n_1764, QN => n21155);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n5572, CK => CLK, Q => 
                           n_1765, QN => n21156);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n5571, CK => CLK, Q => 
                           n_1766, QN => n21157);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n5570, CK => CLK, Q => 
                           n_1767, QN => n21158);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n5569, CK => CLK, Q => 
                           n_1768, QN => n21159);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n5568, CK => CLK, Q => 
                           n_1769, QN => n21160);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n5567, CK => CLK, Q => 
                           n_1770, QN => n21161);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => n5818, CK => CLK, Q => 
                           n_1771, QN => n21162);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => n5817, CK => CLK, Q => 
                           n_1772, QN => n21163);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => n5816, CK => CLK, Q => 
                           n_1773, QN => n21164);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => n5815, CK => CLK, Q => 
                           n_1774, QN => n21165);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => n5814, CK => CLK, Q => 
                           n_1775, QN => n21166);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => n5813, CK => CLK, Q => 
                           n_1776, QN => n21167);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => n5812, CK => CLK, Q => 
                           n_1777, QN => n21168);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => n5811, CK => CLK, Q => 
                           n_1778, QN => n21169);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => n5810, CK => CLK, Q => 
                           n_1779, QN => n21170);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => n5809, CK => CLK, Q => 
                           n_1780, QN => n21171);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => n5808, CK => CLK, Q => 
                           n_1781, QN => n21172);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => n5807, CK => CLK, Q => 
                           n_1782, QN => n21173);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => n5806, CK => CLK, Q => 
                           n_1783, QN => n21174);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => n5805, CK => CLK, Q => 
                           n_1784, QN => n21175);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => n5804, CK => CLK, Q => 
                           n_1785, QN => n21176);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => n5803, CK => CLK, Q => 
                           n_1786, QN => n21177);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => n5802, CK => CLK, Q => 
                           n_1787, QN => n21178);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => n5801, CK => CLK, Q => 
                           n_1788, QN => n21179);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => n5800, CK => CLK, Q => 
                           n_1789, QN => n21180);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => n5799, CK => CLK, Q => 
                           n_1790, QN => n21181);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => n5798, CK => CLK, Q => 
                           n_1791, QN => n21182);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => n5797, CK => CLK, Q => 
                           n_1792, QN => n21183);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => n5796, CK => CLK, Q => 
                           n_1793, QN => n21184);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => n5795, CK => CLK, Q => 
                           n_1794, QN => n21185);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => n5794, CK => CLK, Q => 
                           n_1795, QN => n21186);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => n5793, CK => CLK, Q => 
                           n_1796, QN => n21187);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => n5792, CK => CLK, Q => 
                           n_1797, QN => n21188);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => n5791, CK => CLK, Q => 
                           n_1798, QN => n21189);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n5790, CK => CLK, Q => 
                           n_1799, QN => n21190);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n5789, CK => CLK, Q => 
                           n_1800, QN => n21191);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n5788, CK => CLK, Q => 
                           n_1801, QN => n21192);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n5787, CK => CLK, Q => 
                           n_1802, QN => n21193);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n5786, CK => CLK, Q => 
                           n_1803, QN => n21194);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n5785, CK => CLK, Q => 
                           n_1804, QN => n21195);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n5784, CK => CLK, Q => 
                           n_1805, QN => n21196);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n5783, CK => CLK, Q => 
                           n_1806, QN => n21197);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n5782, CK => CLK, Q => 
                           n_1807, QN => n21198);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n5781, CK => CLK, Q => 
                           n_1808, QN => n21199);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n5780, CK => CLK, Q => 
                           n_1809, QN => n21200);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n5779, CK => CLK, Q => 
                           n_1810, QN => n21201);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n5778, CK => CLK, Q => 
                           n_1811, QN => n21202);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n5777, CK => CLK, Q => 
                           n_1812, QN => n21203);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n5776, CK => CLK, Q => 
                           n_1813, QN => n21204);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n5775, CK => CLK, Q => 
                           n_1814, QN => n21205);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n5774, CK => CLK, Q => 
                           n_1815, QN => n21206);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n5773, CK => CLK, Q => 
                           n_1816, QN => n21207);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n5772, CK => CLK, Q => 
                           n_1817, QN => n21208);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n5771, CK => CLK, Q => 
                           n_1818, QN => n21209);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n5770, CK => CLK, Q => 
                           n_1819, QN => n21210);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n5769, CK => CLK, Q => 
                           n_1820, QN => n21211);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n5768, CK => CLK, Q => 
                           n_1821, QN => n21212);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n5767, CK => CLK, Q => 
                           n_1822, QN => n21213);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n5766, CK => CLK, Q => 
                           n_1823, QN => n21214);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n5765, CK => CLK, Q => 
                           n_1824, QN => n21215);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n5764, CK => CLK, Q => 
                           n_1825, QN => n21216);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n5763, CK => CLK, Q => 
                           n_1826, QN => n21217);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n5762, CK => CLK, Q => 
                           n_1827, QN => n21218);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n5761, CK => CLK, Q => 
                           n_1828, QN => n21219);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n5760, CK => CLK, Q => 
                           n_1829, QN => n21220);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n5759, CK => CLK, Q => 
                           n_1830, QN => n21221);
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => n6782, CK => CLK, Q => 
                           n_1831, QN => n21222);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => n6781, CK => CLK, Q => 
                           n_1832, QN => n21223);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => n6780, CK => CLK, Q => 
                           n_1833, QN => n21224);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => n6779, CK => CLK, Q => 
                           n_1834, QN => n21225);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => n6778, CK => CLK, Q => 
                           n_1835, QN => n21226);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => n6777, CK => CLK, Q => 
                           n_1836, QN => n21227);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => n6776, CK => CLK, Q => 
                           n_1837, QN => n21228);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => n6775, CK => CLK, Q => 
                           n_1838, QN => n21229);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => n6774, CK => CLK, Q => 
                           n_1839, QN => n21230);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => n6773, CK => CLK, Q => 
                           n_1840, QN => n21231);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => n6772, CK => CLK, Q => 
                           n_1841, QN => n21232);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => n6771, CK => CLK, Q => 
                           n_1842, QN => n21233);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => n6770, CK => CLK, Q => 
                           n_1843, QN => n21234);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => n6769, CK => CLK, Q => 
                           n_1844, QN => n21235);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => n6768, CK => CLK, Q => 
                           n_1845, QN => n21236);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => n6767, CK => CLK, Q => 
                           n_1846, QN => n21237);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => n6766, CK => CLK, Q => 
                           n_1847, QN => n21238);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => n6765, CK => CLK, Q => 
                           n_1848, QN => n21239);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => n6764, CK => CLK, Q => 
                           n_1849, QN => n21240);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => n6763, CK => CLK, Q => 
                           n_1850, QN => n21241);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => n6762, CK => CLK, Q => 
                           n_1851, QN => n21242);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => n6761, CK => CLK, Q => 
                           n_1852, QN => n21243);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => n6760, CK => CLK, Q => 
                           n_1853, QN => n21244);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => n6759, CK => CLK, Q => 
                           n_1854, QN => n21245);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => n6758, CK => CLK, Q => 
                           n_1855, QN => n21246);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => n6757, CK => CLK, Q => 
                           n_1856, QN => n21247);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => n6756, CK => CLK, Q => 
                           n_1857, QN => n21248);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => n6755, CK => CLK, Q => 
                           n_1858, QN => n21249);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => n6754, CK => CLK, Q => 
                           n_1859, QN => n21250);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => n6753, CK => CLK, Q => 
                           n_1860, QN => n21251);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => n6752, CK => CLK, Q => 
                           n_1861, QN => n21252);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => n6751, CK => CLK, Q => 
                           n_1862, QN => n21253);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n6750, CK => CLK, Q => 
                           n_1863, QN => n21254);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n6749, CK => CLK, Q => 
                           n_1864, QN => n21255);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n6748, CK => CLK, Q => 
                           n_1865, QN => n21256);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n6747, CK => CLK, Q => 
                           n_1866, QN => n21257);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n6746, CK => CLK, Q => 
                           n_1867, QN => n21258);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n6745, CK => CLK, Q => 
                           n_1868, QN => n21259);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n6744, CK => CLK, Q => 
                           n_1869, QN => n21260);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n6743, CK => CLK, Q => 
                           n_1870, QN => n21261);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n6742, CK => CLK, Q => 
                           n_1871, QN => n21262);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n6741, CK => CLK, Q => 
                           n_1872, QN => n21263);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n6740, CK => CLK, Q => 
                           n_1873, QN => n21264);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n6739, CK => CLK, Q => 
                           n_1874, QN => n21265);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n6738, CK => CLK, Q => 
                           n_1875, QN => n21266);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n6737, CK => CLK, Q => 
                           n_1876, QN => n21267);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n6736, CK => CLK, Q => 
                           n_1877, QN => n21268);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n6735, CK => CLK, Q => 
                           n_1878, QN => n21269);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n6734, CK => CLK, Q => 
                           n_1879, QN => n21270);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n6733, CK => CLK, Q => 
                           n_1880, QN => n21271);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n6732, CK => CLK, Q => 
                           n_1881, QN => n21272);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n6731, CK => CLK, Q => 
                           n_1882, QN => n21273);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n6730, CK => CLK, Q => 
                           n_1883, QN => n21274);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n6729, CK => CLK, Q => 
                           n_1884, QN => n21275);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n6728, CK => CLK, Q => 
                           n_1885, QN => n21276);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n6727, CK => CLK, Q => 
                           n_1886, QN => n21277);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n6726, CK => CLK, Q => 
                           n_1887, QN => n21278);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n6725, CK => CLK, Q => 
                           n_1888, QN => n21279);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n6724, CK => CLK, Q => 
                           n_1889, QN => n21280);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n6723, CK => CLK, Q => 
                           n_1890, QN => n21281);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n6722, CK => CLK, Q => 
                           n_1891, QN => n21282);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n6721, CK => CLK, Q => 
                           n_1892, QN => n21283);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n6720, CK => CLK, Q => 
                           n_1893, QN => n21284);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n6719, CK => CLK, Q => 
                           n_1894, QN => n21285);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => n6910, CK => CLK, Q => 
                           n_1895, QN => n20133);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => n6909, CK => CLK, Q => 
                           n_1896, QN => n19750);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => n6908, CK => CLK, Q => 
                           n_1897, QN => n19751);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => n6907, CK => CLK, Q => 
                           n_1898, QN => n19752);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => n6906, CK => CLK, Q => 
                           n_1899, QN => n19753);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => n6905, CK => CLK, Q => 
                           n_1900, QN => n19754);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => n6904, CK => CLK, Q => 
                           n_1901, QN => n19755);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => n6903, CK => CLK, Q => 
                           n_1902, QN => n19756);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => n6902, CK => CLK, Q => 
                           n_1903, QN => n19757);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => n6901, CK => CLK, Q => 
                           n_1904, QN => n19758);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => n6900, CK => CLK, Q => 
                           n_1905, QN => n19759);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => n6899, CK => CLK, Q => 
                           n_1906, QN => n19760);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => n6898, CK => CLK, Q => 
                           n_1907, QN => n19761);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => n6897, CK => CLK, Q => 
                           n_1908, QN => n19762);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => n6896, CK => CLK, Q => 
                           n_1909, QN => n19763);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => n6895, CK => CLK, Q => 
                           n_1910, QN => n19764);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => n6894, CK => CLK, Q => 
                           n_1911, QN => n19765);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => n6893, CK => CLK, Q => 
                           n_1912, QN => n19766);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => n6892, CK => CLK, Q => 
                           n_1913, QN => n19767);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => n6891, CK => CLK, Q => 
                           n_1914, QN => n19768);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => n6890, CK => CLK, Q => 
                           n_1915, QN => n19769);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => n6889, CK => CLK, Q => 
                           n_1916, QN => n19770);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => n6888, CK => CLK, Q => 
                           n_1917, QN => n19771);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => n6887, CK => CLK, Q => 
                           n_1918, QN => n19772);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => n6886, CK => CLK, Q => 
                           n_1919, QN => n19773);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => n6885, CK => CLK, Q => 
                           n_1920, QN => n19774);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => n6884, CK => CLK, Q => 
                           n_1921, QN => n19775);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => n6883, CK => CLK, Q => 
                           n_1922, QN => n19776);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => n6882, CK => CLK, Q => 
                           n_1923, QN => n19777);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => n6881, CK => CLK, Q => 
                           n_1924, QN => n19778);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => n6880, CK => CLK, Q => 
                           n_1925, QN => n19779);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => n6879, CK => CLK, Q => 
                           n_1926, QN => n19780);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n6878, CK => CLK, Q => 
                           n_1927, QN => n19781);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n6877, CK => CLK, Q => 
                           n_1928, QN => n19782);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n6876, CK => CLK, Q => 
                           n_1929, QN => n19783);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n6875, CK => CLK, Q => 
                           n_1930, QN => n19784);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n6874, CK => CLK, Q => 
                           n_1931, QN => n19785);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n6873, CK => CLK, Q => 
                           n_1932, QN => n19786);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n6872, CK => CLK, Q => 
                           n_1933, QN => n19787);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n6871, CK => CLK, Q => 
                           n_1934, QN => n19788);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n6870, CK => CLK, Q => 
                           n_1935, QN => n19789);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n6869, CK => CLK, Q => 
                           n_1936, QN => n19790);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n6868, CK => CLK, Q => 
                           n_1937, QN => n19791);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n6867, CK => CLK, Q => 
                           n_1938, QN => n19792);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n6866, CK => CLK, Q => 
                           n_1939, QN => n19793);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n6865, CK => CLK, Q => 
                           n_1940, QN => n19794);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n6864, CK => CLK, Q => 
                           n_1941, QN => n19795);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n6863, CK => CLK, Q => 
                           n_1942, QN => n19796);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n6862, CK => CLK, Q => 
                           n_1943, QN => n19797);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n6861, CK => CLK, Q => 
                           n_1944, QN => n19798);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n6860, CK => CLK, Q => 
                           n_1945, QN => n19799);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n6859, CK => CLK, Q => 
                           n_1946, QN => n19800);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n6858, CK => CLK, Q => 
                           n_1947, QN => n19801);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n6857, CK => CLK, Q => 
                           n_1948, QN => n19802);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n6856, CK => CLK, Q => n_1949
                           , QN => n19803);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n6855, CK => CLK, Q => n_1950
                           , QN => n19804);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n6854, CK => CLK, Q => n_1951
                           , QN => n19805);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n6853, CK => CLK, Q => n_1952
                           , QN => n19806);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n6852, CK => CLK, Q => n_1953
                           , QN => n19807);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n6851, CK => CLK, Q => n_1954
                           , QN => n19808);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n6850, CK => CLK, Q => n_1955
                           , QN => n19809);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n6849, CK => CLK, Q => n_1956
                           , QN => n19810);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n6848, CK => CLK, Q => n_1957
                           , QN => n19811);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n6847, CK => CLK, Q => n_1958
                           , QN => n19812);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => n7230, CK => CLK, Q => 
                           n_1959, QN => n20646);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => n7229, CK => CLK, Q => 
                           n_1960, QN => n20647);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => n7228, CK => CLK, Q => 
                           n_1961, QN => n20648);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => n7227, CK => CLK, Q => 
                           n_1962, QN => n20649);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => n7226, CK => CLK, Q => 
                           n_1963, QN => n20650);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => n7225, CK => CLK, Q => 
                           n_1964, QN => n20651);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => n7224, CK => CLK, Q => 
                           n_1965, QN => n20652);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => n7223, CK => CLK, Q => 
                           n_1966, QN => n20653);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => n7222, CK => CLK, Q => 
                           n_1967, QN => n20654);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => n7221, CK => CLK, Q => 
                           n_1968, QN => n20655);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => n7220, CK => CLK, Q => 
                           n_1969, QN => n20656);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => n7219, CK => CLK, Q => 
                           n_1970, QN => n20657);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => n7218, CK => CLK, Q => 
                           n_1971, QN => n20658);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => n7217, CK => CLK, Q => 
                           n_1972, QN => n20659);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => n7216, CK => CLK, Q => 
                           n_1973, QN => n20660);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => n7215, CK => CLK, Q => 
                           n_1974, QN => n20661);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => n7214, CK => CLK, Q => 
                           n_1975, QN => n20662);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => n7213, CK => CLK, Q => 
                           n_1976, QN => n20663);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => n7212, CK => CLK, Q => 
                           n_1977, QN => n20664);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => n7211, CK => CLK, Q => 
                           n_1978, QN => n20665);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => n7210, CK => CLK, Q => 
                           n_1979, QN => n20666);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => n7209, CK => CLK, Q => 
                           n_1980, QN => n20667);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => n7208, CK => CLK, Q => 
                           n_1981, QN => n20668);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => n7207, CK => CLK, Q => 
                           n_1982, QN => n20669);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => n7206, CK => CLK, Q => 
                           n_1983, QN => n20670);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => n7205, CK => CLK, Q => 
                           n_1984, QN => n20671);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => n7204, CK => CLK, Q => 
                           n_1985, QN => n20672);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => n7203, CK => CLK, Q => 
                           n_1986, QN => n20673);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => n7202, CK => CLK, Q => 
                           n_1987, QN => n20674);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => n7201, CK => CLK, Q => 
                           n_1988, QN => n20675);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => n7200, CK => CLK, Q => 
                           n_1989, QN => n20676);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => n7199, CK => CLK, Q => 
                           n_1990, QN => n20677);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n7198, CK => CLK, Q => 
                           n_1991, QN => n20678);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n7197, CK => CLK, Q => 
                           n_1992, QN => n20679);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n7196, CK => CLK, Q => 
                           n_1993, QN => n20680);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n7195, CK => CLK, Q => 
                           n_1994, QN => n20681);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n7194, CK => CLK, Q => 
                           n_1995, QN => n20682);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n7193, CK => CLK, Q => 
                           n_1996, QN => n20683);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n7192, CK => CLK, Q => 
                           n_1997, QN => n20684);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n7191, CK => CLK, Q => 
                           n_1998, QN => n20685);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n7190, CK => CLK, Q => 
                           n_1999, QN => n20686);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n7189, CK => CLK, Q => 
                           n_2000, QN => n20687);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n7188, CK => CLK, Q => 
                           n_2001, QN => n20688);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n7187, CK => CLK, Q => 
                           n_2002, QN => n20689);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n7186, CK => CLK, Q => 
                           n_2003, QN => n20690);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n7185, CK => CLK, Q => 
                           n_2004, QN => n20691);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n7184, CK => CLK, Q => 
                           n_2005, QN => n20692);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n7183, CK => CLK, Q => 
                           n_2006, QN => n20693);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n7182, CK => CLK, Q => 
                           n_2007, QN => n20694);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n7181, CK => CLK, Q => 
                           n_2008, QN => n20695);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n7180, CK => CLK, Q => 
                           n_2009, QN => n20696);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n7179, CK => CLK, Q => 
                           n_2010, QN => n20697);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n7178, CK => CLK, Q => 
                           n_2011, QN => n20698);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n7177, CK => CLK, Q => 
                           n_2012, QN => n20699);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n7176, CK => CLK, Q => n_2013
                           , QN => n20700);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n7175, CK => CLK, Q => n_2014
                           , QN => n20701);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n7174, CK => CLK, Q => n_2015
                           , QN => n20702);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n7173, CK => CLK, Q => n_2016
                           , QN => n20703);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n7172, CK => CLK, Q => n_2017
                           , QN => n20704);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n7171, CK => CLK, Q => n_2018
                           , QN => n20705);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n7170, CK => CLK, Q => n_2019
                           , QN => n20706);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n7169, CK => CLK, Q => n_2020
                           , QN => n20707);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n7168, CK => CLK, Q => n_2021
                           , QN => n20708);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n7167, CK => CLK, Q => n_2022
                           , QN => n20709);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => n6270, CK => CLK, Q => 
                           n_2023, QN => n20710);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => n6269, CK => CLK, Q => 
                           n_2024, QN => n20711);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => n6268, CK => CLK, Q => 
                           n_2025, QN => n20712);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => n6267, CK => CLK, Q => 
                           n_2026, QN => n20713);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => n6266, CK => CLK, Q => 
                           n_2027, QN => n20714);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => n6265, CK => CLK, Q => 
                           n_2028, QN => n20715);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => n6264, CK => CLK, Q => 
                           n_2029, QN => n20716);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => n6263, CK => CLK, Q => 
                           n_2030, QN => n20717);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => n6262, CK => CLK, Q => 
                           n_2031, QN => n20718);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => n6261, CK => CLK, Q => 
                           n_2032, QN => n20719);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => n6260, CK => CLK, Q => 
                           n_2033, QN => n20720);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => n6259, CK => CLK, Q => 
                           n_2034, QN => n20721);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => n6258, CK => CLK, Q => 
                           n_2035, QN => n20722);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => n6257, CK => CLK, Q => 
                           n_2036, QN => n20723);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => n6256, CK => CLK, Q => 
                           n_2037, QN => n20724);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => n6255, CK => CLK, Q => 
                           n_2038, QN => n20725);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => n6254, CK => CLK, Q => 
                           n_2039, QN => n20726);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => n6253, CK => CLK, Q => 
                           n_2040, QN => n20727);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => n6252, CK => CLK, Q => 
                           n_2041, QN => n20728);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => n6251, CK => CLK, Q => 
                           n_2042, QN => n20729);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => n6250, CK => CLK, Q => 
                           n_2043, QN => n20730);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => n6249, CK => CLK, Q => 
                           n_2044, QN => n20731);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => n6248, CK => CLK, Q => 
                           n_2045, QN => n20732);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => n6247, CK => CLK, Q => 
                           n_2046, QN => n20733);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => n6246, CK => CLK, Q => 
                           n_2047, QN => n20734);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => n6245, CK => CLK, Q => 
                           n_2048, QN => n20735);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => n6244, CK => CLK, Q => 
                           n_2049, QN => n20736);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => n6243, CK => CLK, Q => 
                           n_2050, QN => n20737);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => n6242, CK => CLK, Q => 
                           n_2051, QN => n20738);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => n6241, CK => CLK, Q => 
                           n_2052, QN => n20739);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => n6240, CK => CLK, Q => 
                           n_2053, QN => n20740);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => n6239, CK => CLK, Q => 
                           n_2054, QN => n20741);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n6238, CK => CLK, Q => 
                           n_2055, QN => n20742);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n6237, CK => CLK, Q => 
                           n_2056, QN => n20743);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n6236, CK => CLK, Q => 
                           n_2057, QN => n20744);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n6235, CK => CLK, Q => 
                           n_2058, QN => n20745);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n6234, CK => CLK, Q => 
                           n_2059, QN => n20746);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n6233, CK => CLK, Q => 
                           n_2060, QN => n20747);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n6232, CK => CLK, Q => 
                           n_2061, QN => n20748);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n6231, CK => CLK, Q => 
                           n_2062, QN => n20749);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n6230, CK => CLK, Q => 
                           n_2063, QN => n20750);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n6229, CK => CLK, Q => 
                           n_2064, QN => n20751);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n6228, CK => CLK, Q => 
                           n_2065, QN => n20752);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n6227, CK => CLK, Q => 
                           n_2066, QN => n20753);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n6226, CK => CLK, Q => 
                           n_2067, QN => n20754);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n6225, CK => CLK, Q => 
                           n_2068, QN => n20755);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n6224, CK => CLK, Q => 
                           n_2069, QN => n20756);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n6223, CK => CLK, Q => 
                           n_2070, QN => n20757);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n6222, CK => CLK, Q => 
                           n_2071, QN => n20758);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n6221, CK => CLK, Q => 
                           n_2072, QN => n20759);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n6220, CK => CLK, Q => 
                           n_2073, QN => n20760);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n6219, CK => CLK, Q => 
                           n_2074, QN => n20761);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n6218, CK => CLK, Q => 
                           n_2075, QN => n20762);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n6217, CK => CLK, Q => 
                           n_2076, QN => n20763);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n6216, CK => CLK, Q => 
                           n_2077, QN => n20764);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n6215, CK => CLK, Q => 
                           n_2078, QN => n20765);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n6214, CK => CLK, Q => 
                           n_2079, QN => n20766);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n6213, CK => CLK, Q => 
                           n_2080, QN => n20767);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n6212, CK => CLK, Q => 
                           n_2081, QN => n20768);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n6211, CK => CLK, Q => 
                           n_2082, QN => n20769);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n6210, CK => CLK, Q => 
                           n_2083, QN => n20770);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n6209, CK => CLK, Q => 
                           n_2084, QN => n20771);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n6208, CK => CLK, Q => 
                           n_2085, QN => n20772);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n6207, CK => CLK, Q => 
                           n_2086, QN => n20773);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => n6398, CK => CLK, Q => 
                           n_2087, QN => n21350);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => n6397, CK => CLK, Q => 
                           n_2088, QN => n21351);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => n6396, CK => CLK, Q => 
                           n_2089, QN => n21352);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => n6395, CK => CLK, Q => 
                           n_2090, QN => n21353);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => n6394, CK => CLK, Q => 
                           n_2091, QN => n21354);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => n6393, CK => CLK, Q => 
                           n_2092, QN => n21355);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => n6392, CK => CLK, Q => 
                           n_2093, QN => n21356);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => n6391, CK => CLK, Q => 
                           n_2094, QN => n21357);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => n6390, CK => CLK, Q => 
                           n_2095, QN => n21358);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => n6389, CK => CLK, Q => 
                           n_2096, QN => n21359);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => n6388, CK => CLK, Q => 
                           n_2097, QN => n21360);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => n6387, CK => CLK, Q => 
                           n_2098, QN => n21361);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => n6386, CK => CLK, Q => 
                           n_2099, QN => n21362);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => n6385, CK => CLK, Q => 
                           n_2100, QN => n21363);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => n6384, CK => CLK, Q => 
                           n_2101, QN => n21364);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => n6383, CK => CLK, Q => 
                           n_2102, QN => n21365);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => n6382, CK => CLK, Q => 
                           n_2103, QN => n21366);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => n6381, CK => CLK, Q => 
                           n_2104, QN => n21367);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => n6380, CK => CLK, Q => 
                           n_2105, QN => n21368);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => n6379, CK => CLK, Q => 
                           n_2106, QN => n21369);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => n6378, CK => CLK, Q => 
                           n_2107, QN => n21370);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => n6377, CK => CLK, Q => 
                           n_2108, QN => n21371);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => n6376, CK => CLK, Q => 
                           n_2109, QN => n21372);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => n6375, CK => CLK, Q => 
                           n_2110, QN => n21373);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => n6374, CK => CLK, Q => 
                           n_2111, QN => n21374);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => n6373, CK => CLK, Q => 
                           n_2112, QN => n21375);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => n6372, CK => CLK, Q => 
                           n_2113, QN => n21376);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => n6371, CK => CLK, Q => 
                           n_2114, QN => n21377);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => n6370, CK => CLK, Q => 
                           n_2115, QN => n21378);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => n6369, CK => CLK, Q => 
                           n_2116, QN => n21379);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => n6368, CK => CLK, Q => 
                           n_2117, QN => n21380);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => n6367, CK => CLK, Q => 
                           n_2118, QN => n21381);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n6366, CK => CLK, Q => 
                           n_2119, QN => n21382);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n6365, CK => CLK, Q => 
                           n_2120, QN => n21383);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n6364, CK => CLK, Q => 
                           n_2121, QN => n21384);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n6363, CK => CLK, Q => 
                           n_2122, QN => n21385);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n6362, CK => CLK, Q => 
                           n_2123, QN => n21386);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n6361, CK => CLK, Q => 
                           n_2124, QN => n21387);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n6360, CK => CLK, Q => 
                           n_2125, QN => n21388);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n6359, CK => CLK, Q => 
                           n_2126, QN => n21389);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n6358, CK => CLK, Q => 
                           n_2127, QN => n21390);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n6357, CK => CLK, Q => 
                           n_2128, QN => n21391);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n6356, CK => CLK, Q => 
                           n_2129, QN => n21392);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n6355, CK => CLK, Q => 
                           n_2130, QN => n21393);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n6354, CK => CLK, Q => 
                           n_2131, QN => n21394);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n6353, CK => CLK, Q => 
                           n_2132, QN => n21395);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n6352, CK => CLK, Q => 
                           n_2133, QN => n21396);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n6351, CK => CLK, Q => 
                           n_2134, QN => n21397);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n6350, CK => CLK, Q => 
                           n_2135, QN => n21398);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n6349, CK => CLK, Q => 
                           n_2136, QN => n21399);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n6348, CK => CLK, Q => 
                           n_2137, QN => n21400);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n6347, CK => CLK, Q => 
                           n_2138, QN => n21401);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n6346, CK => CLK, Q => 
                           n_2139, QN => n21402);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n6345, CK => CLK, Q => 
                           n_2140, QN => n21403);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n6344, CK => CLK, Q => 
                           n_2141, QN => n21404);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n6343, CK => CLK, Q => 
                           n_2142, QN => n21405);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n6342, CK => CLK, Q => 
                           n_2143, QN => n21406);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n6341, CK => CLK, Q => 
                           n_2144, QN => n21407);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n6340, CK => CLK, Q => 
                           n_2145, QN => n21408);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n6339, CK => CLK, Q => 
                           n_2146, QN => n21409);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n6338, CK => CLK, Q => 
                           n_2147, QN => n21410);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n6337, CK => CLK, Q => 
                           n_2148, QN => n21411);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n6336, CK => CLK, Q => 
                           n_2149, QN => n21412);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n6335, CK => CLK, Q => 
                           n_2150, QN => n21413);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => n5502, CK => CLK, Q => 
                           n17163, QN => n20774);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => n5501, CK => CLK, Q => 
                           n17184, QN => n20775);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => n5500, CK => CLK, Q => 
                           n17205, QN => n20776);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => n5499, CK => CLK, Q => 
                           n17226, QN => n20777);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => n5886, CK => CLK, Q => 
                           n17161, QN => n20778);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => n5885, CK => CLK, Q => 
                           n17182, QN => n20779);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => n5884, CK => CLK, Q => 
                           n17203, QN => n20780);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => n5883, CK => CLK, Q => 
                           n17224, QN => n20781);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => n5498, CK => CLK, Q => 
                           n17247, QN => n20782);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => n5497, CK => CLK, Q => 
                           n17268, QN => n20783);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => n5496, CK => CLK, Q => 
                           n17289, QN => n20784);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => n5495, CK => CLK, Q => 
                           n17310, QN => n20785);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => n5494, CK => CLK, Q => 
                           n17331, QN => n20786);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => n5493, CK => CLK, Q => 
                           n17352, QN => n20787);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => n5492, CK => CLK, Q => 
                           n17373, QN => n20788);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => n5491, CK => CLK, Q => 
                           n17394, QN => n20789);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => n5490, CK => CLK, Q => 
                           n17415, QN => n20790);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => n5489, CK => CLK, Q => 
                           n17436, QN => n20791);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => n5488, CK => CLK, Q => 
                           n17457, QN => n20792);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => n5487, CK => CLK, Q => 
                           n17478, QN => n20793);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => n5486, CK => CLK, Q => 
                           n17499, QN => n20794);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => n5485, CK => CLK, Q => 
                           n17520, QN => n20795);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => n5484, CK => CLK, Q => 
                           n17541, QN => n20796);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => n5483, CK => CLK, Q => 
                           n17562, QN => n20797);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => n5482, CK => CLK, Q => 
                           n17583, QN => n20798);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => n5481, CK => CLK, Q => 
                           n17604, QN => n20799);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => n5480, CK => CLK, Q => 
                           n17625, QN => n20800);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => n5479, CK => CLK, Q => 
                           n17646, QN => n20801);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => n5478, CK => CLK, Q => 
                           n17667, QN => n20802);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => n5477, CK => CLK, Q => 
                           n17688, QN => n20803);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => n5476, CK => CLK, Q => 
                           n17709, QN => n20804);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => n5475, CK => CLK, Q => 
                           n17730, QN => n20805);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => n5474, CK => CLK, Q => 
                           n17751, QN => n20806);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => n5473, CK => CLK, Q => 
                           n17772, QN => n20807);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => n5472, CK => CLK, Q => 
                           n17793, QN => n20808);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => n5471, CK => CLK, Q => 
                           n17814, QN => n20809);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n5470, CK => CLK, Q => 
                           n17835, QN => n20810);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n5469, CK => CLK, Q => 
                           n17856, QN => n20811);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n5468, CK => CLK, Q => 
                           n17877, QN => n20812);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n5467, CK => CLK, Q => 
                           n17898, QN => n20813);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n5466, CK => CLK, Q => 
                           n17919, QN => n20814);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n5465, CK => CLK, Q => 
                           n17940, QN => n20815);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n5464, CK => CLK, Q => 
                           n17961, QN => n20816);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n5463, CK => CLK, Q => 
                           n17982, QN => n20817);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n5462, CK => CLK, Q => 
                           n18003, QN => n20818);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n5461, CK => CLK, Q => 
                           n18024, QN => n20819);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n5460, CK => CLK, Q => 
                           n18045, QN => n20820);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n5459, CK => CLK, Q => 
                           n18066, QN => n20821);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n5458, CK => CLK, Q => 
                           n18087, QN => n20822);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n5457, CK => CLK, Q => 
                           n18108, QN => n20823);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n5456, CK => CLK, Q => 
                           n18129, QN => n20824);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n5455, CK => CLK, Q => 
                           n18150, QN => n20825);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n5454, CK => CLK, Q => 
                           n18171, QN => n20826);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n5453, CK => CLK, Q => 
                           n18192, QN => n20827);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n5452, CK => CLK, Q => 
                           n18213, QN => n20828);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n5451, CK => CLK, Q => 
                           n18234, QN => n20829);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n5450, CK => CLK, Q => 
                           n18255, QN => n20830);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n5449, CK => CLK, Q => 
                           n18276, QN => n20831);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n5448, CK => CLK, Q => 
                           n18297, QN => n20832);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n5447, CK => CLK, Q => 
                           n18318, QN => n20833);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n5446, CK => CLK, Q => 
                           n18339, QN => n20834);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n5445, CK => CLK, Q => 
                           n18360, QN => n20835);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n5444, CK => CLK, Q => 
                           n18381, QN => n20836);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n5443, CK => CLK, Q => 
                           n18402, QN => n20837);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n5442, CK => CLK, Q => 
                           n18423, QN => n20838);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n5441, CK => CLK, Q => 
                           n18444, QN => n20839);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n5440, CK => CLK, Q => 
                           n18465, QN => n20840);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n5439, CK => CLK, Q => 
                           n18486, QN => n20841);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => n5882, CK => CLK, Q => 
                           n17245, QN => n20842);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => n5881, CK => CLK, Q => 
                           n17266, QN => n20843);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => n5880, CK => CLK, Q => 
                           n17287, QN => n20844);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => n5879, CK => CLK, Q => 
                           n17308, QN => n20845);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => n5878, CK => CLK, Q => 
                           n17329, QN => n20846);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => n5877, CK => CLK, Q => 
                           n17350, QN => n20847);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => n5876, CK => CLK, Q => 
                           n17371, QN => n20848);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => n5875, CK => CLK, Q => 
                           n17392, QN => n20849);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => n5874, CK => CLK, Q => 
                           n17413, QN => n20850);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => n5873, CK => CLK, Q => 
                           n17434, QN => n20851);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => n5872, CK => CLK, Q => 
                           n17455, QN => n20852);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => n5871, CK => CLK, Q => 
                           n17476, QN => n20853);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => n5870, CK => CLK, Q => 
                           n17497, QN => n20854);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => n5869, CK => CLK, Q => 
                           n17518, QN => n20855);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => n5868, CK => CLK, Q => 
                           n17539, QN => n20856);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => n5867, CK => CLK, Q => 
                           n17560, QN => n20857);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => n5866, CK => CLK, Q => 
                           n17581, QN => n20858);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => n5865, CK => CLK, Q => 
                           n17602, QN => n20859);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => n5864, CK => CLK, Q => 
                           n17623, QN => n20860);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => n5863, CK => CLK, Q => 
                           n17644, QN => n20861);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => n5862, CK => CLK, Q => 
                           n17665, QN => n20862);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => n5861, CK => CLK, Q => 
                           n17686, QN => n20863);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => n5860, CK => CLK, Q => 
                           n17707, QN => n20864);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => n5859, CK => CLK, Q => 
                           n17728, QN => n20865);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => n5858, CK => CLK, Q => 
                           n17749, QN => n20866);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => n5857, CK => CLK, Q => 
                           n17770, QN => n20867);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => n5856, CK => CLK, Q => 
                           n17791, QN => n20868);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => n5855, CK => CLK, Q => 
                           n17812, QN => n20869);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n5854, CK => CLK, Q => 
                           n17833, QN => n20870);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n5853, CK => CLK, Q => 
                           n17854, QN => n20871);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n5852, CK => CLK, Q => 
                           n17875, QN => n20872);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n5851, CK => CLK, Q => 
                           n17896, QN => n20873);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n5850, CK => CLK, Q => 
                           n17917, QN => n20874);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n5849, CK => CLK, Q => 
                           n17938, QN => n20875);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n5848, CK => CLK, Q => 
                           n17959, QN => n20876);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n5847, CK => CLK, Q => 
                           n17980, QN => n20877);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n5846, CK => CLK, Q => 
                           n18001, QN => n20878);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n5845, CK => CLK, Q => 
                           n18022, QN => n20879);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n5844, CK => CLK, Q => 
                           n18043, QN => n20880);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n5843, CK => CLK, Q => 
                           n18064, QN => n20881);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n5842, CK => CLK, Q => 
                           n18085, QN => n20882);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n5841, CK => CLK, Q => 
                           n18106, QN => n20883);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n5840, CK => CLK, Q => 
                           n18127, QN => n20884);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n5839, CK => CLK, Q => 
                           n18148, QN => n20885);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n5838, CK => CLK, Q => 
                           n18169, QN => n20886);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n5837, CK => CLK, Q => 
                           n18190, QN => n20887);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n5836, CK => CLK, Q => 
                           n18211, QN => n20888);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n5835, CK => CLK, Q => 
                           n18232, QN => n20889);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n5834, CK => CLK, Q => 
                           n18253, QN => n20890);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n5833, CK => CLK, Q => 
                           n18274, QN => n20891);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n5832, CK => CLK, Q => 
                           n18295, QN => n20892);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n5831, CK => CLK, Q => 
                           n18316, QN => n20893);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n5830, CK => CLK, Q => 
                           n18337, QN => n20894);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n5829, CK => CLK, Q => 
                           n18358, QN => n20895);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n5828, CK => CLK, Q => 
                           n18379, QN => n20896);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n5827, CK => CLK, Q => 
                           n18400, QN => n20897);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n5826, CK => CLK, Q => 
                           n18421, QN => n20898);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n5825, CK => CLK, Q => 
                           n18442, QN => n20899);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n5824, CK => CLK, Q => 
                           n18463, QN => n20900);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n5823, CK => CLK, Q => 
                           n18484, QN => n20901);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => n5950, CK => CLK, Q => 
                           n17156, QN => n21286);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => n5949, CK => CLK, Q => 
                           n17177, QN => n21287);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => n5948, CK => CLK, Q => 
                           n17198, QN => n21288);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => n5947, CK => CLK, Q => 
                           n17219, QN => n21289);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => n5946, CK => CLK, Q => 
                           n17240, QN => n21290);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => n5945, CK => CLK, Q => 
                           n17261, QN => n21291);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => n5944, CK => CLK, Q => 
                           n17282, QN => n21292);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => n5943, CK => CLK, Q => 
                           n17303, QN => n21293);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => n5942, CK => CLK, Q => 
                           n17324, QN => n21294);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => n5941, CK => CLK, Q => 
                           n17345, QN => n21295);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => n5940, CK => CLK, Q => 
                           n17366, QN => n21296);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => n5939, CK => CLK, Q => 
                           n17387, QN => n21297);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => n5938, CK => CLK, Q => 
                           n17408, QN => n21298);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => n5937, CK => CLK, Q => 
                           n17429, QN => n21299);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => n5936, CK => CLK, Q => 
                           n17450, QN => n21300);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => n5935, CK => CLK, Q => 
                           n17471, QN => n21301);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => n5934, CK => CLK, Q => 
                           n17492, QN => n21302);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => n5933, CK => CLK, Q => 
                           n17513, QN => n21303);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => n5932, CK => CLK, Q => 
                           n17534, QN => n21304);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => n5931, CK => CLK, Q => 
                           n17555, QN => n21305);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => n5930, CK => CLK, Q => 
                           n17576, QN => n21306);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => n5929, CK => CLK, Q => 
                           n17597, QN => n21307);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => n5928, CK => CLK, Q => 
                           n17618, QN => n21308);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => n5927, CK => CLK, Q => 
                           n17639, QN => n21309);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => n5926, CK => CLK, Q => 
                           n17660, QN => n21310);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => n5925, CK => CLK, Q => 
                           n17681, QN => n21311);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => n5924, CK => CLK, Q => 
                           n17702, QN => n21312);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => n5923, CK => CLK, Q => 
                           n17723, QN => n21313);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => n5922, CK => CLK, Q => 
                           n17744, QN => n21314);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => n5921, CK => CLK, Q => 
                           n17765, QN => n21315);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => n5920, CK => CLK, Q => 
                           n17786, QN => n21316);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => n5919, CK => CLK, Q => 
                           n17807, QN => n21317);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n5918, CK => CLK, Q => 
                           n17828, QN => n21318);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n5917, CK => CLK, Q => 
                           n17849, QN => n21319);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n5916, CK => CLK, Q => 
                           n17870, QN => n21320);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n5915, CK => CLK, Q => 
                           n17891, QN => n21321);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n5914, CK => CLK, Q => 
                           n17912, QN => n21322);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n5913, CK => CLK, Q => 
                           n17933, QN => n21323);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n5912, CK => CLK, Q => 
                           n17954, QN => n21324);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n5911, CK => CLK, Q => 
                           n17975, QN => n21325);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n5910, CK => CLK, Q => 
                           n17996, QN => n21326);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n5909, CK => CLK, Q => 
                           n18017, QN => n21327);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n5908, CK => CLK, Q => 
                           n18038, QN => n21328);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n5907, CK => CLK, Q => 
                           n18059, QN => n21329);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n5906, CK => CLK, Q => 
                           n18080, QN => n21330);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n5905, CK => CLK, Q => 
                           n18101, QN => n21331);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n5904, CK => CLK, Q => 
                           n18122, QN => n21332);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n5903, CK => CLK, Q => 
                           n18143, QN => n21333);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n5902, CK => CLK, Q => 
                           n18164, QN => n21334);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n5901, CK => CLK, Q => 
                           n18185, QN => n21335);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n5900, CK => CLK, Q => 
                           n18206, QN => n21336);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n5899, CK => CLK, Q => 
                           n18227, QN => n21337);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n5898, CK => CLK, Q => 
                           n18248, QN => n21338);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n5897, CK => CLK, Q => 
                           n18269, QN => n21339);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n5896, CK => CLK, Q => 
                           n18290, QN => n21340);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n5895, CK => CLK, Q => 
                           n18311, QN => n21341);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n5894, CK => CLK, Q => 
                           n18332, QN => n21342);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n5893, CK => CLK, Q => 
                           n18353, QN => n21343);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n5892, CK => CLK, Q => 
                           n18374, QN => n21344);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n5891, CK => CLK, Q => 
                           n18395, QN => n21345);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n5890, CK => CLK, Q => 
                           n18416, QN => n21346);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n5889, CK => CLK, Q => 
                           n18437, QN => n21347);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n5888, CK => CLK, Q => 
                           n18458, QN => n21348);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n5887, CK => CLK, Q => 
                           n18479, QN => n21349);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => n6974, CK => CLK, Q => 
                           n24477, QN => n19686);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => n6973, CK => CLK, Q => 
                           n24476, QN => n19687);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => n6972, CK => CLK, Q => 
                           n24475, QN => n19688);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => n6971, CK => CLK, Q => 
                           n24474, QN => n19689);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => n6970, CK => CLK, Q => 
                           n24853, QN => n19690);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => n6969, CK => CLK, Q => 
                           n24852, QN => n19691);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => n6968, CK => CLK, Q => 
                           n24851, QN => n19692);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => n6967, CK => CLK, Q => 
                           n24850, QN => n19693);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => n6966, CK => CLK, Q => 
                           n24849, QN => n19694);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => n6965, CK => CLK, Q => 
                           n24848, QN => n19695);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => n6964, CK => CLK, Q => 
                           n24847, QN => n19696);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => n6963, CK => CLK, Q => 
                           n24846, QN => n19697);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => n6962, CK => CLK, Q => 
                           n24845, QN => n19698);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => n6961, CK => CLK, Q => 
                           n24844, QN => n19699);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => n6960, CK => CLK, Q => 
                           n24843, QN => n19700);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => n6959, CK => CLK, Q => 
                           n24842, QN => n19701);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => n6958, CK => CLK, Q => 
                           n24841, QN => n19702);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => n6957, CK => CLK, Q => 
                           n24840, QN => n19703);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => n6956, CK => CLK, Q => 
                           n24839, QN => n19704);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => n6955, CK => CLK, Q => 
                           n24838, QN => n19705);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => n6954, CK => CLK, Q => 
                           n24837, QN => n19706);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => n6953, CK => CLK, Q => 
                           n24836, QN => n19707);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => n6952, CK => CLK, Q => 
                           n24835, QN => n19708);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => n6951, CK => CLK, Q => 
                           n24834, QN => n19709);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => n6950, CK => CLK, Q => 
                           n24833, QN => n19710);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => n6949, CK => CLK, Q => 
                           n24832, QN => n19711);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => n6948, CK => CLK, Q => 
                           n24831, QN => n19712);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => n6947, CK => CLK, Q => 
                           n24830, QN => n19713);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => n6946, CK => CLK, Q => 
                           n24829, QN => n19714);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => n6945, CK => CLK, Q => 
                           n24828, QN => n19715);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => n6944, CK => CLK, Q => 
                           n24827, QN => n19716);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => n6943, CK => CLK, Q => 
                           n24826, QN => n19717);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n6942, CK => CLK, Q => 
                           n24825, QN => n19718);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n6941, CK => CLK, Q => 
                           n24824, QN => n19719);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n6940, CK => CLK, Q => 
                           n24823, QN => n19720);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n6939, CK => CLK, Q => 
                           n24822, QN => n19721);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n6938, CK => CLK, Q => 
                           n24821, QN => n19722);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n6937, CK => CLK, Q => 
                           n24820, QN => n19723);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n6936, CK => CLK, Q => 
                           n24819, QN => n19724);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n6935, CK => CLK, Q => 
                           n24818, QN => n19725);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n6934, CK => CLK, Q => 
                           n24817, QN => n19726);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n6933, CK => CLK, Q => 
                           n24816, QN => n19727);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n6932, CK => CLK, Q => 
                           n24815, QN => n19728);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n6931, CK => CLK, Q => 
                           n24814, QN => n19729);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n6930, CK => CLK, Q => 
                           n24813, QN => n19730);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n6929, CK => CLK, Q => 
                           n24812, QN => n19731);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n6928, CK => CLK, Q => 
                           n24811, QN => n19732);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n6927, CK => CLK, Q => 
                           n24810, QN => n19733);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n6926, CK => CLK, Q => 
                           n24809, QN => n19734);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n6925, CK => CLK, Q => 
                           n24808, QN => n19735);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n6924, CK => CLK, Q => 
                           n24807, QN => n19736);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n6923, CK => CLK, Q => 
                           n24806, QN => n19737);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n6922, CK => CLK, Q => 
                           n24805, QN => n19738);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n6921, CK => CLK, Q => 
                           n24804, QN => n19739);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n6920, CK => CLK, Q => n24803
                           , QN => n19740);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n6919, CK => CLK, Q => n24802
                           , QN => n19741);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n6918, CK => CLK, Q => n24801
                           , QN => n19742);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n6917, CK => CLK, Q => n24800
                           , QN => n19743);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n6916, CK => CLK, Q => n24799
                           , QN => n19744);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n6915, CK => CLK, Q => n24798
                           , QN => n19745);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n6914, CK => CLK, Q => n24797
                           , QN => n19746);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n6913, CK => CLK, Q => n24796
                           , QN => n19747);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n6912, CK => CLK, Q => n24795
                           , QN => n19748);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n6911, CK => CLK, Q => n24794
                           , QN => n19749);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => n6014, CK => CLK, Q => 
                           n17157, QN => n21030);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => n6013, CK => CLK, Q => 
                           n17178, QN => n21031);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => n6012, CK => CLK, Q => 
                           n17199, QN => n21032);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => n6011, CK => CLK, Q => 
                           n17220, QN => n21033);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => n6010, CK => CLK, Q => 
                           n17241, QN => n21034);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => n6009, CK => CLK, Q => 
                           n17262, QN => n21035);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => n6008, CK => CLK, Q => 
                           n17283, QN => n21036);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => n6007, CK => CLK, Q => 
                           n17304, QN => n21037);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => n6006, CK => CLK, Q => 
                           n17325, QN => n21038);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => n6005, CK => CLK, Q => 
                           n17346, QN => n21039);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => n6004, CK => CLK, Q => 
                           n17367, QN => n21040);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => n6003, CK => CLK, Q => 
                           n17388, QN => n21041);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => n6002, CK => CLK, Q => 
                           n17409, QN => n21042);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => n6001, CK => CLK, Q => 
                           n17430, QN => n21043);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => n6000, CK => CLK, Q => 
                           n17451, QN => n21044);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => n5999, CK => CLK, Q => 
                           n17472, QN => n21045);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => n5998, CK => CLK, Q => 
                           n17493, QN => n21046);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => n5997, CK => CLK, Q => 
                           n17514, QN => n21047);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => n5996, CK => CLK, Q => 
                           n17535, QN => n21048);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => n5995, CK => CLK, Q => 
                           n17556, QN => n21049);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => n5994, CK => CLK, Q => 
                           n17577, QN => n21050);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => n5993, CK => CLK, Q => 
                           n17598, QN => n21051);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => n5992, CK => CLK, Q => 
                           n17619, QN => n21052);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => n5991, CK => CLK, Q => 
                           n17640, QN => n21053);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => n5990, CK => CLK, Q => 
                           n17661, QN => n21054);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => n5989, CK => CLK, Q => 
                           n17682, QN => n21055);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => n5988, CK => CLK, Q => 
                           n17703, QN => n21056);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => n5987, CK => CLK, Q => 
                           n17724, QN => n21057);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => n5986, CK => CLK, Q => 
                           n17745, QN => n21058);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => n5985, CK => CLK, Q => 
                           n17766, QN => n21059);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => n5984, CK => CLK, Q => 
                           n17787, QN => n21060);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => n5983, CK => CLK, Q => 
                           n17808, QN => n21061);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n5982, CK => CLK, Q => 
                           n17829, QN => n21062);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n5981, CK => CLK, Q => 
                           n17850, QN => n21063);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n5980, CK => CLK, Q => 
                           n17871, QN => n21064);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n5979, CK => CLK, Q => 
                           n17892, QN => n21065);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n5978, CK => CLK, Q => 
                           n17913, QN => n21066);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n5977, CK => CLK, Q => 
                           n17934, QN => n21067);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n5976, CK => CLK, Q => 
                           n17955, QN => n21068);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n5975, CK => CLK, Q => 
                           n17976, QN => n21069);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n5974, CK => CLK, Q => 
                           n17997, QN => n21070);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n5973, CK => CLK, Q => 
                           n18018, QN => n21071);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n5972, CK => CLK, Q => 
                           n18039, QN => n21072);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n5971, CK => CLK, Q => 
                           n18060, QN => n21073);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n5970, CK => CLK, Q => 
                           n18081, QN => n21074);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n5969, CK => CLK, Q => 
                           n18102, QN => n21075);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n5968, CK => CLK, Q => 
                           n18123, QN => n21076);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n5967, CK => CLK, Q => 
                           n18144, QN => n21077);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n5966, CK => CLK, Q => 
                           n18165, QN => n21078);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n5965, CK => CLK, Q => 
                           n18186, QN => n21079);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n5964, CK => CLK, Q => 
                           n18207, QN => n21080);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n5963, CK => CLK, Q => 
                           n18228, QN => n21081);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n5962, CK => CLK, Q => 
                           n18249, QN => n21082);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n5961, CK => CLK, Q => 
                           n18270, QN => n21083);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n5960, CK => CLK, Q => 
                           n18291, QN => n21084);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n5959, CK => CLK, Q => 
                           n18312, QN => n21085);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n5958, CK => CLK, Q => 
                           n18333, QN => n21086);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n5957, CK => CLK, Q => 
                           n18354, QN => n21087);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n5956, CK => CLK, Q => 
                           n18375, QN => n21088);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n5955, CK => CLK, Q => 
                           n18396, QN => n21089);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n5954, CK => CLK, Q => 
                           n18417, QN => n21090);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n5953, CK => CLK, Q => 
                           n18438, QN => n21091);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n5952, CK => CLK, Q => 
                           n18459, QN => n21092);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n5951, CK => CLK, Q => 
                           n18480, QN => n21093);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => n6462, CK => CLK, Q => 
                           n17148, QN => n20902);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => n6461, CK => CLK, Q => 
                           n17169, QN => n20903);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => n6460, CK => CLK, Q => 
                           n17190, QN => n20904);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => n6459, CK => CLK, Q => 
                           n17211, QN => n20905);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => n6458, CK => CLK, Q => 
                           n17232, QN => n20906);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => n6457, CK => CLK, Q => 
                           n17253, QN => n20907);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => n6456, CK => CLK, Q => 
                           n17274, QN => n20908);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => n6455, CK => CLK, Q => 
                           n17295, QN => n20909);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => n6454, CK => CLK, Q => 
                           n17316, QN => n20910);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => n6453, CK => CLK, Q => 
                           n17337, QN => n20911);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => n6452, CK => CLK, Q => 
                           n17358, QN => n20912);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => n6451, CK => CLK, Q => 
                           n17379, QN => n20913);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => n6450, CK => CLK, Q => 
                           n17400, QN => n20914);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => n6449, CK => CLK, Q => 
                           n17421, QN => n20915);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => n6448, CK => CLK, Q => 
                           n17442, QN => n20916);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => n6447, CK => CLK, Q => 
                           n17463, QN => n20917);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => n6446, CK => CLK, Q => 
                           n17484, QN => n20918);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => n6445, CK => CLK, Q => 
                           n17505, QN => n20919);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => n6444, CK => CLK, Q => 
                           n17526, QN => n20920);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => n6443, CK => CLK, Q => 
                           n17547, QN => n20921);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => n6442, CK => CLK, Q => 
                           n17568, QN => n20922);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => n6441, CK => CLK, Q => 
                           n17589, QN => n20923);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => n6440, CK => CLK, Q => 
                           n17610, QN => n20924);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => n6439, CK => CLK, Q => 
                           n17631, QN => n20925);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => n6438, CK => CLK, Q => 
                           n17652, QN => n20926);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => n6437, CK => CLK, Q => 
                           n17673, QN => n20927);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => n6436, CK => CLK, Q => 
                           n17694, QN => n20928);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => n6435, CK => CLK, Q => 
                           n17715, QN => n20929);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => n6434, CK => CLK, Q => 
                           n17736, QN => n20930);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => n6433, CK => CLK, Q => 
                           n17757, QN => n20931);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => n6432, CK => CLK, Q => 
                           n17778, QN => n20932);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => n6431, CK => CLK, Q => 
                           n17799, QN => n20933);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n6430, CK => CLK, Q => 
                           n17820, QN => n20934);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n6429, CK => CLK, Q => 
                           n17841, QN => n20935);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n6428, CK => CLK, Q => 
                           n17862, QN => n20936);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n6427, CK => CLK, Q => 
                           n17883, QN => n20937);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n6426, CK => CLK, Q => 
                           n17904, QN => n20938);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n6425, CK => CLK, Q => 
                           n17925, QN => n20939);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n6424, CK => CLK, Q => 
                           n17946, QN => n20940);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n6423, CK => CLK, Q => 
                           n17967, QN => n20941);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n6422, CK => CLK, Q => 
                           n17988, QN => n20942);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n6421, CK => CLK, Q => 
                           n18009, QN => n20943);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n6420, CK => CLK, Q => 
                           n18030, QN => n20944);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n6419, CK => CLK, Q => 
                           n18051, QN => n20945);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n6418, CK => CLK, Q => 
                           n18072, QN => n20946);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n6417, CK => CLK, Q => 
                           n18093, QN => n20947);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n6416, CK => CLK, Q => 
                           n18114, QN => n20948);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n6415, CK => CLK, Q => 
                           n18135, QN => n20949);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n6414, CK => CLK, Q => 
                           n18156, QN => n20950);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n6413, CK => CLK, Q => 
                           n18177, QN => n20951);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n6412, CK => CLK, Q => 
                           n18198, QN => n20952);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n6411, CK => CLK, Q => 
                           n18219, QN => n20953);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n6410, CK => CLK, Q => 
                           n18240, QN => n20954);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n6409, CK => CLK, Q => 
                           n18261, QN => n20955);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n6408, CK => CLK, Q => 
                           n18282, QN => n20956);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n6407, CK => CLK, Q => 
                           n18303, QN => n20957);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n6406, CK => CLK, Q => 
                           n18324, QN => n20958);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n6405, CK => CLK, Q => 
                           n18345, QN => n20959);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n6404, CK => CLK, Q => 
                           n18366, QN => n20960);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n6403, CK => CLK, Q => 
                           n18387, QN => n20961);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n6402, CK => CLK, Q => 
                           n18408, QN => n20962);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n6401, CK => CLK, Q => 
                           n18429, QN => n20963);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n6400, CK => CLK, Q => 
                           n18450, QN => n20964);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n6399, CK => CLK, Q => 
                           n18471, QN => n20965);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => n6590, CK => CLK, Q => 
                           n17149, QN => n21414);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => n6589, CK => CLK, Q => 
                           n17170, QN => n21415);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => n6588, CK => CLK, Q => 
                           n17191, QN => n21416);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => n6587, CK => CLK, Q => 
                           n17212, QN => n21417);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => n6586, CK => CLK, Q => 
                           n17233, QN => n21418);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => n6585, CK => CLK, Q => 
                           n17254, QN => n21419);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => n6584, CK => CLK, Q => 
                           n17275, QN => n21420);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => n6583, CK => CLK, Q => 
                           n17296, QN => n21421);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => n6582, CK => CLK, Q => 
                           n17317, QN => n21422);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => n6581, CK => CLK, Q => 
                           n17338, QN => n21423);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => n6580, CK => CLK, Q => 
                           n17359, QN => n21424);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => n6579, CK => CLK, Q => 
                           n17380, QN => n21425);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => n6578, CK => CLK, Q => 
                           n17401, QN => n21426);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => n6577, CK => CLK, Q => 
                           n17422, QN => n21427);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => n6576, CK => CLK, Q => 
                           n17443, QN => n21428);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => n6575, CK => CLK, Q => 
                           n17464, QN => n21429);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => n6574, CK => CLK, Q => 
                           n17485, QN => n21430);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => n6573, CK => CLK, Q => 
                           n17506, QN => n21431);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => n6572, CK => CLK, Q => 
                           n17527, QN => n21432);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => n6571, CK => CLK, Q => 
                           n17548, QN => n21433);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => n6570, CK => CLK, Q => 
                           n17569, QN => n21434);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => n6569, CK => CLK, Q => 
                           n17590, QN => n21435);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => n6568, CK => CLK, Q => 
                           n17611, QN => n21436);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => n6567, CK => CLK, Q => 
                           n17632, QN => n21437);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => n6566, CK => CLK, Q => 
                           n17653, QN => n21438);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => n6565, CK => CLK, Q => 
                           n17674, QN => n21439);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => n6564, CK => CLK, Q => 
                           n17695, QN => n21440);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => n6563, CK => CLK, Q => 
                           n17716, QN => n21441);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => n6562, CK => CLK, Q => 
                           n17737, QN => n21442);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => n6561, CK => CLK, Q => 
                           n17758, QN => n21443);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => n6560, CK => CLK, Q => 
                           n17779, QN => n21444);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => n6559, CK => CLK, Q => 
                           n17800, QN => n21445);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n6558, CK => CLK, Q => 
                           n17821, QN => n21446);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n6557, CK => CLK, Q => 
                           n17842, QN => n21447);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n6556, CK => CLK, Q => 
                           n17863, QN => n21448);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n6555, CK => CLK, Q => 
                           n17884, QN => n21449);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n6554, CK => CLK, Q => 
                           n17905, QN => n21450);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n6553, CK => CLK, Q => 
                           n17926, QN => n21451);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n6552, CK => CLK, Q => 
                           n17947, QN => n21452);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n6551, CK => CLK, Q => 
                           n17968, QN => n21453);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n6550, CK => CLK, Q => 
                           n17989, QN => n21454);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n6549, CK => CLK, Q => 
                           n18010, QN => n21455);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n6548, CK => CLK, Q => 
                           n18031, QN => n21456);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n6547, CK => CLK, Q => 
                           n18052, QN => n21457);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n6546, CK => CLK, Q => 
                           n18073, QN => n21458);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n6545, CK => CLK, Q => 
                           n18094, QN => n21459);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n6544, CK => CLK, Q => 
                           n18115, QN => n21460);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n6543, CK => CLK, Q => 
                           n18136, QN => n21461);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n6542, CK => CLK, Q => 
                           n18157, QN => n21462);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n6541, CK => CLK, Q => 
                           n18178, QN => n21463);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n6540, CK => CLK, Q => 
                           n18199, QN => n21464);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n6539, CK => CLK, Q => 
                           n18220, QN => n21465);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n6538, CK => CLK, Q => 
                           n18241, QN => n21466);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n6537, CK => CLK, Q => 
                           n18262, QN => n21467);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n6536, CK => CLK, Q => 
                           n18283, QN => n21468);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n6535, CK => CLK, Q => 
                           n18304, QN => n21469);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n6534, CK => CLK, Q => 
                           n18325, QN => n21470);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n6533, CK => CLK, Q => 
                           n18346, QN => n21471);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n6532, CK => CLK, Q => 
                           n18367, QN => n21472);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n6531, CK => CLK, Q => 
                           n18388, QN => n21473);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n6530, CK => CLK, Q => 
                           n18409, QN => n21474);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n6529, CK => CLK, Q => 
                           n18430, QN => n21475);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n6528, CK => CLK, Q => 
                           n18451, QN => n21476);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n6527, CK => CLK, Q => 
                           n18472, QN => n21477);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => n5566, CK => CLK, Q => 
                           n24441, QN => n20262);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => n5565, CK => CLK, Q => 
                           n24439, QN => n20263);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => n5564, CK => CLK, Q => 
                           n24437, QN => n20264);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => n5563, CK => CLK, Q => 
                           n24435, QN => n20265);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => n5694, CK => CLK, Q => 
                           n24085, QN => n20266);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => n5693, CK => CLK, Q => 
                           n24083, QN => n20267);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => n5692, CK => CLK, Q => 
                           n24081, QN => n20268);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => n5691, CK => CLK, Q => 
                           n24079, QN => n20269);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => n5562, CK => CLK, Q => 
                           n24433, QN => n20462);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => n5561, CK => CLK, Q => 
                           n24431, QN => n20463);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => n5560, CK => CLK, Q => 
                           n24429, QN => n20464);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => n5559, CK => CLK, Q => 
                           n24427, QN => n20465);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => n5558, CK => CLK, Q => 
                           n24425, QN => n20466);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => n5557, CK => CLK, Q => 
                           n24423, QN => n20467);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => n5556, CK => CLK, Q => 
                           n24421, QN => n20468);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => n5555, CK => CLK, Q => 
                           n24419, QN => n20469);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => n5554, CK => CLK, Q => 
                           n24417, QN => n20470);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => n5553, CK => CLK, Q => 
                           n24415, QN => n20471);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => n5552, CK => CLK, Q => 
                           n24413, QN => n20472);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => n5551, CK => CLK, Q => 
                           n24411, QN => n20473);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => n5550, CK => CLK, Q => 
                           n24409, QN => n20474);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => n5549, CK => CLK, Q => 
                           n24407, QN => n20475);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => n5548, CK => CLK, Q => 
                           n24405, QN => n20476);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => n5547, CK => CLK, Q => 
                           n24403, QN => n20477);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => n5546, CK => CLK, Q => 
                           n24401, QN => n20478);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => n5545, CK => CLK, Q => 
                           n24399, QN => n20479);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => n5544, CK => CLK, Q => 
                           n24397, QN => n20480);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => n5543, CK => CLK, Q => 
                           n24395, QN => n20481);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => n5542, CK => CLK, Q => 
                           n24393, QN => n20482);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => n5541, CK => CLK, Q => 
                           n24391, QN => n20483);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => n5540, CK => CLK, Q => 
                           n24389, QN => n20484);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => n5539, CK => CLK, Q => 
                           n24387, QN => n20485);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => n5538, CK => CLK, Q => 
                           n24385, QN => n20486);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => n5537, CK => CLK, Q => 
                           n24383, QN => n20487);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => n5536, CK => CLK, Q => 
                           n24381, QN => n20488);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => n5535, CK => CLK, Q => 
                           n24379, QN => n20489);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n5534, CK => CLK, Q => 
                           n24377, QN => n20490);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n5533, CK => CLK, Q => 
                           n24375, QN => n20491);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n5532, CK => CLK, Q => 
                           n24373, QN => n20492);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n5531, CK => CLK, Q => 
                           n24371, QN => n20493);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n5530, CK => CLK, Q => 
                           n24369, QN => n20494);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n5529, CK => CLK, Q => 
                           n24367, QN => n20495);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n5528, CK => CLK, Q => 
                           n24365, QN => n20496);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n5527, CK => CLK, Q => 
                           n24363, QN => n20497);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n5526, CK => CLK, Q => 
                           n24361, QN => n20498);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n5525, CK => CLK, Q => 
                           n24359, QN => n20499);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n5524, CK => CLK, Q => 
                           n24357, QN => n20500);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n5523, CK => CLK, Q => 
                           n24355, QN => n20501);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n5522, CK => CLK, Q => 
                           n24353, QN => n20502);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n5521, CK => CLK, Q => 
                           n24351, QN => n20503);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n5520, CK => CLK, Q => 
                           n24349, QN => n20504);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n5519, CK => CLK, Q => 
                           n24347, QN => n20505);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n5518, CK => CLK, Q => 
                           n24345, QN => n20506);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n5517, CK => CLK, Q => 
                           n24343, QN => n20507);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n5516, CK => CLK, Q => 
                           n24341, QN => n20508);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n5515, CK => CLK, Q => 
                           n24339, QN => n20509);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n5514, CK => CLK, Q => 
                           n24465, QN => n20510);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n5513, CK => CLK, Q => 
                           n24463, QN => n20511);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n5512, CK => CLK, Q => 
                           n24461, QN => n20512);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n5511, CK => CLK, Q => 
                           n24459, QN => n20513);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n5510, CK => CLK, Q => 
                           n24457, QN => n20514);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n5509, CK => CLK, Q => 
                           n24455, QN => n20515);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n5508, CK => CLK, Q => 
                           n24453, QN => n20516);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n5507, CK => CLK, Q => 
                           n24451, QN => n20517);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n5506, CK => CLK, Q => 
                           n24449, QN => n20518);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n5505, CK => CLK, Q => 
                           n24447, QN => n20519);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n5504, CK => CLK, Q => 
                           n24445, QN => n20520);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n5503, CK => CLK, Q => 
                           n24443, QN => n20521);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => n5690, CK => CLK, Q => 
                           n24205, QN => n20522);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => n5689, CK => CLK, Q => 
                           n24203, QN => n20523);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => n5688, CK => CLK, Q => 
                           n24201, QN => n20524);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => n5687, CK => CLK, Q => 
                           n24199, QN => n20525);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => n5686, CK => CLK, Q => 
                           n24197, QN => n20526);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => n5685, CK => CLK, Q => 
                           n24195, QN => n20527);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => n5684, CK => CLK, Q => 
                           n24193, QN => n20528);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => n5683, CK => CLK, Q => 
                           n24191, QN => n20529);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => n5682, CK => CLK, Q => 
                           n24189, QN => n20530);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => n5681, CK => CLK, Q => 
                           n24187, QN => n20531);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => n5680, CK => CLK, Q => 
                           n24185, QN => n20532);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => n5679, CK => CLK, Q => 
                           n24183, QN => n20533);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => n5678, CK => CLK, Q => 
                           n24181, QN => n20534);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => n5677, CK => CLK, Q => 
                           n24179, QN => n20535);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => n5676, CK => CLK, Q => 
                           n24177, QN => n20536);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => n5675, CK => CLK, Q => 
                           n24175, QN => n20537);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => n5674, CK => CLK, Q => 
                           n24173, QN => n20538);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => n5673, CK => CLK, Q => 
                           n24171, QN => n20539);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => n5672, CK => CLK, Q => 
                           n24169, QN => n20540);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => n5671, CK => CLK, Q => 
                           n24167, QN => n20541);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => n5670, CK => CLK, Q => 
                           n24165, QN => n20542);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => n5669, CK => CLK, Q => 
                           n24163, QN => n20543);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => n5668, CK => CLK, Q => 
                           n24161, QN => n20544);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => n5667, CK => CLK, Q => 
                           n24159, QN => n20545);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => n5666, CK => CLK, Q => 
                           n24157, QN => n20546);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => n5665, CK => CLK, Q => 
                           n24155, QN => n20547);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => n5664, CK => CLK, Q => 
                           n24153, QN => n20548);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => n5663, CK => CLK, Q => 
                           n24151, QN => n20549);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n5662, CK => CLK, Q => 
                           n24149, QN => n20550);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n5661, CK => CLK, Q => 
                           n24147, QN => n20551);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n5660, CK => CLK, Q => 
                           n24145, QN => n20552);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n5659, CK => CLK, Q => 
                           n24143, QN => n20553);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n5658, CK => CLK, Q => 
                           n24141, QN => n20554);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n5657, CK => CLK, Q => 
                           n24139, QN => n20555);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n5656, CK => CLK, Q => 
                           n24137, QN => n20556);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n5655, CK => CLK, Q => 
                           n24135, QN => n20557);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n5654, CK => CLK, Q => 
                           n24133, QN => n20558);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n5653, CK => CLK, Q => 
                           n24131, QN => n20559);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n5652, CK => CLK, Q => 
                           n24129, QN => n20560);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n5651, CK => CLK, Q => 
                           n24127, QN => n20561);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n5650, CK => CLK, Q => 
                           n24125, QN => n20562);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n5649, CK => CLK, Q => 
                           n24123, QN => n20563);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n5648, CK => CLK, Q => 
                           n24121, QN => n20564);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n5647, CK => CLK, Q => 
                           n24119, QN => n20565);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n5646, CK => CLK, Q => 
                           n24117, QN => n20566);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n5645, CK => CLK, Q => 
                           n24115, QN => n20567);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n5644, CK => CLK, Q => 
                           n24113, QN => n20568);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n5643, CK => CLK, Q => 
                           n24111, QN => n20569);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n5642, CK => CLK, Q => 
                           n24109, QN => n20570);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n5641, CK => CLK, Q => 
                           n24107, QN => n20571);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n5640, CK => CLK, Q => 
                           n24105, QN => n20572);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n5639, CK => CLK, Q => 
                           n24103, QN => n20573);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n5638, CK => CLK, Q => 
                           n24101, QN => n20574);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n5637, CK => CLK, Q => 
                           n24099, QN => n20575);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n5636, CK => CLK, Q => 
                           n24097, QN => n20576);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n5635, CK => CLK, Q => 
                           n24095, QN => n20577);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n5634, CK => CLK, Q => 
                           n24093, QN => n20578);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n5633, CK => CLK, Q => 
                           n24091, QN => n20579);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n5632, CK => CLK, Q => 
                           n24089, QN => n20580);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n5631, CK => CLK, Q => 
                           n24087, QN => n20581);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => n6846, CK => CLK, Q => 
                           n23957, QN => n20582);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => n6845, CK => CLK, Q => 
                           n23956, QN => n20583);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => n6844, CK => CLK, Q => 
                           n23955, QN => n20584);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => n6843, CK => CLK, Q => 
                           n23954, QN => n20585);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => n6842, CK => CLK, Q => 
                           n24077, QN => n20586);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => n6841, CK => CLK, Q => 
                           n24076, QN => n20587);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => n6840, CK => CLK, Q => 
                           n24075, QN => n20588);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => n6839, CK => CLK, Q => 
                           n24074, QN => n20589);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => n6838, CK => CLK, Q => 
                           n24073, QN => n20590);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => n6837, CK => CLK, Q => 
                           n24072, QN => n20591);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => n6836, CK => CLK, Q => 
                           n24071, QN => n20592);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => n6835, CK => CLK, Q => 
                           n24070, QN => n20593);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => n6834, CK => CLK, Q => 
                           n24069, QN => n20594);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => n6833, CK => CLK, Q => 
                           n24068, QN => n20595);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => n6832, CK => CLK, Q => 
                           n24067, QN => n20596);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => n6831, CK => CLK, Q => 
                           n24066, QN => n20597);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => n6830, CK => CLK, Q => 
                           n24065, QN => n20598);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => n6829, CK => CLK, Q => 
                           n24064, QN => n20599);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => n6828, CK => CLK, Q => 
                           n24063, QN => n20600);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => n6827, CK => CLK, Q => 
                           n24062, QN => n20601);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => n6826, CK => CLK, Q => 
                           n24061, QN => n20602);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => n6825, CK => CLK, Q => 
                           n24060, QN => n20603);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => n6824, CK => CLK, Q => 
                           n24059, QN => n20604);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => n6823, CK => CLK, Q => 
                           n24058, QN => n20605);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => n6822, CK => CLK, Q => 
                           n24057, QN => n20606);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => n6821, CK => CLK, Q => 
                           n24056, QN => n20607);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => n6820, CK => CLK, Q => 
                           n24055, QN => n20608);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => n6819, CK => CLK, Q => 
                           n24054, QN => n20609);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => n6818, CK => CLK, Q => 
                           n24053, QN => n20610);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => n6817, CK => CLK, Q => 
                           n24052, QN => n20611);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => n6816, CK => CLK, Q => 
                           n24051, QN => n20612);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => n6815, CK => CLK, Q => 
                           n24050, QN => n20613);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n6814, CK => CLK, Q => 
                           n24049, QN => n20614);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n6813, CK => CLK, Q => 
                           n24048, QN => n20615);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n6812, CK => CLK, Q => 
                           n24047, QN => n20616);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n6811, CK => CLK, Q => 
                           n24046, QN => n20617);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n6810, CK => CLK, Q => 
                           n24045, QN => n20618);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n6809, CK => CLK, Q => 
                           n24044, QN => n20619);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n6808, CK => CLK, Q => 
                           n24043, QN => n20620);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n6807, CK => CLK, Q => 
                           n24042, QN => n20621);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n6806, CK => CLK, Q => 
                           n24041, QN => n20622);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n6805, CK => CLK, Q => 
                           n24040, QN => n20623);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n6804, CK => CLK, Q => 
                           n24039, QN => n20624);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n6803, CK => CLK, Q => 
                           n24038, QN => n20625);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n6802, CK => CLK, Q => 
                           n24037, QN => n20626);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n6801, CK => CLK, Q => 
                           n24036, QN => n20627);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n6800, CK => CLK, Q => 
                           n24035, QN => n20628);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n6799, CK => CLK, Q => 
                           n24034, QN => n20629);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n6798, CK => CLK, Q => 
                           n24033, QN => n20630);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n6797, CK => CLK, Q => 
                           n24032, QN => n20631);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n6796, CK => CLK, Q => 
                           n24031, QN => n20632);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n6795, CK => CLK, Q => 
                           n24030, QN => n20633);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n6794, CK => CLK, Q => 
                           n24029, QN => n20634);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n6793, CK => CLK, Q => 
                           n24028, QN => n20635);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n6792, CK => CLK, Q => 
                           n24027, QN => n20636);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n6791, CK => CLK, Q => 
                           n24026, QN => n20637);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n6790, CK => CLK, Q => 
                           n24025, QN => n20638);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n6789, CK => CLK, Q => 
                           n24024, QN => n20639);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n6788, CK => CLK, Q => 
                           n24023, QN => n20640);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n6787, CK => CLK, Q => 
                           n24022, QN => n20641);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n6786, CK => CLK, Q => 
                           n24021, QN => n20642);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n6785, CK => CLK, Q => 
                           n24020, QN => n20643);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n6784, CK => CLK, Q => 
                           n24019, QN => n20644);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n6783, CK => CLK, Q => 
                           n24018, QN => n20645);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => n7102, CK => CLK, Q => 
                           n24481, QN => n19622);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => n7101, CK => CLK, Q => 
                           n24480, QN => n19623);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => n7100, CK => CLK, Q => 
                           n24479, QN => n19624);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => n7099, CK => CLK, Q => 
                           n24478, QN => n19625);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => n7098, CK => CLK, Q => 
                           n24913, QN => n19626);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => n7097, CK => CLK, Q => 
                           n24912, QN => n19627);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => n7096, CK => CLK, Q => 
                           n24911, QN => n19628);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => n7095, CK => CLK, Q => 
                           n24910, QN => n19629);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => n7094, CK => CLK, Q => 
                           n24909, QN => n19630);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => n7093, CK => CLK, Q => 
                           n24908, QN => n19631);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => n7092, CK => CLK, Q => 
                           n24907, QN => n19632);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => n7091, CK => CLK, Q => 
                           n24906, QN => n19633);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => n7090, CK => CLK, Q => 
                           n24905, QN => n19634);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => n7089, CK => CLK, Q => 
                           n24904, QN => n19635);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => n7088, CK => CLK, Q => 
                           n24903, QN => n19636);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => n7087, CK => CLK, Q => 
                           n24902, QN => n19637);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => n7086, CK => CLK, Q => 
                           n24901, QN => n19638);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => n7085, CK => CLK, Q => 
                           n24900, QN => n19639);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => n7084, CK => CLK, Q => 
                           n24899, QN => n19640);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => n7083, CK => CLK, Q => 
                           n24898, QN => n19641);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => n7082, CK => CLK, Q => 
                           n24897, QN => n19642);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => n7081, CK => CLK, Q => 
                           n24896, QN => n19643);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => n7080, CK => CLK, Q => 
                           n24895, QN => n19644);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => n7079, CK => CLK, Q => 
                           n24894, QN => n19645);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => n7078, CK => CLK, Q => 
                           n24893, QN => n19646);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => n7077, CK => CLK, Q => 
                           n24892, QN => n19647);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => n7076, CK => CLK, Q => 
                           n24891, QN => n19648);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => n7075, CK => CLK, Q => 
                           n24890, QN => n19649);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => n7074, CK => CLK, Q => 
                           n24889, QN => n19650);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => n7073, CK => CLK, Q => 
                           n24888, QN => n19651);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => n7072, CK => CLK, Q => 
                           n24887, QN => n19652);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => n7071, CK => CLK, Q => 
                           n24886, QN => n19653);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n7070, CK => CLK, Q => 
                           n24885, QN => n19654);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n7069, CK => CLK, Q => 
                           n24884, QN => n19655);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n7068, CK => CLK, Q => 
                           n24883, QN => n19656);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n7067, CK => CLK, Q => 
                           n24882, QN => n19657);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n7066, CK => CLK, Q => 
                           n24881, QN => n19658);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n7065, CK => CLK, Q => 
                           n24880, QN => n19659);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n7064, CK => CLK, Q => 
                           n24879, QN => n19660);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n7063, CK => CLK, Q => 
                           n24878, QN => n19661);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n7062, CK => CLK, Q => 
                           n24877, QN => n19662);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n7061, CK => CLK, Q => 
                           n24876, QN => n19663);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n7060, CK => CLK, Q => 
                           n24875, QN => n19664);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n7059, CK => CLK, Q => 
                           n24874, QN => n19665);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n7058, CK => CLK, Q => 
                           n24873, QN => n19666);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n7057, CK => CLK, Q => 
                           n24872, QN => n19667);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n7056, CK => CLK, Q => 
                           n24871, QN => n19668);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n7055, CK => CLK, Q => 
                           n24870, QN => n19669);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n7054, CK => CLK, Q => 
                           n24869, QN => n19670);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n7053, CK => CLK, Q => 
                           n24868, QN => n19671);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n7052, CK => CLK, Q => 
                           n24867, QN => n19672);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n7051, CK => CLK, Q => 
                           n24866, QN => n19673);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n7050, CK => CLK, Q => 
                           n24865, QN => n19674);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n7049, CK => CLK, Q => 
                           n24864, QN => n19675);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n7048, CK => CLK, Q => n24863
                           , QN => n19676);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n7047, CK => CLK, Q => n24862
                           , QN => n19677);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n7046, CK => CLK, Q => n24861
                           , QN => n19678);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n7045, CK => CLK, Q => n24860
                           , QN => n19679);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n7044, CK => CLK, Q => n24859
                           , QN => n19680);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n7043, CK => CLK, Q => n24858
                           , QN => n19681);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n7042, CK => CLK, Q => n24857
                           , QN => n19682);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n7041, CK => CLK, Q => n24856
                           , QN => n19683);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n7040, CK => CLK, Q => n24855
                           , QN => n19684);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n7039, CK => CLK, Q => n24854
                           , QN => n19685);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n7294, CK => CLK, Q => 
                           n24311, QN => n20198);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n7293, CK => CLK, Q => 
                           n24308, QN => n20199);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n7292, CK => CLK, Q => 
                           n24305, QN => n20200);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n7291, CK => CLK, Q => 
                           n24302, QN => n20201);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n7290, CK => CLK, Q => 
                           n24300, QN => n20202);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n7289, CK => CLK, Q => 
                           n24298, QN => n20203);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n7288, CK => CLK, Q => 
                           n24296, QN => n20204);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n7287, CK => CLK, Q => 
                           n24294, QN => n20205);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n7286, CK => CLK, Q => 
                           n24292, QN => n20206);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n7285, CK => CLK, Q => 
                           n24290, QN => n20207);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n7284, CK => CLK, Q => 
                           n24288, QN => n20208);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n7283, CK => CLK, Q => 
                           n24286, QN => n20209);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n7282, CK => CLK, Q => 
                           n24284, QN => n20210);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n7281, CK => CLK, Q => 
                           n24282, QN => n20211);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n7280, CK => CLK, Q => 
                           n24280, QN => n20212);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n7279, CK => CLK, Q => 
                           n24278, QN => n20213);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n7278, CK => CLK, Q => 
                           n24276, QN => n20214);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n7277, CK => CLK, Q => 
                           n24274, QN => n20215);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n7276, CK => CLK, Q => 
                           n24272, QN => n20216);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n7275, CK => CLK, Q => 
                           n24270, QN => n20217);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n7274, CK => CLK, Q => 
                           n24268, QN => n20218);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n7273, CK => CLK, Q => 
                           n24266, QN => n20219);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n7272, CK => CLK, Q => 
                           n24264, QN => n20220);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n7271, CK => CLK, Q => 
                           n24262, QN => n20221);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n7270, CK => CLK, Q => 
                           n24260, QN => n20222);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n7269, CK => CLK, Q => 
                           n24258, QN => n20223);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n7268, CK => CLK, Q => 
                           n24256, QN => n20224);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n7267, CK => CLK, Q => 
                           n24254, QN => n20225);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n7266, CK => CLK, Q => 
                           n24252, QN => n20226);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n7265, CK => CLK, Q => 
                           n24250, QN => n20227);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n7264, CK => CLK, Q => 
                           n24248, QN => n20228);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n7263, CK => CLK, Q => 
                           n24246, QN => n20229);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n7262, CK => CLK, Q => 
                           n24244, QN => n20230);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n7261, CK => CLK, Q => 
                           n24242, QN => n20231);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n7260, CK => CLK, Q => 
                           n24240, QN => n20232);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n7259, CK => CLK, Q => 
                           n24238, QN => n20233);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n7258, CK => CLK, Q => 
                           n24236, QN => n20234);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n7257, CK => CLK, Q => 
                           n24234, QN => n20235);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n7256, CK => CLK, Q => 
                           n24232, QN => n20236);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n7255, CK => CLK, Q => 
                           n24230, QN => n20237);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n7254, CK => CLK, Q => 
                           n24228, QN => n20238);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n7253, CK => CLK, Q => 
                           n24226, QN => n20239);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n7252, CK => CLK, Q => 
                           n24224, QN => n20240);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n7251, CK => CLK, Q => 
                           n24222, QN => n20241);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n7250, CK => CLK, Q => 
                           n24220, QN => n20242);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n7249, CK => CLK, Q => 
                           n24218, QN => n20243);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n7248, CK => CLK, Q => 
                           n24216, QN => n20244);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n7247, CK => CLK, Q => 
                           n24214, QN => n20245);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n7246, CK => CLK, Q => 
                           n24212, QN => n20246);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n7245, CK => CLK, Q => 
                           n24210, QN => n20247);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n7244, CK => CLK, Q => 
                           n24208, QN => n20248);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n7243, CK => CLK, Q => 
                           n24206, QN => n20249);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n7242, CK => CLK, Q => 
                           n24336, QN => n20250);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n7241, CK => CLK, Q => 
                           n24334, QN => n20251);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n7240, CK => CLK, Q => n24332
                           , QN => n20252);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n7239, CK => CLK, Q => n24330
                           , QN => n20253);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n7238, CK => CLK, Q => n24328
                           , QN => n20254);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n7237, CK => CLK, Q => n24326
                           , QN => n20255);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n7236, CK => CLK, Q => n24324
                           , QN => n20256);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n7235, CK => CLK, Q => n24322
                           , QN => n20257);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n7234, CK => CLK, Q => n24320
                           , QN => n20258);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n7233, CK => CLK, Q => n24318
                           , QN => n20259);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n7232, CK => CLK, Q => n24316
                           , QN => n20260);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n7231, CK => CLK, Q => n24314
                           , QN => n20261);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => n6078, CK => CLK, Q => 
                           n24613, QN => n19877);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => n6077, CK => CLK, Q => 
                           n24611, QN => n19878);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => n6076, CK => CLK, Q => 
                           n24609, QN => n19879);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => n6075, CK => CLK, Q => 
                           n24607, QN => n19880);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => n6074, CK => CLK, Q => 
                           n24673, QN => n19881);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => n6073, CK => CLK, Q => 
                           n24672, QN => n19882);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => n6072, CK => CLK, Q => 
                           n24671, QN => n19883);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => n6071, CK => CLK, Q => 
                           n24670, QN => n19884);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => n6070, CK => CLK, Q => 
                           n24669, QN => n19885);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => n6069, CK => CLK, Q => 
                           n24668, QN => n19886);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => n6068, CK => CLK, Q => 
                           n24667, QN => n19887);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => n6067, CK => CLK, Q => 
                           n24666, QN => n19888);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => n6066, CK => CLK, Q => 
                           n24665, QN => n19889);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => n6065, CK => CLK, Q => 
                           n24664, QN => n19890);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => n6064, CK => CLK, Q => 
                           n24663, QN => n19891);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => n6063, CK => CLK, Q => 
                           n24662, QN => n19892);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => n6062, CK => CLK, Q => 
                           n24661, QN => n19893);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => n6061, CK => CLK, Q => 
                           n24660, QN => n19894);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => n6060, CK => CLK, Q => 
                           n24659, QN => n19895);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => n6059, CK => CLK, Q => 
                           n24658, QN => n19896);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => n6058, CK => CLK, Q => 
                           n24657, QN => n19897);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => n6057, CK => CLK, Q => 
                           n24656, QN => n19898);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => n6056, CK => CLK, Q => 
                           n24655, QN => n19899);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => n6055, CK => CLK, Q => 
                           n24654, QN => n19900);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => n6054, CK => CLK, Q => 
                           n24653, QN => n19901);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => n6053, CK => CLK, Q => 
                           n24652, QN => n19902);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => n6052, CK => CLK, Q => 
                           n24651, QN => n19903);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => n6051, CK => CLK, Q => 
                           n24650, QN => n19904);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => n6050, CK => CLK, Q => 
                           n24649, QN => n19905);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => n6049, CK => CLK, Q => 
                           n24648, QN => n19906);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => n6048, CK => CLK, Q => 
                           n24647, QN => n19907);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => n6047, CK => CLK, Q => 
                           n24646, QN => n19908);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n6046, CK => CLK, Q => 
                           n24645, QN => n19909);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n6045, CK => CLK, Q => 
                           n24644, QN => n19910);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n6044, CK => CLK, Q => 
                           n24643, QN => n19911);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n6043, CK => CLK, Q => 
                           n24642, QN => n19912);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n6042, CK => CLK, Q => 
                           n24641, QN => n19913);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n6041, CK => CLK, Q => 
                           n24640, QN => n19914);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n6040, CK => CLK, Q => 
                           n24639, QN => n19915);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n6039, CK => CLK, Q => 
                           n24638, QN => n19916);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n6038, CK => CLK, Q => 
                           n24637, QN => n19917);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n6037, CK => CLK, Q => 
                           n24636, QN => n19918);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n6036, CK => CLK, Q => 
                           n24635, QN => n19919);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n6035, CK => CLK, Q => 
                           n24634, QN => n19920);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n6034, CK => CLK, Q => 
                           n24633, QN => n19921);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n6033, CK => CLK, Q => 
                           n24632, QN => n19922);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n6032, CK => CLK, Q => 
                           n24631, QN => n19923);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n6031, CK => CLK, Q => 
                           n24630, QN => n19924);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n6030, CK => CLK, Q => 
                           n24629, QN => n19925);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n6029, CK => CLK, Q => 
                           n24628, QN => n19926);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n6028, CK => CLK, Q => 
                           n24627, QN => n19927);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n6027, CK => CLK, Q => 
                           n24626, QN => n19928);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n6026, CK => CLK, Q => 
                           n24625, QN => n19929);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n6025, CK => CLK, Q => 
                           n24624, QN => n19930);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n6024, CK => CLK, Q => 
                           n24623, QN => n19931);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n6023, CK => CLK, Q => 
                           n24622, QN => n19932);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n6022, CK => CLK, Q => 
                           n24621, QN => n19933);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n6021, CK => CLK, Q => 
                           n24620, QN => n19934);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n6020, CK => CLK, Q => 
                           n24619, QN => n19935);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n6019, CK => CLK, Q => 
                           n24618, QN => n19936);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n6018, CK => CLK, Q => 
                           n24617, QN => n19937);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n6017, CK => CLK, Q => 
                           n24616, QN => n19938);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n6016, CK => CLK, Q => 
                           n24615, QN => n19939);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n6015, CK => CLK, Q => 
                           n24614, QN => n19940);
   OUT2_reg_63_inst : DFF_X1 port map( D => n5374, CK => CLK, Q => OUT2_63_port
                           , QN => n_2151);
   U18481 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n25046,
                           ZN => n23931);
   U18482 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n25244,
                           ZN => n22734);
   U18483 : NOR3_X1 port map( A1 => n25046, A2 => ADD_RD2(2), A3 => n19492, ZN 
                           => n23934);
   U18484 : NOR3_X1 port map( A1 => n25244, A2 => ADD_RD1(2), A3 => n19487, ZN 
                           => n22737);
   U18485 : BUF_X1 port map( A => n25570, Z => n25572);
   U18486 : BUF_X1 port map( A => n25570, Z => n25573);
   U18487 : BUF_X1 port map( A => n25570, Z => n25574);
   U18488 : BUF_X1 port map( A => n25571, Z => n25575);
   U18489 : BUF_X1 port map( A => n25571, Z => n25576);
   U18490 : BUF_X1 port map( A => n21479, Z => n25770);
   U18491 : BUF_X1 port map( A => n21479, Z => n25771);
   U18492 : BUF_X1 port map( A => n21479, Z => n25772);
   U18493 : BUF_X1 port map( A => n21479, Z => n25773);
   U18494 : BUF_X1 port map( A => n22798, Z => n24998);
   U18495 : BUF_X1 port map( A => n22798, Z => n24999);
   U18496 : BUF_X1 port map( A => n22798, Z => n25000);
   U18497 : BUF_X1 port map( A => n22798, Z => n25001);
   U18498 : BUF_X1 port map( A => n22798, Z => n25002);
   U18499 : BUF_X1 port map( A => n21601, Z => n25196);
   U18500 : BUF_X1 port map( A => n21601, Z => n25197);
   U18501 : BUF_X1 port map( A => n21601, Z => n25198);
   U18502 : BUF_X1 port map( A => n21601, Z => n25199);
   U18503 : BUF_X1 port map( A => n21601, Z => n25200);
   U18504 : BUF_X1 port map( A => n25595, Z => n25597);
   U18505 : BUF_X1 port map( A => n25557, Z => n25559);
   U18506 : BUF_X1 port map( A => n25467, Z => n25469);
   U18507 : BUF_X1 port map( A => n25634, Z => n25636);
   U18508 : BUF_X1 port map( A => n25441, Z => n25443);
   U18509 : BUF_X1 port map( A => n25402, Z => n25404);
   U18510 : BUF_X1 port map( A => n25480, Z => n25482);
   U18511 : BUF_X1 port map( A => n25762, Z => n25764);
   U18512 : BUF_X1 port map( A => n25454, Z => n25456);
   U18513 : BUF_X1 port map( A => n25376, Z => n25378);
   U18514 : BUF_X1 port map( A => n25531, Z => n25533);
   U18515 : BUF_X1 port map( A => n25724, Z => n25726);
   U18516 : BUF_X1 port map( A => n25647, Z => n25649);
   U18517 : BUF_X1 port map( A => n25415, Z => n25417);
   U18518 : BUF_X1 port map( A => n25389, Z => n25391);
   U18519 : BUF_X1 port map( A => n25621, Z => n25623);
   U18520 : BUF_X1 port map( A => n25544, Z => n25546);
   U18521 : BUF_X1 port map( A => n25518, Z => n25520);
   U18522 : BUF_X1 port map( A => n25737, Z => n25739);
   U18523 : BUF_X1 port map( A => n25428, Z => n25430);
   U18524 : BUF_X1 port map( A => n25493, Z => n25495);
   U18525 : BUF_X1 port map( A => n25608, Z => n25610);
   U18526 : BUF_X1 port map( A => n25660, Z => n25662);
   U18527 : BUF_X1 port map( A => n25673, Z => n25675);
   U18528 : BUF_X1 port map( A => n25698, Z => n25700);
   U18529 : BUF_X1 port map( A => n25711, Z => n25713);
   U18530 : BUF_X1 port map( A => n25595, Z => n25598);
   U18531 : BUF_X1 port map( A => n25595, Z => n25599);
   U18532 : BUF_X1 port map( A => n25596, Z => n25600);
   U18533 : BUF_X1 port map( A => n25596, Z => n25601);
   U18534 : BUF_X1 port map( A => n25557, Z => n25560);
   U18535 : BUF_X1 port map( A => n25557, Z => n25561);
   U18536 : BUF_X1 port map( A => n25558, Z => n25562);
   U18537 : BUF_X1 port map( A => n25558, Z => n25563);
   U18538 : BUF_X1 port map( A => n25467, Z => n25470);
   U18539 : BUF_X1 port map( A => n25467, Z => n25471);
   U18540 : BUF_X1 port map( A => n25468, Z => n25472);
   U18541 : BUF_X1 port map( A => n25468, Z => n25473);
   U18542 : BUF_X1 port map( A => n25634, Z => n25637);
   U18543 : BUF_X1 port map( A => n25634, Z => n25638);
   U18544 : BUF_X1 port map( A => n25635, Z => n25639);
   U18545 : BUF_X1 port map( A => n25635, Z => n25640);
   U18546 : BUF_X1 port map( A => n25441, Z => n25444);
   U18547 : BUF_X1 port map( A => n25441, Z => n25445);
   U18548 : BUF_X1 port map( A => n25442, Z => n25446);
   U18549 : BUF_X1 port map( A => n25402, Z => n25405);
   U18550 : BUF_X1 port map( A => n25402, Z => n25406);
   U18551 : BUF_X1 port map( A => n25403, Z => n25407);
   U18552 : BUF_X1 port map( A => n25442, Z => n25447);
   U18553 : BUF_X1 port map( A => n25403, Z => n25408);
   U18554 : BUF_X1 port map( A => n25480, Z => n25483);
   U18555 : BUF_X1 port map( A => n25480, Z => n25484);
   U18556 : BUF_X1 port map( A => n25481, Z => n25485);
   U18557 : BUF_X1 port map( A => n25481, Z => n25486);
   U18558 : BUF_X1 port map( A => n25762, Z => n25765);
   U18559 : BUF_X1 port map( A => n25762, Z => n25766);
   U18560 : BUF_X1 port map( A => n25763, Z => n25767);
   U18561 : BUF_X1 port map( A => n25763, Z => n25768);
   U18562 : BUF_X1 port map( A => n25454, Z => n25457);
   U18563 : BUF_X1 port map( A => n25454, Z => n25458);
   U18564 : BUF_X1 port map( A => n25455, Z => n25459);
   U18565 : BUF_X1 port map( A => n25376, Z => n25379);
   U18566 : BUF_X1 port map( A => n25376, Z => n25380);
   U18567 : BUF_X1 port map( A => n25377, Z => n25381);
   U18568 : BUF_X1 port map( A => n25455, Z => n25460);
   U18569 : BUF_X1 port map( A => n25377, Z => n25382);
   U18570 : BUF_X1 port map( A => n25531, Z => n25534);
   U18571 : BUF_X1 port map( A => n25531, Z => n25535);
   U18572 : BUF_X1 port map( A => n25532, Z => n25536);
   U18573 : BUF_X1 port map( A => n25532, Z => n25537);
   U18574 : BUF_X1 port map( A => n25724, Z => n25727);
   U18575 : BUF_X1 port map( A => n25724, Z => n25728);
   U18576 : BUF_X1 port map( A => n25725, Z => n25729);
   U18577 : BUF_X1 port map( A => n25725, Z => n25730);
   U18578 : BUF_X1 port map( A => n25647, Z => n25650);
   U18579 : BUF_X1 port map( A => n25647, Z => n25651);
   U18580 : BUF_X1 port map( A => n25648, Z => n25652);
   U18581 : BUF_X1 port map( A => n25648, Z => n25653);
   U18582 : BUF_X1 port map( A => n25415, Z => n25418);
   U18583 : BUF_X1 port map( A => n25415, Z => n25419);
   U18584 : BUF_X1 port map( A => n25416, Z => n25420);
   U18585 : BUF_X1 port map( A => n25389, Z => n25392);
   U18586 : BUF_X1 port map( A => n25389, Z => n25393);
   U18587 : BUF_X1 port map( A => n25390, Z => n25394);
   U18588 : BUF_X1 port map( A => n25621, Z => n25624);
   U18589 : BUF_X1 port map( A => n25621, Z => n25625);
   U18590 : BUF_X1 port map( A => n25622, Z => n25626);
   U18591 : BUF_X1 port map( A => n25622, Z => n25627);
   U18592 : BUF_X1 port map( A => n25544, Z => n25547);
   U18593 : BUF_X1 port map( A => n25544, Z => n25548);
   U18594 : BUF_X1 port map( A => n25545, Z => n25549);
   U18595 : BUF_X1 port map( A => n25545, Z => n25550);
   U18596 : BUF_X1 port map( A => n25518, Z => n25521);
   U18597 : BUF_X1 port map( A => n25518, Z => n25522);
   U18598 : BUF_X1 port map( A => n25519, Z => n25523);
   U18599 : BUF_X1 port map( A => n25519, Z => n25524);
   U18600 : BUF_X1 port map( A => n25416, Z => n25421);
   U18601 : BUF_X1 port map( A => n25390, Z => n25395);
   U18602 : BUF_X1 port map( A => n25737, Z => n25740);
   U18603 : BUF_X1 port map( A => n25737, Z => n25741);
   U18604 : BUF_X1 port map( A => n25738, Z => n25742);
   U18605 : BUF_X1 port map( A => n25738, Z => n25743);
   U18606 : BUF_X1 port map( A => n25428, Z => n25431);
   U18607 : BUF_X1 port map( A => n25428, Z => n25432);
   U18608 : BUF_X1 port map( A => n25429, Z => n25433);
   U18609 : BUF_X1 port map( A => n25429, Z => n25434);
   U18610 : BUF_X1 port map( A => n25493, Z => n25496);
   U18611 : BUF_X1 port map( A => n25493, Z => n25497);
   U18612 : BUF_X1 port map( A => n25494, Z => n25498);
   U18613 : BUF_X1 port map( A => n25494, Z => n25499);
   U18614 : BUF_X1 port map( A => n25608, Z => n25611);
   U18615 : BUF_X1 port map( A => n25608, Z => n25612);
   U18616 : BUF_X1 port map( A => n25609, Z => n25613);
   U18617 : BUF_X1 port map( A => n25609, Z => n25614);
   U18618 : BUF_X1 port map( A => n25660, Z => n25663);
   U18619 : BUF_X1 port map( A => n25660, Z => n25664);
   U18620 : BUF_X1 port map( A => n25661, Z => n25665);
   U18621 : BUF_X1 port map( A => n25661, Z => n25666);
   U18622 : BUF_X1 port map( A => n25673, Z => n25676);
   U18623 : BUF_X1 port map( A => n25673, Z => n25677);
   U18624 : BUF_X1 port map( A => n25674, Z => n25678);
   U18625 : BUF_X1 port map( A => n25674, Z => n25679);
   U18626 : BUF_X1 port map( A => n25698, Z => n25701);
   U18627 : BUF_X1 port map( A => n25698, Z => n25702);
   U18628 : BUF_X1 port map( A => n25699, Z => n25703);
   U18629 : BUF_X1 port map( A => n25699, Z => n25704);
   U18630 : BUF_X1 port map( A => n25711, Z => n25714);
   U18631 : BUF_X1 port map( A => n25711, Z => n25715);
   U18632 : BUF_X1 port map( A => n25712, Z => n25716);
   U18633 : BUF_X1 port map( A => n25712, Z => n25717);
   U18634 : BUF_X1 port map( A => n21478, Z => n25775);
   U18635 : BUF_X1 port map( A => n21478, Z => n25776);
   U18636 : BUF_X1 port map( A => n21478, Z => n25777);
   U18637 : BUF_X1 port map( A => n21478, Z => n25778);
   U18638 : BUF_X1 port map( A => n21478, Z => n25779);
   U18639 : BUF_X1 port map( A => n21483, Z => n25756);
   U18640 : BUF_X1 port map( A => n21483, Z => n25757);
   U18641 : BUF_X1 port map( A => n21483, Z => n25758);
   U18642 : BUF_X1 port map( A => n21483, Z => n25759);
   U18643 : BUF_X1 port map( A => n21483, Z => n25760);
   U18644 : BUF_X1 port map( A => n21555, Z => n25370);
   U18645 : BUF_X1 port map( A => n21555, Z => n25371);
   U18646 : BUF_X1 port map( A => n21555, Z => n25372);
   U18647 : BUF_X1 port map( A => n21555, Z => n25373);
   U18648 : BUF_X1 port map( A => n21555, Z => n25374);
   U18649 : BUF_X1 port map( A => n21486, Z => n25744);
   U18650 : BUF_X1 port map( A => n21486, Z => n25745);
   U18651 : BUF_X1 port map( A => n21486, Z => n25746);
   U18652 : BUF_X1 port map( A => n21486, Z => n25747);
   U18653 : BUF_X1 port map( A => n21486, Z => n25748);
   U18654 : BUF_X1 port map( A => n21516, Z => n25589);
   U18655 : BUF_X1 port map( A => n21516, Z => n25590);
   U18656 : BUF_X1 port map( A => n21516, Z => n25591);
   U18657 : BUF_X1 port map( A => n21516, Z => n25592);
   U18658 : BUF_X1 port map( A => n21516, Z => n25593);
   U18659 : BUF_X1 port map( A => n21523, Z => n25551);
   U18660 : BUF_X1 port map( A => n21523, Z => n25552);
   U18661 : BUF_X1 port map( A => n21523, Z => n25553);
   U18662 : BUF_X1 port map( A => n21523, Z => n25554);
   U18663 : BUF_X1 port map( A => n21523, Z => n25555);
   U18664 : BUF_X1 port map( A => n21539, Z => n25461);
   U18665 : BUF_X1 port map( A => n21539, Z => n25462);
   U18666 : BUF_X1 port map( A => n21539, Z => n25463);
   U18667 : BUF_X1 port map( A => n21539, Z => n25464);
   U18668 : BUF_X1 port map( A => n21539, Z => n25465);
   U18669 : BUF_X1 port map( A => n21509, Z => n25628);
   U18670 : BUF_X1 port map( A => n21509, Z => n25629);
   U18671 : BUF_X1 port map( A => n21509, Z => n25630);
   U18672 : BUF_X1 port map( A => n21509, Z => n25631);
   U18673 : BUF_X1 port map( A => n21509, Z => n25632);
   U18674 : BUF_X1 port map( A => n21544, Z => n25435);
   U18675 : BUF_X1 port map( A => n21544, Z => n25436);
   U18676 : BUF_X1 port map( A => n21544, Z => n25437);
   U18677 : BUF_X1 port map( A => n21544, Z => n25438);
   U18678 : BUF_X1 port map( A => n21544, Z => n25439);
   U18679 : BUF_X1 port map( A => n21551, Z => n25396);
   U18680 : BUF_X1 port map( A => n21551, Z => n25397);
   U18681 : BUF_X1 port map( A => n21551, Z => n25398);
   U18682 : BUF_X1 port map( A => n21551, Z => n25399);
   U18683 : BUF_X1 port map( A => n21551, Z => n25400);
   U18684 : BUF_X1 port map( A => n21537, Z => n25474);
   U18685 : BUF_X1 port map( A => n21537, Z => n25475);
   U18686 : BUF_X1 port map( A => n21537, Z => n25476);
   U18687 : BUF_X1 port map( A => n21537, Z => n25477);
   U18688 : BUF_X1 port map( A => n21537, Z => n25478);
   U18689 : BUF_X1 port map( A => n21520, Z => n25564);
   U18690 : BUF_X1 port map( A => n21520, Z => n25565);
   U18691 : BUF_X1 port map( A => n21520, Z => n25566);
   U18692 : BUF_X1 port map( A => n21520, Z => n25567);
   U18693 : BUF_X1 port map( A => n21520, Z => n25568);
   U18694 : BUF_X1 port map( A => n21542, Z => n25448);
   U18695 : BUF_X1 port map( A => n21542, Z => n25449);
   U18696 : BUF_X1 port map( A => n21542, Z => n25450);
   U18697 : BUF_X1 port map( A => n21542, Z => n25451);
   U18698 : BUF_X1 port map( A => n21542, Z => n25452);
   U18699 : BUF_X1 port map( A => n21527, Z => n25525);
   U18700 : BUF_X1 port map( A => n21527, Z => n25526);
   U18701 : BUF_X1 port map( A => n21527, Z => n25527);
   U18702 : BUF_X1 port map( A => n21527, Z => n25528);
   U18703 : BUF_X1 port map( A => n21527, Z => n25529);
   U18704 : BUF_X1 port map( A => n21493, Z => n25718);
   U18705 : BUF_X1 port map( A => n21493, Z => n25719);
   U18706 : BUF_X1 port map( A => n21493, Z => n25720);
   U18707 : BUF_X1 port map( A => n21493, Z => n25721);
   U18708 : BUF_X1 port map( A => n21493, Z => n25722);
   U18709 : BUF_X1 port map( A => n21507, Z => n25641);
   U18710 : BUF_X1 port map( A => n21507, Z => n25642);
   U18711 : BUF_X1 port map( A => n21507, Z => n25643);
   U18712 : BUF_X1 port map( A => n21507, Z => n25644);
   U18713 : BUF_X1 port map( A => n21507, Z => n25645);
   U18714 : BUF_X1 port map( A => n21548, Z => n25409);
   U18715 : BUF_X1 port map( A => n21548, Z => n25410);
   U18716 : BUF_X1 port map( A => n21548, Z => n25411);
   U18717 : BUF_X1 port map( A => n21548, Z => n25412);
   U18718 : BUF_X1 port map( A => n21548, Z => n25413);
   U18719 : BUF_X1 port map( A => n21553, Z => n25383);
   U18720 : BUF_X1 port map( A => n21553, Z => n25384);
   U18721 : BUF_X1 port map( A => n21553, Z => n25385);
   U18722 : BUF_X1 port map( A => n21553, Z => n25386);
   U18723 : BUF_X1 port map( A => n21553, Z => n25387);
   U18724 : BUF_X1 port map( A => n21511, Z => n25615);
   U18725 : BUF_X1 port map( A => n21511, Z => n25616);
   U18726 : BUF_X1 port map( A => n21511, Z => n25617);
   U18727 : BUF_X1 port map( A => n21511, Z => n25618);
   U18728 : BUF_X1 port map( A => n21511, Z => n25619);
   U18729 : BUF_X1 port map( A => n21525, Z => n25538);
   U18730 : BUF_X1 port map( A => n21525, Z => n25539);
   U18731 : BUF_X1 port map( A => n21525, Z => n25540);
   U18732 : BUF_X1 port map( A => n21525, Z => n25541);
   U18733 : BUF_X1 port map( A => n21525, Z => n25542);
   U18734 : BUF_X1 port map( A => n21530, Z => n25512);
   U18735 : BUF_X1 port map( A => n21530, Z => n25513);
   U18736 : BUF_X1 port map( A => n21530, Z => n25514);
   U18737 : BUF_X1 port map( A => n21530, Z => n25515);
   U18738 : BUF_X1 port map( A => n21530, Z => n25516);
   U18739 : BUF_X1 port map( A => n21489, Z => n25731);
   U18740 : BUF_X1 port map( A => n21489, Z => n25732);
   U18741 : BUF_X1 port map( A => n21489, Z => n25733);
   U18742 : BUF_X1 port map( A => n21489, Z => n25734);
   U18743 : BUF_X1 port map( A => n21489, Z => n25735);
   U18744 : BUF_X1 port map( A => n21546, Z => n25422);
   U18745 : BUF_X1 port map( A => n21546, Z => n25423);
   U18746 : BUF_X1 port map( A => n21546, Z => n25424);
   U18747 : BUF_X1 port map( A => n21546, Z => n25425);
   U18748 : BUF_X1 port map( A => n21546, Z => n25426);
   U18749 : BUF_X1 port map( A => n21518, Z => n25577);
   U18750 : BUF_X1 port map( A => n21518, Z => n25578);
   U18751 : BUF_X1 port map( A => n21518, Z => n25579);
   U18752 : BUF_X1 port map( A => n21518, Z => n25580);
   U18753 : BUF_X1 port map( A => n21518, Z => n25581);
   U18754 : BUF_X1 port map( A => n21533, Z => n25500);
   U18755 : BUF_X1 port map( A => n21533, Z => n25501);
   U18756 : BUF_X1 port map( A => n21533, Z => n25502);
   U18757 : BUF_X1 port map( A => n21533, Z => n25503);
   U18758 : BUF_X1 port map( A => n21533, Z => n25504);
   U18759 : BUF_X1 port map( A => n21500, Z => n25680);
   U18760 : BUF_X1 port map( A => n21500, Z => n25681);
   U18761 : BUF_X1 port map( A => n21500, Z => n25682);
   U18762 : BUF_X1 port map( A => n21500, Z => n25683);
   U18763 : BUF_X1 port map( A => n21500, Z => n25684);
   U18764 : BUF_X1 port map( A => n21535, Z => n25487);
   U18765 : BUF_X1 port map( A => n21535, Z => n25488);
   U18766 : BUF_X1 port map( A => n21535, Z => n25489);
   U18767 : BUF_X1 port map( A => n21535, Z => n25490);
   U18768 : BUF_X1 port map( A => n21535, Z => n25491);
   U18769 : BUF_X1 port map( A => n21514, Z => n25602);
   U18770 : BUF_X1 port map( A => n21514, Z => n25603);
   U18771 : BUF_X1 port map( A => n21514, Z => n25604);
   U18772 : BUF_X1 port map( A => n21514, Z => n25605);
   U18773 : BUF_X1 port map( A => n21514, Z => n25606);
   U18774 : BUF_X1 port map( A => n21505, Z => n25654);
   U18775 : BUF_X1 port map( A => n21505, Z => n25655);
   U18776 : BUF_X1 port map( A => n21505, Z => n25656);
   U18777 : BUF_X1 port map( A => n21505, Z => n25657);
   U18778 : BUF_X1 port map( A => n21505, Z => n25658);
   U18779 : BUF_X1 port map( A => n21502, Z => n25667);
   U18780 : BUF_X1 port map( A => n21502, Z => n25668);
   U18781 : BUF_X1 port map( A => n21502, Z => n25669);
   U18782 : BUF_X1 port map( A => n21502, Z => n25670);
   U18783 : BUF_X1 port map( A => n21502, Z => n25671);
   U18784 : BUF_X1 port map( A => n21498, Z => n25692);
   U18785 : BUF_X1 port map( A => n21498, Z => n25693);
   U18786 : BUF_X1 port map( A => n21498, Z => n25694);
   U18787 : BUF_X1 port map( A => n21498, Z => n25695);
   U18788 : BUF_X1 port map( A => n21498, Z => n25696);
   U18789 : BUF_X1 port map( A => n21496, Z => n25705);
   U18790 : BUF_X1 port map( A => n21496, Z => n25706);
   U18791 : BUF_X1 port map( A => n21496, Z => n25707);
   U18792 : BUF_X1 port map( A => n21496, Z => n25708);
   U18793 : BUF_X1 port map( A => n21496, Z => n25709);
   U18794 : BUF_X1 port map( A => n21479, Z => n25769);
   U18795 : BUF_X1 port map( A => n21519, Z => n25570);
   U18796 : BUF_X1 port map( A => n21519, Z => n25571);
   U18797 : OAI21_X1 port map( B1 => n21480, B2 => n21481, A => n25973, ZN => 
                           n21478);
   U18798 : BUF_X1 port map( A => n22777, Z => n25082);
   U18799 : BUF_X1 port map( A => n22777, Z => n25083);
   U18800 : BUF_X1 port map( A => n22777, Z => n25084);
   U18801 : BUF_X1 port map( A => n22777, Z => n25085);
   U18802 : BUF_X1 port map( A => n22777, Z => n25086);
   U18803 : BUF_X1 port map( A => n21580, Z => n25280);
   U18804 : BUF_X1 port map( A => n21580, Z => n25281);
   U18805 : BUF_X1 port map( A => n21580, Z => n25282);
   U18806 : BUF_X1 port map( A => n21580, Z => n25283);
   U18807 : BUF_X1 port map( A => n21580, Z => n25284);
   U18808 : BUF_X1 port map( A => n22787, Z => n25052);
   U18809 : BUF_X1 port map( A => n22787, Z => n25053);
   U18810 : BUF_X1 port map( A => n22787, Z => n25054);
   U18811 : BUF_X1 port map( A => n22787, Z => n25055);
   U18812 : BUF_X1 port map( A => n22787, Z => n25056);
   U18813 : BUF_X1 port map( A => n21590, Z => n25250);
   U18814 : BUF_X1 port map( A => n21590, Z => n25251);
   U18815 : BUF_X1 port map( A => n21590, Z => n25252);
   U18816 : BUF_X1 port map( A => n21590, Z => n25253);
   U18817 : BUF_X1 port map( A => n21590, Z => n25254);
   U18818 : BUF_X1 port map( A => n22767, Z => n25130);
   U18819 : BUF_X1 port map( A => n22767, Z => n25131);
   U18820 : BUF_X1 port map( A => n22767, Z => n25132);
   U18821 : BUF_X1 port map( A => n22767, Z => n25133);
   U18822 : BUF_X1 port map( A => n22767, Z => n25134);
   U18823 : BUF_X1 port map( A => n21570, Z => n25328);
   U18824 : BUF_X1 port map( A => n21570, Z => n25329);
   U18825 : BUF_X1 port map( A => n21570, Z => n25330);
   U18826 : BUF_X1 port map( A => n21570, Z => n25331);
   U18827 : BUF_X1 port map( A => n21570, Z => n25332);
   U18828 : BUF_X1 port map( A => n22762, Z => n25154);
   U18829 : BUF_X1 port map( A => n22772, Z => n25106);
   U18830 : BUF_X1 port map( A => n22792, Z => n25028);
   U18831 : BUF_X1 port map( A => n22797, Z => n25004);
   U18832 : BUF_X1 port map( A => n22802, Z => n24980);
   U18833 : BUF_X1 port map( A => n22762, Z => n25155);
   U18834 : BUF_X1 port map( A => n22772, Z => n25107);
   U18835 : BUF_X1 port map( A => n22792, Z => n25029);
   U18836 : BUF_X1 port map( A => n22797, Z => n25005);
   U18837 : BUF_X1 port map( A => n22802, Z => n24981);
   U18838 : BUF_X1 port map( A => n22762, Z => n25156);
   U18839 : BUF_X1 port map( A => n22772, Z => n25108);
   U18840 : BUF_X1 port map( A => n22792, Z => n25030);
   U18841 : BUF_X1 port map( A => n22797, Z => n25006);
   U18842 : BUF_X1 port map( A => n22802, Z => n24982);
   U18843 : BUF_X1 port map( A => n22762, Z => n25157);
   U18844 : BUF_X1 port map( A => n22772, Z => n25109);
   U18845 : BUF_X1 port map( A => n22792, Z => n25031);
   U18846 : BUF_X1 port map( A => n22797, Z => n25007);
   U18847 : BUF_X1 port map( A => n22802, Z => n24983);
   U18848 : BUF_X1 port map( A => n22762, Z => n25158);
   U18849 : BUF_X1 port map( A => n22772, Z => n25110);
   U18850 : BUF_X1 port map( A => n22792, Z => n25032);
   U18851 : BUF_X1 port map( A => n22797, Z => n25008);
   U18852 : BUF_X1 port map( A => n22802, Z => n24984);
   U18853 : BUF_X1 port map( A => n21565, Z => n25352);
   U18854 : BUF_X1 port map( A => n21575, Z => n25304);
   U18855 : BUF_X1 port map( A => n21595, Z => n25226);
   U18856 : BUF_X1 port map( A => n21600, Z => n25202);
   U18857 : BUF_X1 port map( A => n21605, Z => n25178);
   U18858 : BUF_X1 port map( A => n21565, Z => n25353);
   U18859 : BUF_X1 port map( A => n21575, Z => n25305);
   U18860 : BUF_X1 port map( A => n21595, Z => n25227);
   U18861 : BUF_X1 port map( A => n21600, Z => n25203);
   U18862 : BUF_X1 port map( A => n21605, Z => n25179);
   U18863 : BUF_X1 port map( A => n21565, Z => n25354);
   U18864 : BUF_X1 port map( A => n21575, Z => n25306);
   U18865 : BUF_X1 port map( A => n21595, Z => n25228);
   U18866 : BUF_X1 port map( A => n21600, Z => n25204);
   U18867 : BUF_X1 port map( A => n21605, Z => n25180);
   U18868 : BUF_X1 port map( A => n21565, Z => n25355);
   U18869 : BUF_X1 port map( A => n21575, Z => n25307);
   U18870 : BUF_X1 port map( A => n21595, Z => n25229);
   U18871 : BUF_X1 port map( A => n21600, Z => n25205);
   U18872 : BUF_X1 port map( A => n21605, Z => n25181);
   U18873 : BUF_X1 port map( A => n21565, Z => n25356);
   U18874 : BUF_X1 port map( A => n21575, Z => n25308);
   U18875 : BUF_X1 port map( A => n21595, Z => n25230);
   U18876 : BUF_X1 port map( A => n21600, Z => n25206);
   U18877 : BUF_X1 port map( A => n21605, Z => n25182);
   U18878 : BUF_X1 port map( A => n22759, Z => n25167);
   U18879 : BUF_X1 port map( A => n22769, Z => n25119);
   U18880 : BUF_X1 port map( A => n22764, Z => n25143);
   U18881 : BUF_X1 port map( A => n22789, Z => n25041);
   U18882 : BUF_X1 port map( A => n22759, Z => n25168);
   U18883 : BUF_X1 port map( A => n22769, Z => n25120);
   U18884 : BUF_X1 port map( A => n22764, Z => n25144);
   U18885 : BUF_X1 port map( A => n22789, Z => n25042);
   U18886 : BUF_X1 port map( A => n22759, Z => n25169);
   U18887 : BUF_X1 port map( A => n22769, Z => n25121);
   U18888 : BUF_X1 port map( A => n22764, Z => n25145);
   U18889 : BUF_X1 port map( A => n22789, Z => n25043);
   U18890 : BUF_X1 port map( A => n22759, Z => n25170);
   U18891 : BUF_X1 port map( A => n22769, Z => n25122);
   U18892 : BUF_X1 port map( A => n22764, Z => n25146);
   U18893 : BUF_X1 port map( A => n22789, Z => n25044);
   U18894 : BUF_X1 port map( A => n21562, Z => n25365);
   U18895 : BUF_X1 port map( A => n21572, Z => n25317);
   U18896 : BUF_X1 port map( A => n21567, Z => n25341);
   U18897 : BUF_X1 port map( A => n21592, Z => n25239);
   U18898 : BUF_X1 port map( A => n21562, Z => n25366);
   U18899 : BUF_X1 port map( A => n21572, Z => n25318);
   U18900 : BUF_X1 port map( A => n21567, Z => n25342);
   U18901 : BUF_X1 port map( A => n21592, Z => n25240);
   U18902 : BUF_X1 port map( A => n21562, Z => n25367);
   U18903 : BUF_X1 port map( A => n21572, Z => n25319);
   U18904 : BUF_X1 port map( A => n21567, Z => n25343);
   U18905 : BUF_X1 port map( A => n21592, Z => n25241);
   U18906 : BUF_X1 port map( A => n21562, Z => n25368);
   U18907 : BUF_X1 port map( A => n21572, Z => n25320);
   U18908 : BUF_X1 port map( A => n21567, Z => n25344);
   U18909 : BUF_X1 port map( A => n21592, Z => n25242);
   U18910 : BUF_X1 port map( A => n22774, Z => n25095);
   U18911 : BUF_X1 port map( A => n22794, Z => n25017);
   U18912 : BUF_X1 port map( A => n22774, Z => n25096);
   U18913 : BUF_X1 port map( A => n22774, Z => n25097);
   U18914 : BUF_X1 port map( A => n22799, Z => n24993);
   U18915 : BUF_X1 port map( A => n22794, Z => n25018);
   U18916 : BUF_X1 port map( A => n22794, Z => n25019);
   U18917 : BUF_X1 port map( A => n22774, Z => n25098);
   U18918 : BUF_X1 port map( A => n22794, Z => n25020);
   U18919 : BUF_X1 port map( A => n21577, Z => n25293);
   U18920 : BUF_X1 port map( A => n21577, Z => n25294);
   U18921 : BUF_X1 port map( A => n21577, Z => n25296);
   U18922 : BUF_X1 port map( A => n22784, Z => n25065);
   U18923 : BUF_X1 port map( A => n22784, Z => n25066);
   U18924 : BUF_X1 port map( A => n22799, Z => n24994);
   U18925 : BUF_X1 port map( A => n22784, Z => n25067);
   U18926 : BUF_X1 port map( A => n22799, Z => n24995);
   U18927 : BUF_X1 port map( A => n22784, Z => n25068);
   U18928 : BUF_X1 port map( A => n22799, Z => n24996);
   U18929 : BUF_X1 port map( A => n21587, Z => n25263);
   U18930 : BUF_X1 port map( A => n21597, Z => n25215);
   U18931 : BUF_X1 port map( A => n21577, Z => n25295);
   U18932 : BUF_X1 port map( A => n21602, Z => n25191);
   U18933 : BUF_X1 port map( A => n21587, Z => n25264);
   U18934 : BUF_X1 port map( A => n21597, Z => n25216);
   U18935 : BUF_X1 port map( A => n21602, Z => n25192);
   U18936 : BUF_X1 port map( A => n21587, Z => n25265);
   U18937 : BUF_X1 port map( A => n21597, Z => n25217);
   U18938 : BUF_X1 port map( A => n21602, Z => n25193);
   U18939 : BUF_X1 port map( A => n21587, Z => n25266);
   U18940 : BUF_X1 port map( A => n21597, Z => n25218);
   U18941 : BUF_X1 port map( A => n21602, Z => n25194);
   U18942 : BUF_X1 port map( A => n22778, Z => n25076);
   U18943 : BUF_X1 port map( A => n22778, Z => n25077);
   U18944 : BUF_X1 port map( A => n22778, Z => n25078);
   U18945 : BUF_X1 port map( A => n22778, Z => n25079);
   U18946 : BUF_X1 port map( A => n22778, Z => n25080);
   U18947 : BUF_X1 port map( A => n21581, Z => n25274);
   U18948 : BUF_X1 port map( A => n21581, Z => n25275);
   U18949 : BUF_X1 port map( A => n21581, Z => n25276);
   U18950 : BUF_X1 port map( A => n21581, Z => n25277);
   U18951 : BUF_X1 port map( A => n21581, Z => n25278);
   U18952 : BUF_X1 port map( A => n22773, Z => n25100);
   U18953 : BUF_X1 port map( A => n22768, Z => n25124);
   U18954 : BUF_X1 port map( A => n22793, Z => n25022);
   U18955 : BUF_X1 port map( A => n22803, Z => n24974);
   U18956 : BUF_X1 port map( A => n22773, Z => n25101);
   U18957 : BUF_X1 port map( A => n22768, Z => n25125);
   U18958 : BUF_X1 port map( A => n22793, Z => n25023);
   U18959 : BUF_X1 port map( A => n22803, Z => n24975);
   U18960 : BUF_X1 port map( A => n22773, Z => n25102);
   U18961 : BUF_X1 port map( A => n22768, Z => n25126);
   U18962 : BUF_X1 port map( A => n22793, Z => n25024);
   U18963 : BUF_X1 port map( A => n22803, Z => n24976);
   U18964 : BUF_X1 port map( A => n22773, Z => n25103);
   U18965 : BUF_X1 port map( A => n22768, Z => n25127);
   U18966 : BUF_X1 port map( A => n22793, Z => n25025);
   U18967 : BUF_X1 port map( A => n22803, Z => n24977);
   U18968 : BUF_X1 port map( A => n22773, Z => n25104);
   U18969 : BUF_X1 port map( A => n22768, Z => n25128);
   U18970 : BUF_X1 port map( A => n22793, Z => n25026);
   U18971 : BUF_X1 port map( A => n22803, Z => n24978);
   U18972 : BUF_X1 port map( A => n21576, Z => n25298);
   U18973 : BUF_X1 port map( A => n21571, Z => n25322);
   U18974 : BUF_X1 port map( A => n21596, Z => n25220);
   U18975 : BUF_X1 port map( A => n21606, Z => n25172);
   U18976 : BUF_X1 port map( A => n21576, Z => n25299);
   U18977 : BUF_X1 port map( A => n21571, Z => n25323);
   U18978 : BUF_X1 port map( A => n21596, Z => n25221);
   U18979 : BUF_X1 port map( A => n21606, Z => n25173);
   U18980 : BUF_X1 port map( A => n21576, Z => n25300);
   U18981 : BUF_X1 port map( A => n21571, Z => n25324);
   U18982 : BUF_X1 port map( A => n21596, Z => n25222);
   U18983 : BUF_X1 port map( A => n21606, Z => n25174);
   U18984 : BUF_X1 port map( A => n21576, Z => n25301);
   U18985 : BUF_X1 port map( A => n21571, Z => n25325);
   U18986 : BUF_X1 port map( A => n21596, Z => n25223);
   U18987 : BUF_X1 port map( A => n21606, Z => n25175);
   U18988 : BUF_X1 port map( A => n21576, Z => n25302);
   U18989 : BUF_X1 port map( A => n21571, Z => n25326);
   U18990 : BUF_X1 port map( A => n21596, Z => n25224);
   U18991 : BUF_X1 port map( A => n21606, Z => n25176);
   U18992 : BUF_X1 port map( A => n22763, Z => n25148);
   U18993 : BUF_X1 port map( A => n22763, Z => n25149);
   U18994 : BUF_X1 port map( A => n22763, Z => n25150);
   U18995 : BUF_X1 port map( A => n22763, Z => n25151);
   U18996 : BUF_X1 port map( A => n22763, Z => n25152);
   U18997 : BUF_X1 port map( A => n21566, Z => n25346);
   U18998 : BUF_X1 port map( A => n21566, Z => n25347);
   U18999 : BUF_X1 port map( A => n21566, Z => n25348);
   U19000 : BUF_X1 port map( A => n21566, Z => n25349);
   U19001 : BUF_X1 port map( A => n21566, Z => n25350);
   U19002 : BUF_X1 port map( A => n22779, Z => n25070);
   U19003 : BUF_X1 port map( A => n22779, Z => n25071);
   U19004 : BUF_X1 port map( A => n22779, Z => n25072);
   U19005 : BUF_X1 port map( A => n22779, Z => n25073);
   U19006 : BUF_X1 port map( A => n22779, Z => n25074);
   U19007 : BUF_X1 port map( A => n21582, Z => n25268);
   U19008 : BUF_X1 port map( A => n21582, Z => n25269);
   U19009 : BUF_X1 port map( A => n21582, Z => n25270);
   U19010 : BUF_X1 port map( A => n21582, Z => n25271);
   U19011 : BUF_X1 port map( A => n21582, Z => n25272);
   U19012 : NAND2_X1 port map( A1 => n25978, A2 => n25764, ZN => n21483);
   U19013 : NAND2_X1 port map( A1 => n25978, A2 => n25378, ZN => n21555);
   U19014 : NAND2_X1 port map( A1 => n25978, A2 => n25750, ZN => n21486);
   U19015 : BUF_X1 port map( A => n21517, Z => n25583);
   U19016 : BUF_X1 port map( A => n21532, Z => n25506);
   U19017 : BUF_X1 port map( A => n21485, Z => n25750);
   U19018 : BUF_X1 port map( A => n21499, Z => n25686);
   U19019 : BUF_X1 port map( A => n21517, Z => n25584);
   U19020 : BUF_X1 port map( A => n21517, Z => n25585);
   U19021 : BUF_X1 port map( A => n21517, Z => n25586);
   U19022 : BUF_X1 port map( A => n21517, Z => n25587);
   U19023 : BUF_X1 port map( A => n21532, Z => n25507);
   U19024 : BUF_X1 port map( A => n21532, Z => n25508);
   U19025 : BUF_X1 port map( A => n21532, Z => n25509);
   U19026 : BUF_X1 port map( A => n21532, Z => n25510);
   U19027 : BUF_X1 port map( A => n21485, Z => n25751);
   U19028 : BUF_X1 port map( A => n21485, Z => n25752);
   U19029 : BUF_X1 port map( A => n21485, Z => n25753);
   U19030 : BUF_X1 port map( A => n21485, Z => n25754);
   U19031 : BUF_X1 port map( A => n21499, Z => n25687);
   U19032 : BUF_X1 port map( A => n21499, Z => n25688);
   U19033 : BUF_X1 port map( A => n21499, Z => n25689);
   U19034 : BUF_X1 port map( A => n21499, Z => n25690);
   U19035 : NAND2_X1 port map( A1 => n25975, A2 => n25546, ZN => n21525);
   U19036 : NAND2_X1 port map( A1 => n25975, A2 => n25520, ZN => n21530);
   U19037 : NAND2_X1 port map( A1 => n25975, A2 => n25506, ZN => n21533);
   U19038 : NAND2_X1 port map( A1 => n25975, A2 => n25495, ZN => n21535);
   U19039 : NAND2_X1 port map( A1 => n25976, A2 => n25597, ZN => n21516);
   U19040 : NAND2_X1 port map( A1 => n25976, A2 => n25559, ZN => n21523);
   U19041 : NAND2_X1 port map( A1 => n25976, A2 => n25469, ZN => n21539);
   U19042 : NAND2_X1 port map( A1 => n25976, A2 => n25636, ZN => n21509);
   U19043 : NAND2_X1 port map( A1 => n25976, A2 => n25443, ZN => n21544);
   U19044 : NAND2_X1 port map( A1 => n25977, A2 => n25404, ZN => n21551);
   U19045 : NAND2_X1 port map( A1 => n25976, A2 => n25482, ZN => n21537);
   U19046 : NAND2_X1 port map( A1 => n25976, A2 => n25572, ZN => n21520);
   U19047 : NAND2_X1 port map( A1 => n25977, A2 => n25456, ZN => n21542);
   U19048 : NAND2_X1 port map( A1 => n25976, A2 => n25533, ZN => n21527);
   U19049 : NAND2_X1 port map( A1 => n25977, A2 => n25726, ZN => n21493);
   U19050 : NAND2_X1 port map( A1 => n25976, A2 => n25649, ZN => n21507);
   U19051 : NAND2_X1 port map( A1 => n25976, A2 => n25623, ZN => n21511);
   U19052 : NAND2_X1 port map( A1 => n25977, A2 => n25417, ZN => n21548);
   U19053 : NAND2_X1 port map( A1 => n25977, A2 => n25391, ZN => n21553);
   U19054 : NAND2_X1 port map( A1 => n25977, A2 => n25739, ZN => n21489);
   U19055 : NAND2_X1 port map( A1 => n25977, A2 => n25430, ZN => n21546);
   U19056 : NAND2_X1 port map( A1 => n25976, A2 => n25583, ZN => n21518);
   U19057 : NAND2_X1 port map( A1 => n25977, A2 => n25686, ZN => n21500);
   U19058 : NAND2_X1 port map( A1 => n25976, A2 => n25610, ZN => n21514);
   U19059 : NAND2_X1 port map( A1 => n25977, A2 => n25662, ZN => n21505);
   U19060 : NAND2_X1 port map( A1 => n25977, A2 => n25675, ZN => n21502);
   U19061 : NAND2_X1 port map( A1 => n25977, A2 => n25700, ZN => n21498);
   U19062 : NAND2_X1 port map( A1 => n25977, A2 => n25713, ZN => n21496);
   U19063 : BUF_X1 port map( A => n22775, Z => n25088);
   U19064 : BUF_X1 port map( A => n22760, Z => n25160);
   U19065 : BUF_X1 port map( A => n22765, Z => n25136);
   U19066 : BUF_X1 port map( A => n22795, Z => n25010);
   U19067 : BUF_X1 port map( A => n22775, Z => n25089);
   U19068 : BUF_X1 port map( A => n22760, Z => n25161);
   U19069 : BUF_X1 port map( A => n22765, Z => n25137);
   U19070 : BUF_X1 port map( A => n22795, Z => n25011);
   U19071 : BUF_X1 port map( A => n22760, Z => n25162);
   U19072 : BUF_X1 port map( A => n22795, Z => n25012);
   U19073 : BUF_X1 port map( A => n22785, Z => n25059);
   U19074 : BUF_X1 port map( A => n22775, Z => n25090);
   U19075 : BUF_X1 port map( A => n22765, Z => n25138);
   U19076 : BUF_X1 port map( A => n22775, Z => n25091);
   U19077 : BUF_X1 port map( A => n22760, Z => n25163);
   U19078 : BUF_X1 port map( A => n22765, Z => n25139);
   U19079 : BUF_X1 port map( A => n22795, Z => n25013);
   U19080 : BUF_X1 port map( A => n22765, Z => n25140);
   U19081 : BUF_X1 port map( A => n22795, Z => n25014);
   U19082 : BUF_X1 port map( A => n21578, Z => n25286);
   U19083 : BUF_X1 port map( A => n21563, Z => n25358);
   U19084 : BUF_X1 port map( A => n21568, Z => n25334);
   U19085 : BUF_X1 port map( A => n21598, Z => n25208);
   U19086 : BUF_X1 port map( A => n21563, Z => n25359);
   U19087 : BUF_X1 port map( A => n21568, Z => n25335);
   U19088 : BUF_X1 port map( A => n21598, Z => n25209);
   U19089 : BUF_X1 port map( A => n21563, Z => n25360);
   U19090 : BUF_X1 port map( A => n21568, Z => n25336);
   U19091 : BUF_X1 port map( A => n21598, Z => n25210);
   U19092 : BUF_X1 port map( A => n21563, Z => n25361);
   U19093 : BUF_X1 port map( A => n21598, Z => n25211);
   U19094 : BUF_X1 port map( A => n21563, Z => n25362);
   U19095 : BUF_X1 port map( A => n21568, Z => n25338);
   U19096 : BUF_X1 port map( A => n21598, Z => n25212);
   U19097 : BUF_X1 port map( A => n22790, Z => n25034);
   U19098 : BUF_X1 port map( A => n22785, Z => n25058);
   U19099 : BUF_X1 port map( A => n22790, Z => n25035);
   U19100 : BUF_X1 port map( A => n22785, Z => n25060);
   U19101 : BUF_X1 port map( A => n22790, Z => n25037);
   U19102 : BUF_X1 port map( A => n22785, Z => n25061);
   U19103 : BUF_X1 port map( A => n22775, Z => n25092);
   U19104 : BUF_X1 port map( A => n22760, Z => n25164);
   U19105 : BUF_X1 port map( A => n22790, Z => n25038);
   U19106 : BUF_X1 port map( A => n22785, Z => n25062);
   U19107 : BUF_X1 port map( A => n21593, Z => n25232);
   U19108 : BUF_X1 port map( A => n21588, Z => n25256);
   U19109 : BUF_X1 port map( A => n21578, Z => n25287);
   U19110 : BUF_X1 port map( A => n21568, Z => n25337);
   U19111 : BUF_X1 port map( A => n22790, Z => n25036);
   U19112 : BUF_X1 port map( A => n21593, Z => n25233);
   U19113 : BUF_X1 port map( A => n21588, Z => n25257);
   U19114 : BUF_X1 port map( A => n21578, Z => n25288);
   U19115 : BUF_X1 port map( A => n21593, Z => n25234);
   U19116 : BUF_X1 port map( A => n21588, Z => n25258);
   U19117 : BUF_X1 port map( A => n21578, Z => n25289);
   U19118 : BUF_X1 port map( A => n21593, Z => n25235);
   U19119 : BUF_X1 port map( A => n21588, Z => n25259);
   U19120 : BUF_X1 port map( A => n21578, Z => n25290);
   U19121 : BUF_X1 port map( A => n21593, Z => n25236);
   U19122 : BUF_X1 port map( A => n21588, Z => n25260);
   U19123 : BUF_X1 port map( A => n22770, Z => n25112);
   U19124 : BUF_X1 port map( A => n22800, Z => n24986);
   U19125 : BUF_X1 port map( A => n22770, Z => n25113);
   U19126 : BUF_X1 port map( A => n22800, Z => n24987);
   U19127 : BUF_X1 port map( A => n22770, Z => n25114);
   U19128 : BUF_X1 port map( A => n22800, Z => n24988);
   U19129 : BUF_X1 port map( A => n22770, Z => n25115);
   U19130 : BUF_X1 port map( A => n22800, Z => n24989);
   U19131 : BUF_X1 port map( A => n22770, Z => n25116);
   U19132 : BUF_X1 port map( A => n22800, Z => n24990);
   U19133 : BUF_X1 port map( A => n21573, Z => n25310);
   U19134 : BUF_X1 port map( A => n21603, Z => n25184);
   U19135 : BUF_X1 port map( A => n21573, Z => n25311);
   U19136 : BUF_X1 port map( A => n21603, Z => n25185);
   U19137 : BUF_X1 port map( A => n21573, Z => n25312);
   U19138 : BUF_X1 port map( A => n21603, Z => n25186);
   U19139 : BUF_X1 port map( A => n21573, Z => n25313);
   U19140 : BUF_X1 port map( A => n21603, Z => n25187);
   U19141 : BUF_X1 port map( A => n21573, Z => n25314);
   U19142 : BUF_X1 port map( A => n21603, Z => n25188);
   U19143 : BUF_X1 port map( A => n22759, Z => n25166);
   U19144 : BUF_X1 port map( A => n22764, Z => n25142);
   U19145 : BUF_X1 port map( A => n22789, Z => n25040);
   U19146 : BUF_X1 port map( A => n21562, Z => n25364);
   U19147 : BUF_X1 port map( A => n21567, Z => n25340);
   U19148 : BUF_X1 port map( A => n21592, Z => n25238);
   U19149 : BUF_X1 port map( A => n22769, Z => n25118);
   U19150 : BUF_X1 port map( A => n21572, Z => n25316);
   U19151 : BUF_X1 port map( A => n22774, Z => n25094);
   U19152 : BUF_X1 port map( A => n22794, Z => n25016);
   U19153 : BUF_X1 port map( A => n21577, Z => n25292);
   U19154 : BUF_X1 port map( A => n21597, Z => n25214);
   U19155 : BUF_X1 port map( A => n22784, Z => n25064);
   U19156 : BUF_X1 port map( A => n22799, Z => n24992);
   U19157 : BUF_X1 port map( A => n21587, Z => n25262);
   U19158 : BUF_X1 port map( A => n21602, Z => n25190);
   U19159 : NAND2_X1 port map( A1 => n25978, A2 => n25775, ZN => n21479);
   U19160 : OAI21_X1 port map( B1 => n21481, B2 => n21521, A => n25974, ZN => 
                           n21519);
   U19161 : AND2_X1 port map( A1 => n23946, A2 => n23928, ZN => n22798);
   U19162 : AND2_X1 port map( A1 => n22749, A2 => n22731, ZN => n21601);
   U19163 : BUF_X1 port map( A => n21482, Z => n25762);
   U19164 : BUF_X1 port map( A => n21488, Z => n25737);
   U19165 : BUF_X1 port map( A => n21515, Z => n25595);
   U19166 : BUF_X1 port map( A => n21522, Z => n25557);
   U19167 : BUF_X1 port map( A => n21538, Z => n25467);
   U19168 : BUF_X1 port map( A => n21508, Z => n25634);
   U19169 : BUF_X1 port map( A => n21543, Z => n25441);
   U19170 : BUF_X1 port map( A => n21550, Z => n25402);
   U19171 : BUF_X1 port map( A => n21536, Z => n25480);
   U19172 : BUF_X1 port map( A => n21541, Z => n25454);
   U19173 : BUF_X1 port map( A => n21554, Z => n25376);
   U19174 : BUF_X1 port map( A => n21526, Z => n25531);
   U19175 : BUF_X1 port map( A => n21492, Z => n25724);
   U19176 : BUF_X1 port map( A => n21506, Z => n25647);
   U19177 : BUF_X1 port map( A => n21547, Z => n25415);
   U19178 : BUF_X1 port map( A => n21552, Z => n25389);
   U19179 : BUF_X1 port map( A => n21510, Z => n25621);
   U19180 : BUF_X1 port map( A => n21524, Z => n25544);
   U19181 : BUF_X1 port map( A => n21529, Z => n25518);
   U19182 : BUF_X1 port map( A => n21545, Z => n25428);
   U19183 : BUF_X1 port map( A => n21534, Z => n25493);
   U19184 : BUF_X1 port map( A => n21513, Z => n25608);
   U19185 : BUF_X1 port map( A => n21504, Z => n25660);
   U19186 : BUF_X1 port map( A => n21501, Z => n25673);
   U19187 : BUF_X1 port map( A => n21497, Z => n25698);
   U19188 : BUF_X1 port map( A => n21495, Z => n25711);
   U19189 : BUF_X1 port map( A => n21482, Z => n25763);
   U19190 : BUF_X1 port map( A => n21488, Z => n25738);
   U19191 : BUF_X1 port map( A => n21515, Z => n25596);
   U19192 : BUF_X1 port map( A => n21522, Z => n25558);
   U19193 : BUF_X1 port map( A => n21538, Z => n25468);
   U19194 : BUF_X1 port map( A => n21508, Z => n25635);
   U19195 : BUF_X1 port map( A => n21543, Z => n25442);
   U19196 : BUF_X1 port map( A => n21550, Z => n25403);
   U19197 : BUF_X1 port map( A => n21536, Z => n25481);
   U19198 : BUF_X1 port map( A => n21541, Z => n25455);
   U19199 : BUF_X1 port map( A => n21554, Z => n25377);
   U19200 : BUF_X1 port map( A => n21526, Z => n25532);
   U19201 : BUF_X1 port map( A => n21492, Z => n25725);
   U19202 : BUF_X1 port map( A => n21506, Z => n25648);
   U19203 : BUF_X1 port map( A => n21510, Z => n25622);
   U19204 : BUF_X1 port map( A => n21524, Z => n25545);
   U19205 : BUF_X1 port map( A => n21529, Z => n25519);
   U19206 : BUF_X1 port map( A => n21547, Z => n25416);
   U19207 : BUF_X1 port map( A => n21552, Z => n25390);
   U19208 : BUF_X1 port map( A => n21545, Z => n25429);
   U19209 : BUF_X1 port map( A => n21534, Z => n25494);
   U19210 : BUF_X1 port map( A => n21513, Z => n25609);
   U19211 : BUF_X1 port map( A => n21504, Z => n25661);
   U19212 : BUF_X1 port map( A => n21501, Z => n25674);
   U19213 : BUF_X1 port map( A => n21497, Z => n25699);
   U19214 : BUF_X1 port map( A => n21495, Z => n25712);
   U19215 : OAI22_X1 port map( A1 => n25563, A2 => n21353, B1 => n25962, B2 => 
                           n25556, ZN => n6395);
   U19216 : OAI22_X1 port map( A1 => n25563, A2 => n21352, B1 => n25965, B2 => 
                           n25556, ZN => n6396);
   U19217 : OAI22_X1 port map( A1 => n25563, A2 => n21351, B1 => n25968, B2 => 
                           n25556, ZN => n6397);
   U19218 : OAI22_X1 port map( A1 => n25563, A2 => n21350, B1 => n25971, B2 => 
                           n25556, ZN => n6398);
   U19219 : OAI22_X1 port map( A1 => n25640, A2 => n21225, B1 => n25961, B2 => 
                           n25633, ZN => n6779);
   U19220 : OAI22_X1 port map( A1 => n25640, A2 => n21224, B1 => n25964, B2 => 
                           n25633, ZN => n6780);
   U19221 : OAI22_X1 port map( A1 => n25640, A2 => n21223, B1 => n25967, B2 => 
                           n25633, ZN => n6781);
   U19222 : OAI22_X1 port map( A1 => n25640, A2 => n21222, B1 => n25970, B2 => 
                           n25633, ZN => n6782);
   U19223 : OAI22_X1 port map( A1 => n25447, A2 => n21101, B1 => n25963, B2 => 
                           n25440, ZN => n5819);
   U19224 : OAI22_X1 port map( A1 => n25447, A2 => n21100, B1 => n25966, B2 => 
                           n25440, ZN => n5820);
   U19225 : OAI22_X1 port map( A1 => n25447, A2 => n21099, B1 => n25969, B2 => 
                           n25440, ZN => n5821);
   U19226 : OAI22_X1 port map( A1 => n25447, A2 => n21098, B1 => n25972, B2 => 
                           n25440, ZN => n5822);
   U19227 : OAI22_X1 port map( A1 => n25408, A2 => n21097, B1 => n25963, B2 => 
                           n25401, ZN => n5627);
   U19228 : OAI22_X1 port map( A1 => n25408, A2 => n21096, B1 => n25966, B2 => 
                           n25401, ZN => n5628);
   U19229 : OAI22_X1 port map( A1 => n25408, A2 => n21095, B1 => n25969, B2 => 
                           n25401, ZN => n5629);
   U19230 : OAI22_X1 port map( A1 => n25408, A2 => n21094, B1 => n25972, B2 => 
                           n25401, ZN => n5630);
   U19231 : OAI22_X1 port map( A1 => n25768, A2 => n20969, B1 => n25961, B2 => 
                           n25761, ZN => n7419);
   U19232 : OAI22_X1 port map( A1 => n25768, A2 => n20968, B1 => n25964, B2 => 
                           n25761, ZN => n7420);
   U19233 : OAI22_X1 port map( A1 => n25768, A2 => n20967, B1 => n25967, B2 => 
                           n25761, ZN => n7421);
   U19234 : OAI22_X1 port map( A1 => n25768, A2 => n20966, B1 => n25970, B2 => 
                           n25761, ZN => n7422);
   U19235 : OAI22_X1 port map( A1 => n25537, A2 => n20713, B1 => n25962, B2 => 
                           n25530, ZN => n6267);
   U19236 : OAI22_X1 port map( A1 => n25537, A2 => n20712, B1 => n25965, B2 => 
                           n25530, ZN => n6268);
   U19237 : OAI22_X1 port map( A1 => n25537, A2 => n20711, B1 => n25968, B2 => 
                           n25530, ZN => n6269);
   U19238 : OAI22_X1 port map( A1 => n25537, A2 => n20710, B1 => n25971, B2 => 
                           n25530, ZN => n6270);
   U19239 : OAI22_X1 port map( A1 => n25730, A2 => n20649, B1 => n25961, B2 => 
                           n25723, ZN => n7227);
   U19240 : OAI22_X1 port map( A1 => n25730, A2 => n20648, B1 => n25964, B2 => 
                           n25723, ZN => n7228);
   U19241 : OAI22_X1 port map( A1 => n25730, A2 => n20647, B1 => n25967, B2 => 
                           n25723, ZN => n7229);
   U19242 : OAI22_X1 port map( A1 => n25730, A2 => n20646, B1 => n25970, B2 => 
                           n25723, ZN => n7230);
   U19243 : OAI22_X1 port map( A1 => n25627, A2 => n20401, B1 => n25962, B2 => 
                           n25620, ZN => n6715);
   U19244 : OAI22_X1 port map( A1 => n25627, A2 => n20400, B1 => n25965, B2 => 
                           n25620, ZN => n6716);
   U19245 : OAI22_X1 port map( A1 => n25627, A2 => n20399, B1 => n25968, B2 => 
                           n25620, ZN => n6717);
   U19246 : OAI22_X1 port map( A1 => n25627, A2 => n20398, B1 => n25971, B2 => 
                           n25620, ZN => n6718);
   U19247 : OAI22_X1 port map( A1 => n25550, A2 => n20337, B1 => n25962, B2 => 
                           n25543, ZN => n6331);
   U19248 : OAI22_X1 port map( A1 => n25550, A2 => n20336, B1 => n25965, B2 => 
                           n25543, ZN => n6332);
   U19249 : OAI22_X1 port map( A1 => n25550, A2 => n20335, B1 => n25968, B2 => 
                           n25543, ZN => n6333);
   U19250 : OAI22_X1 port map( A1 => n25550, A2 => n20334, B1 => n25971, B2 => 
                           n25543, ZN => n6334);
   U19251 : OAI22_X1 port map( A1 => n25524, A2 => n20273, B1 => n25962, B2 => 
                           n25517, ZN => n6203);
   U19252 : OAI22_X1 port map( A1 => n25524, A2 => n20272, B1 => n25965, B2 => 
                           n25517, ZN => n6204);
   U19253 : OAI22_X1 port map( A1 => n25524, A2 => n20271, B1 => n25968, B2 => 
                           n25517, ZN => n6205);
   U19254 : OAI22_X1 port map( A1 => n25524, A2 => n20270, B1 => n25971, B2 => 
                           n25517, ZN => n6206);
   U19255 : OAI22_X1 port map( A1 => n25434, A2 => n20137, B1 => n25963, B2 => 
                           n25427, ZN => n5755);
   U19256 : OAI22_X1 port map( A1 => n25434, A2 => n20136, B1 => n25966, B2 => 
                           n25427, ZN => n5756);
   U19257 : OAI22_X1 port map( A1 => n25434, A2 => n20135, B1 => n25969, B2 => 
                           n25427, ZN => n5757);
   U19258 : OAI22_X1 port map( A1 => n25434, A2 => n20134, B1 => n25972, B2 => 
                           n25427, ZN => n5758);
   U19259 : OAI22_X1 port map( A1 => n25666, A2 => n20133, B1 => n25970, B2 => 
                           n25659, ZN => n6910);
   U19260 : OAI22_X1 port map( A1 => n25614, A2 => n19816, B1 => n25962, B2 => 
                           n25607, ZN => n6651);
   U19261 : OAI22_X1 port map( A1 => n25614, A2 => n19815, B1 => n25965, B2 => 
                           n25607, ZN => n6652);
   U19262 : OAI22_X1 port map( A1 => n25614, A2 => n19814, B1 => n25968, B2 => 
                           n25607, ZN => n6653);
   U19263 : OAI22_X1 port map( A1 => n25614, A2 => n19813, B1 => n25971, B2 => 
                           n25607, ZN => n6654);
   U19264 : OAI22_X1 port map( A1 => n25666, A2 => n19752, B1 => n25961, B2 => 
                           n25659, ZN => n6907);
   U19265 : OAI22_X1 port map( A1 => n25666, A2 => n19751, B1 => n25964, B2 => 
                           n25659, ZN => n6908);
   U19266 : OAI22_X1 port map( A1 => n25666, A2 => n19750, B1 => n25967, B2 => 
                           n25659, ZN => n6909);
   U19267 : OAI22_X1 port map( A1 => n25717, A2 => n19561, B1 => n25961, B2 => 
                           n25710, ZN => n7163);
   U19268 : OAI22_X1 port map( A1 => n25717, A2 => n19560, B1 => n25964, B2 => 
                           n25710, ZN => n7164);
   U19269 : OAI22_X1 port map( A1 => n25717, A2 => n19559, B1 => n25967, B2 => 
                           n25710, ZN => n7165);
   U19270 : OAI22_X1 port map( A1 => n25717, A2 => n19558, B1 => n25970, B2 => 
                           n25710, ZN => n7166);
   U19271 : OAI22_X1 port map( A1 => n25443, A2 => n21221, B1 => n25783, B2 => 
                           n25435, ZN => n5759);
   U19272 : OAI22_X1 port map( A1 => n25443, A2 => n21220, B1 => n25786, B2 => 
                           n25435, ZN => n5760);
   U19273 : OAI22_X1 port map( A1 => n25443, A2 => n21219, B1 => n25789, B2 => 
                           n25435, ZN => n5761);
   U19274 : OAI22_X1 port map( A1 => n25443, A2 => n21218, B1 => n25792, B2 => 
                           n25435, ZN => n5762);
   U19275 : OAI22_X1 port map( A1 => n25443, A2 => n21217, B1 => n25795, B2 => 
                           n25435, ZN => n5763);
   U19276 : OAI22_X1 port map( A1 => n25443, A2 => n21216, B1 => n25798, B2 => 
                           n25435, ZN => n5764);
   U19277 : OAI22_X1 port map( A1 => n25443, A2 => n21215, B1 => n25801, B2 => 
                           n25435, ZN => n5765);
   U19278 : OAI22_X1 port map( A1 => n25443, A2 => n21214, B1 => n25804, B2 => 
                           n25435, ZN => n5766);
   U19279 : OAI22_X1 port map( A1 => n25443, A2 => n21213, B1 => n25807, B2 => 
                           n25435, ZN => n5767);
   U19280 : OAI22_X1 port map( A1 => n25443, A2 => n21212, B1 => n25810, B2 => 
                           n25435, ZN => n5768);
   U19281 : OAI22_X1 port map( A1 => n25443, A2 => n21211, B1 => n25813, B2 => 
                           n25435, ZN => n5769);
   U19282 : OAI22_X1 port map( A1 => n25443, A2 => n21210, B1 => n25816, B2 => 
                           n25435, ZN => n5770);
   U19283 : OAI22_X1 port map( A1 => n25444, A2 => n21209, B1 => n25819, B2 => 
                           n25436, ZN => n5771);
   U19284 : OAI22_X1 port map( A1 => n25444, A2 => n21208, B1 => n25822, B2 => 
                           n25436, ZN => n5772);
   U19285 : OAI22_X1 port map( A1 => n25444, A2 => n21207, B1 => n25825, B2 => 
                           n25436, ZN => n5773);
   U19286 : OAI22_X1 port map( A1 => n25444, A2 => n21206, B1 => n25828, B2 => 
                           n25436, ZN => n5774);
   U19287 : OAI22_X1 port map( A1 => n25444, A2 => n21205, B1 => n25831, B2 => 
                           n25436, ZN => n5775);
   U19288 : OAI22_X1 port map( A1 => n25444, A2 => n21204, B1 => n25834, B2 => 
                           n25436, ZN => n5776);
   U19289 : OAI22_X1 port map( A1 => n25444, A2 => n21203, B1 => n25837, B2 => 
                           n25436, ZN => n5777);
   U19290 : OAI22_X1 port map( A1 => n25444, A2 => n21202, B1 => n25840, B2 => 
                           n25436, ZN => n5778);
   U19291 : OAI22_X1 port map( A1 => n25444, A2 => n21201, B1 => n25843, B2 => 
                           n25436, ZN => n5779);
   U19292 : OAI22_X1 port map( A1 => n25444, A2 => n21200, B1 => n25846, B2 => 
                           n25436, ZN => n5780);
   U19293 : OAI22_X1 port map( A1 => n25444, A2 => n21199, B1 => n25849, B2 => 
                           n25436, ZN => n5781);
   U19294 : OAI22_X1 port map( A1 => n25444, A2 => n21198, B1 => n25852, B2 => 
                           n25436, ZN => n5782);
   U19295 : OAI22_X1 port map( A1 => n25444, A2 => n21197, B1 => n25855, B2 => 
                           n25437, ZN => n5783);
   U19296 : OAI22_X1 port map( A1 => n25445, A2 => n21196, B1 => n25858, B2 => 
                           n25437, ZN => n5784);
   U19297 : OAI22_X1 port map( A1 => n25445, A2 => n21195, B1 => n25861, B2 => 
                           n25437, ZN => n5785);
   U19298 : OAI22_X1 port map( A1 => n25445, A2 => n21194, B1 => n25864, B2 => 
                           n25437, ZN => n5786);
   U19299 : OAI22_X1 port map( A1 => n25445, A2 => n21193, B1 => n25867, B2 => 
                           n25437, ZN => n5787);
   U19300 : OAI22_X1 port map( A1 => n25445, A2 => n21192, B1 => n25870, B2 => 
                           n25437, ZN => n5788);
   U19301 : OAI22_X1 port map( A1 => n25445, A2 => n21191, B1 => n25873, B2 => 
                           n25437, ZN => n5789);
   U19302 : OAI22_X1 port map( A1 => n25445, A2 => n21190, B1 => n25876, B2 => 
                           n25437, ZN => n5790);
   U19303 : OAI22_X1 port map( A1 => n25445, A2 => n21189, B1 => n25879, B2 => 
                           n25437, ZN => n5791);
   U19304 : OAI22_X1 port map( A1 => n25445, A2 => n21188, B1 => n25882, B2 => 
                           n25437, ZN => n5792);
   U19305 : OAI22_X1 port map( A1 => n25445, A2 => n21187, B1 => n25885, B2 => 
                           n25437, ZN => n5793);
   U19306 : OAI22_X1 port map( A1 => n25445, A2 => n21186, B1 => n25888, B2 => 
                           n25437, ZN => n5794);
   U19307 : OAI22_X1 port map( A1 => n25445, A2 => n21185, B1 => n25891, B2 => 
                           n25438, ZN => n5795);
   U19308 : OAI22_X1 port map( A1 => n25445, A2 => n21184, B1 => n25894, B2 => 
                           n25438, ZN => n5796);
   U19309 : OAI22_X1 port map( A1 => n25446, A2 => n21183, B1 => n25897, B2 => 
                           n25438, ZN => n5797);
   U19310 : OAI22_X1 port map( A1 => n25446, A2 => n21182, B1 => n25900, B2 => 
                           n25438, ZN => n5798);
   U19311 : OAI22_X1 port map( A1 => n25446, A2 => n21181, B1 => n25903, B2 => 
                           n25438, ZN => n5799);
   U19312 : OAI22_X1 port map( A1 => n25446, A2 => n21180, B1 => n25906, B2 => 
                           n25438, ZN => n5800);
   U19313 : OAI22_X1 port map( A1 => n25446, A2 => n21179, B1 => n25909, B2 => 
                           n25438, ZN => n5801);
   U19314 : OAI22_X1 port map( A1 => n25446, A2 => n21178, B1 => n25912, B2 => 
                           n25438, ZN => n5802);
   U19315 : OAI22_X1 port map( A1 => n25446, A2 => n21177, B1 => n25915, B2 => 
                           n25438, ZN => n5803);
   U19316 : OAI22_X1 port map( A1 => n25446, A2 => n21176, B1 => n25918, B2 => 
                           n25438, ZN => n5804);
   U19317 : OAI22_X1 port map( A1 => n25446, A2 => n21175, B1 => n25921, B2 => 
                           n25438, ZN => n5805);
   U19318 : OAI22_X1 port map( A1 => n25446, A2 => n21174, B1 => n25924, B2 => 
                           n25438, ZN => n5806);
   U19319 : OAI22_X1 port map( A1 => n25446, A2 => n21173, B1 => n25927, B2 => 
                           n25439, ZN => n5807);
   U19320 : OAI22_X1 port map( A1 => n25446, A2 => n21172, B1 => n25930, B2 => 
                           n25439, ZN => n5808);
   U19321 : OAI22_X1 port map( A1 => n25446, A2 => n21171, B1 => n25933, B2 => 
                           n25439, ZN => n5809);
   U19322 : OAI22_X1 port map( A1 => n25447, A2 => n21170, B1 => n25936, B2 => 
                           n25439, ZN => n5810);
   U19323 : OAI22_X1 port map( A1 => n25447, A2 => n21169, B1 => n25939, B2 => 
                           n25439, ZN => n5811);
   U19324 : OAI22_X1 port map( A1 => n25447, A2 => n21168, B1 => n25942, B2 => 
                           n25439, ZN => n5812);
   U19325 : OAI22_X1 port map( A1 => n25447, A2 => n21167, B1 => n25945, B2 => 
                           n25439, ZN => n5813);
   U19326 : OAI22_X1 port map( A1 => n25447, A2 => n21166, B1 => n25948, B2 => 
                           n25439, ZN => n5814);
   U19327 : OAI22_X1 port map( A1 => n25447, A2 => n21165, B1 => n25951, B2 => 
                           n25439, ZN => n5815);
   U19328 : OAI22_X1 port map( A1 => n25447, A2 => n21164, B1 => n25954, B2 => 
                           n25439, ZN => n5816);
   U19329 : OAI22_X1 port map( A1 => n25447, A2 => n21163, B1 => n25957, B2 => 
                           n25439, ZN => n5817);
   U19330 : OAI22_X1 port map( A1 => n25447, A2 => n21162, B1 => n25960, B2 => 
                           n25439, ZN => n5818);
   U19331 : OAI22_X1 port map( A1 => n25404, A2 => n21161, B1 => n25783, B2 => 
                           n25396, ZN => n5567);
   U19332 : OAI22_X1 port map( A1 => n25404, A2 => n21160, B1 => n25786, B2 => 
                           n25396, ZN => n5568);
   U19333 : OAI22_X1 port map( A1 => n25404, A2 => n21159, B1 => n25789, B2 => 
                           n25396, ZN => n5569);
   U19334 : OAI22_X1 port map( A1 => n25404, A2 => n21158, B1 => n25792, B2 => 
                           n25396, ZN => n5570);
   U19335 : OAI22_X1 port map( A1 => n25404, A2 => n21157, B1 => n25795, B2 => 
                           n25396, ZN => n5571);
   U19336 : OAI22_X1 port map( A1 => n25404, A2 => n21156, B1 => n25798, B2 => 
                           n25396, ZN => n5572);
   U19337 : OAI22_X1 port map( A1 => n25404, A2 => n21155, B1 => n25801, B2 => 
                           n25396, ZN => n5573);
   U19338 : OAI22_X1 port map( A1 => n25404, A2 => n21154, B1 => n25804, B2 => 
                           n25396, ZN => n5574);
   U19339 : OAI22_X1 port map( A1 => n25404, A2 => n21153, B1 => n25807, B2 => 
                           n25396, ZN => n5575);
   U19340 : OAI22_X1 port map( A1 => n25404, A2 => n21152, B1 => n25810, B2 => 
                           n25396, ZN => n5576);
   U19341 : OAI22_X1 port map( A1 => n25404, A2 => n21151, B1 => n25813, B2 => 
                           n25396, ZN => n5577);
   U19342 : OAI22_X1 port map( A1 => n25404, A2 => n21150, B1 => n25816, B2 => 
                           n25396, ZN => n5578);
   U19343 : OAI22_X1 port map( A1 => n25405, A2 => n21149, B1 => n25819, B2 => 
                           n25397, ZN => n5579);
   U19344 : OAI22_X1 port map( A1 => n25405, A2 => n21148, B1 => n25822, B2 => 
                           n25397, ZN => n5580);
   U19345 : OAI22_X1 port map( A1 => n25405, A2 => n21147, B1 => n25825, B2 => 
                           n25397, ZN => n5581);
   U19346 : OAI22_X1 port map( A1 => n25405, A2 => n21146, B1 => n25828, B2 => 
                           n25397, ZN => n5582);
   U19347 : OAI22_X1 port map( A1 => n25405, A2 => n21145, B1 => n25831, B2 => 
                           n25397, ZN => n5583);
   U19348 : OAI22_X1 port map( A1 => n25405, A2 => n21144, B1 => n25834, B2 => 
                           n25397, ZN => n5584);
   U19349 : OAI22_X1 port map( A1 => n25405, A2 => n21143, B1 => n25837, B2 => 
                           n25397, ZN => n5585);
   U19350 : OAI22_X1 port map( A1 => n25405, A2 => n21142, B1 => n25840, B2 => 
                           n25397, ZN => n5586);
   U19351 : OAI22_X1 port map( A1 => n25405, A2 => n21141, B1 => n25843, B2 => 
                           n25397, ZN => n5587);
   U19352 : OAI22_X1 port map( A1 => n25405, A2 => n21140, B1 => n25846, B2 => 
                           n25397, ZN => n5588);
   U19353 : OAI22_X1 port map( A1 => n25405, A2 => n21139, B1 => n25849, B2 => 
                           n25397, ZN => n5589);
   U19354 : OAI22_X1 port map( A1 => n25405, A2 => n21138, B1 => n25852, B2 => 
                           n25397, ZN => n5590);
   U19355 : OAI22_X1 port map( A1 => n25405, A2 => n21137, B1 => n25855, B2 => 
                           n25398, ZN => n5591);
   U19356 : OAI22_X1 port map( A1 => n25406, A2 => n21136, B1 => n25858, B2 => 
                           n25398, ZN => n5592);
   U19357 : OAI22_X1 port map( A1 => n25406, A2 => n21135, B1 => n25861, B2 => 
                           n25398, ZN => n5593);
   U19358 : OAI22_X1 port map( A1 => n25406, A2 => n21134, B1 => n25864, B2 => 
                           n25398, ZN => n5594);
   U19359 : OAI22_X1 port map( A1 => n25406, A2 => n21133, B1 => n25867, B2 => 
                           n25398, ZN => n5595);
   U19360 : OAI22_X1 port map( A1 => n25406, A2 => n21132, B1 => n25870, B2 => 
                           n25398, ZN => n5596);
   U19361 : OAI22_X1 port map( A1 => n25406, A2 => n21131, B1 => n25873, B2 => 
                           n25398, ZN => n5597);
   U19362 : OAI22_X1 port map( A1 => n25406, A2 => n21130, B1 => n25876, B2 => 
                           n25398, ZN => n5598);
   U19363 : OAI22_X1 port map( A1 => n25406, A2 => n21129, B1 => n25879, B2 => 
                           n25398, ZN => n5599);
   U19364 : OAI22_X1 port map( A1 => n25406, A2 => n21128, B1 => n25882, B2 => 
                           n25398, ZN => n5600);
   U19365 : OAI22_X1 port map( A1 => n25406, A2 => n21127, B1 => n25885, B2 => 
                           n25398, ZN => n5601);
   U19366 : OAI22_X1 port map( A1 => n25406, A2 => n21126, B1 => n25888, B2 => 
                           n25398, ZN => n5602);
   U19367 : OAI22_X1 port map( A1 => n25406, A2 => n21125, B1 => n25891, B2 => 
                           n25399, ZN => n5603);
   U19368 : OAI22_X1 port map( A1 => n25406, A2 => n21124, B1 => n25894, B2 => 
                           n25399, ZN => n5604);
   U19369 : OAI22_X1 port map( A1 => n25407, A2 => n21123, B1 => n25897, B2 => 
                           n25399, ZN => n5605);
   U19370 : OAI22_X1 port map( A1 => n25407, A2 => n21122, B1 => n25900, B2 => 
                           n25399, ZN => n5606);
   U19371 : OAI22_X1 port map( A1 => n25407, A2 => n21121, B1 => n25903, B2 => 
                           n25399, ZN => n5607);
   U19372 : OAI22_X1 port map( A1 => n25407, A2 => n21120, B1 => n25906, B2 => 
                           n25399, ZN => n5608);
   U19373 : OAI22_X1 port map( A1 => n25407, A2 => n21119, B1 => n25909, B2 => 
                           n25399, ZN => n5609);
   U19374 : OAI22_X1 port map( A1 => n25407, A2 => n21118, B1 => n25912, B2 => 
                           n25399, ZN => n5610);
   U19375 : OAI22_X1 port map( A1 => n25407, A2 => n21117, B1 => n25915, B2 => 
                           n25399, ZN => n5611);
   U19376 : OAI22_X1 port map( A1 => n25407, A2 => n21116, B1 => n25918, B2 => 
                           n25399, ZN => n5612);
   U19377 : OAI22_X1 port map( A1 => n25407, A2 => n21115, B1 => n25921, B2 => 
                           n25399, ZN => n5613);
   U19378 : OAI22_X1 port map( A1 => n25407, A2 => n21114, B1 => n25924, B2 => 
                           n25399, ZN => n5614);
   U19379 : OAI22_X1 port map( A1 => n25407, A2 => n21113, B1 => n25927, B2 => 
                           n25400, ZN => n5615);
   U19380 : OAI22_X1 port map( A1 => n25407, A2 => n21112, B1 => n25930, B2 => 
                           n25400, ZN => n5616);
   U19381 : OAI22_X1 port map( A1 => n25407, A2 => n21111, B1 => n25933, B2 => 
                           n25400, ZN => n5617);
   U19382 : OAI22_X1 port map( A1 => n25408, A2 => n21110, B1 => n25936, B2 => 
                           n25400, ZN => n5618);
   U19383 : OAI22_X1 port map( A1 => n25408, A2 => n21109, B1 => n25939, B2 => 
                           n25400, ZN => n5619);
   U19384 : OAI22_X1 port map( A1 => n25408, A2 => n21108, B1 => n25942, B2 => 
                           n25400, ZN => n5620);
   U19385 : OAI22_X1 port map( A1 => n25408, A2 => n21107, B1 => n25945, B2 => 
                           n25400, ZN => n5621);
   U19386 : OAI22_X1 port map( A1 => n25408, A2 => n21106, B1 => n25948, B2 => 
                           n25400, ZN => n5622);
   U19387 : OAI22_X1 port map( A1 => n25408, A2 => n21105, B1 => n25951, B2 => 
                           n25400, ZN => n5623);
   U19388 : OAI22_X1 port map( A1 => n25408, A2 => n21104, B1 => n25954, B2 => 
                           n25400, ZN => n5624);
   U19389 : OAI22_X1 port map( A1 => n25408, A2 => n21103, B1 => n25957, B2 => 
                           n25400, ZN => n5625);
   U19390 : OAI22_X1 port map( A1 => n25408, A2 => n21102, B1 => n25960, B2 => 
                           n25400, ZN => n5626);
   U19391 : OAI22_X1 port map( A1 => n25430, A2 => n20197, B1 => n25783, B2 => 
                           n25422, ZN => n5695);
   U19392 : OAI22_X1 port map( A1 => n25430, A2 => n20196, B1 => n25786, B2 => 
                           n25422, ZN => n5696);
   U19393 : OAI22_X1 port map( A1 => n25430, A2 => n20195, B1 => n25789, B2 => 
                           n25422, ZN => n5697);
   U19394 : OAI22_X1 port map( A1 => n25430, A2 => n20194, B1 => n25792, B2 => 
                           n25422, ZN => n5698);
   U19395 : OAI22_X1 port map( A1 => n25430, A2 => n20193, B1 => n25795, B2 => 
                           n25422, ZN => n5699);
   U19396 : OAI22_X1 port map( A1 => n25430, A2 => n20192, B1 => n25798, B2 => 
                           n25422, ZN => n5700);
   U19397 : OAI22_X1 port map( A1 => n25430, A2 => n20191, B1 => n25801, B2 => 
                           n25422, ZN => n5701);
   U19398 : OAI22_X1 port map( A1 => n25430, A2 => n20190, B1 => n25804, B2 => 
                           n25422, ZN => n5702);
   U19399 : OAI22_X1 port map( A1 => n25430, A2 => n20189, B1 => n25807, B2 => 
                           n25422, ZN => n5703);
   U19400 : OAI22_X1 port map( A1 => n25430, A2 => n20188, B1 => n25810, B2 => 
                           n25422, ZN => n5704);
   U19401 : OAI22_X1 port map( A1 => n25430, A2 => n20187, B1 => n25813, B2 => 
                           n25422, ZN => n5705);
   U19402 : OAI22_X1 port map( A1 => n25430, A2 => n20186, B1 => n25816, B2 => 
                           n25422, ZN => n5706);
   U19403 : OAI22_X1 port map( A1 => n25431, A2 => n20185, B1 => n25819, B2 => 
                           n25423, ZN => n5707);
   U19404 : OAI22_X1 port map( A1 => n25431, A2 => n20184, B1 => n25822, B2 => 
                           n25423, ZN => n5708);
   U19405 : OAI22_X1 port map( A1 => n25431, A2 => n20183, B1 => n25825, B2 => 
                           n25423, ZN => n5709);
   U19406 : OAI22_X1 port map( A1 => n25431, A2 => n20182, B1 => n25828, B2 => 
                           n25423, ZN => n5710);
   U19407 : OAI22_X1 port map( A1 => n25431, A2 => n20181, B1 => n25831, B2 => 
                           n25423, ZN => n5711);
   U19408 : OAI22_X1 port map( A1 => n25431, A2 => n20180, B1 => n25834, B2 => 
                           n25423, ZN => n5712);
   U19409 : OAI22_X1 port map( A1 => n25431, A2 => n20179, B1 => n25837, B2 => 
                           n25423, ZN => n5713);
   U19410 : OAI22_X1 port map( A1 => n25431, A2 => n20178, B1 => n25840, B2 => 
                           n25423, ZN => n5714);
   U19411 : OAI22_X1 port map( A1 => n25431, A2 => n20177, B1 => n25843, B2 => 
                           n25423, ZN => n5715);
   U19412 : OAI22_X1 port map( A1 => n25431, A2 => n20176, B1 => n25846, B2 => 
                           n25423, ZN => n5716);
   U19413 : OAI22_X1 port map( A1 => n25431, A2 => n20175, B1 => n25849, B2 => 
                           n25423, ZN => n5717);
   U19414 : OAI22_X1 port map( A1 => n25431, A2 => n20174, B1 => n25852, B2 => 
                           n25423, ZN => n5718);
   U19415 : OAI22_X1 port map( A1 => n25431, A2 => n20173, B1 => n25855, B2 => 
                           n25424, ZN => n5719);
   U19416 : OAI22_X1 port map( A1 => n25432, A2 => n20172, B1 => n25858, B2 => 
                           n25424, ZN => n5720);
   U19417 : OAI22_X1 port map( A1 => n25432, A2 => n20171, B1 => n25861, B2 => 
                           n25424, ZN => n5721);
   U19418 : OAI22_X1 port map( A1 => n25432, A2 => n20170, B1 => n25864, B2 => 
                           n25424, ZN => n5722);
   U19419 : OAI22_X1 port map( A1 => n25432, A2 => n20169, B1 => n25867, B2 => 
                           n25424, ZN => n5723);
   U19420 : OAI22_X1 port map( A1 => n25432, A2 => n20168, B1 => n25870, B2 => 
                           n25424, ZN => n5724);
   U19421 : OAI22_X1 port map( A1 => n25432, A2 => n20167, B1 => n25873, B2 => 
                           n25424, ZN => n5725);
   U19422 : OAI22_X1 port map( A1 => n25432, A2 => n20166, B1 => n25876, B2 => 
                           n25424, ZN => n5726);
   U19423 : OAI22_X1 port map( A1 => n25432, A2 => n20165, B1 => n25879, B2 => 
                           n25424, ZN => n5727);
   U19424 : OAI22_X1 port map( A1 => n25432, A2 => n20164, B1 => n25882, B2 => 
                           n25424, ZN => n5728);
   U19425 : OAI22_X1 port map( A1 => n25432, A2 => n20163, B1 => n25885, B2 => 
                           n25424, ZN => n5729);
   U19426 : OAI22_X1 port map( A1 => n25432, A2 => n20162, B1 => n25888, B2 => 
                           n25424, ZN => n5730);
   U19427 : OAI22_X1 port map( A1 => n25432, A2 => n20161, B1 => n25891, B2 => 
                           n25425, ZN => n5731);
   U19428 : OAI22_X1 port map( A1 => n25432, A2 => n20160, B1 => n25894, B2 => 
                           n25425, ZN => n5732);
   U19429 : OAI22_X1 port map( A1 => n25433, A2 => n20159, B1 => n25897, B2 => 
                           n25425, ZN => n5733);
   U19430 : OAI22_X1 port map( A1 => n25433, A2 => n20158, B1 => n25900, B2 => 
                           n25425, ZN => n5734);
   U19431 : OAI22_X1 port map( A1 => n25433, A2 => n20157, B1 => n25903, B2 => 
                           n25425, ZN => n5735);
   U19432 : OAI22_X1 port map( A1 => n25433, A2 => n20156, B1 => n25906, B2 => 
                           n25425, ZN => n5736);
   U19433 : OAI22_X1 port map( A1 => n25433, A2 => n20155, B1 => n25909, B2 => 
                           n25425, ZN => n5737);
   U19434 : OAI22_X1 port map( A1 => n25433, A2 => n20154, B1 => n25912, B2 => 
                           n25425, ZN => n5738);
   U19435 : OAI22_X1 port map( A1 => n25433, A2 => n20153, B1 => n25915, B2 => 
                           n25425, ZN => n5739);
   U19436 : OAI22_X1 port map( A1 => n25433, A2 => n20152, B1 => n25918, B2 => 
                           n25425, ZN => n5740);
   U19437 : OAI22_X1 port map( A1 => n25433, A2 => n20151, B1 => n25921, B2 => 
                           n25425, ZN => n5741);
   U19438 : OAI22_X1 port map( A1 => n25433, A2 => n20150, B1 => n25924, B2 => 
                           n25425, ZN => n5742);
   U19439 : OAI22_X1 port map( A1 => n25433, A2 => n20149, B1 => n25927, B2 => 
                           n25426, ZN => n5743);
   U19440 : OAI22_X1 port map( A1 => n25433, A2 => n20148, B1 => n25930, B2 => 
                           n25426, ZN => n5744);
   U19441 : OAI22_X1 port map( A1 => n25433, A2 => n20147, B1 => n25933, B2 => 
                           n25426, ZN => n5745);
   U19442 : OAI22_X1 port map( A1 => n25434, A2 => n20146, B1 => n25936, B2 => 
                           n25426, ZN => n5746);
   U19443 : OAI22_X1 port map( A1 => n25434, A2 => n20145, B1 => n25939, B2 => 
                           n25426, ZN => n5747);
   U19444 : OAI22_X1 port map( A1 => n25434, A2 => n20144, B1 => n25942, B2 => 
                           n25426, ZN => n5748);
   U19445 : OAI22_X1 port map( A1 => n25434, A2 => n20143, B1 => n25945, B2 => 
                           n25426, ZN => n5749);
   U19446 : OAI22_X1 port map( A1 => n25434, A2 => n20142, B1 => n25948, B2 => 
                           n25426, ZN => n5750);
   U19447 : OAI22_X1 port map( A1 => n25434, A2 => n20141, B1 => n25951, B2 => 
                           n25426, ZN => n5751);
   U19448 : OAI22_X1 port map( A1 => n25434, A2 => n20140, B1 => n25954, B2 => 
                           n25426, ZN => n5752);
   U19449 : OAI22_X1 port map( A1 => n25434, A2 => n20139, B1 => n25957, B2 => 
                           n25426, ZN => n5753);
   U19450 : OAI22_X1 port map( A1 => n25434, A2 => n20138, B1 => n25960, B2 => 
                           n25426, ZN => n5754);
   U19451 : OAI22_X1 port map( A1 => n25559, A2 => n21413, B1 => n25782, B2 => 
                           n25551, ZN => n6335);
   U19452 : OAI22_X1 port map( A1 => n25559, A2 => n21412, B1 => n25785, B2 => 
                           n25551, ZN => n6336);
   U19453 : OAI22_X1 port map( A1 => n25559, A2 => n21411, B1 => n25788, B2 => 
                           n25551, ZN => n6337);
   U19454 : OAI22_X1 port map( A1 => n25559, A2 => n21410, B1 => n25791, B2 => 
                           n25551, ZN => n6338);
   U19455 : OAI22_X1 port map( A1 => n25559, A2 => n21409, B1 => n25794, B2 => 
                           n25551, ZN => n6339);
   U19456 : OAI22_X1 port map( A1 => n25559, A2 => n21408, B1 => n25797, B2 => 
                           n25551, ZN => n6340);
   U19457 : OAI22_X1 port map( A1 => n25559, A2 => n21407, B1 => n25800, B2 => 
                           n25551, ZN => n6341);
   U19458 : OAI22_X1 port map( A1 => n25559, A2 => n21406, B1 => n25803, B2 => 
                           n25551, ZN => n6342);
   U19459 : OAI22_X1 port map( A1 => n25559, A2 => n21405, B1 => n25806, B2 => 
                           n25551, ZN => n6343);
   U19460 : OAI22_X1 port map( A1 => n25559, A2 => n21404, B1 => n25809, B2 => 
                           n25551, ZN => n6344);
   U19461 : OAI22_X1 port map( A1 => n25559, A2 => n21403, B1 => n25812, B2 => 
                           n25551, ZN => n6345);
   U19462 : OAI22_X1 port map( A1 => n25559, A2 => n21402, B1 => n25815, B2 => 
                           n25551, ZN => n6346);
   U19463 : OAI22_X1 port map( A1 => n25560, A2 => n21401, B1 => n25818, B2 => 
                           n25552, ZN => n6347);
   U19464 : OAI22_X1 port map( A1 => n25560, A2 => n21400, B1 => n25821, B2 => 
                           n25552, ZN => n6348);
   U19465 : OAI22_X1 port map( A1 => n25560, A2 => n21399, B1 => n25824, B2 => 
                           n25552, ZN => n6349);
   U19466 : OAI22_X1 port map( A1 => n25560, A2 => n21398, B1 => n25827, B2 => 
                           n25552, ZN => n6350);
   U19467 : OAI22_X1 port map( A1 => n25560, A2 => n21397, B1 => n25830, B2 => 
                           n25552, ZN => n6351);
   U19468 : OAI22_X1 port map( A1 => n25560, A2 => n21396, B1 => n25833, B2 => 
                           n25552, ZN => n6352);
   U19469 : OAI22_X1 port map( A1 => n25560, A2 => n21395, B1 => n25836, B2 => 
                           n25552, ZN => n6353);
   U19470 : OAI22_X1 port map( A1 => n25560, A2 => n21394, B1 => n25839, B2 => 
                           n25552, ZN => n6354);
   U19471 : OAI22_X1 port map( A1 => n25560, A2 => n21393, B1 => n25842, B2 => 
                           n25552, ZN => n6355);
   U19472 : OAI22_X1 port map( A1 => n25560, A2 => n21392, B1 => n25845, B2 => 
                           n25552, ZN => n6356);
   U19473 : OAI22_X1 port map( A1 => n25560, A2 => n21391, B1 => n25848, B2 => 
                           n25552, ZN => n6357);
   U19474 : OAI22_X1 port map( A1 => n25560, A2 => n21390, B1 => n25851, B2 => 
                           n25552, ZN => n6358);
   U19475 : OAI22_X1 port map( A1 => n25560, A2 => n21389, B1 => n25854, B2 => 
                           n25553, ZN => n6359);
   U19476 : OAI22_X1 port map( A1 => n25561, A2 => n21388, B1 => n25857, B2 => 
                           n25553, ZN => n6360);
   U19477 : OAI22_X1 port map( A1 => n25561, A2 => n21387, B1 => n25860, B2 => 
                           n25553, ZN => n6361);
   U19478 : OAI22_X1 port map( A1 => n25561, A2 => n21386, B1 => n25863, B2 => 
                           n25553, ZN => n6362);
   U19479 : OAI22_X1 port map( A1 => n25561, A2 => n21385, B1 => n25866, B2 => 
                           n25553, ZN => n6363);
   U19480 : OAI22_X1 port map( A1 => n25561, A2 => n21384, B1 => n25869, B2 => 
                           n25553, ZN => n6364);
   U19481 : OAI22_X1 port map( A1 => n25561, A2 => n21383, B1 => n25872, B2 => 
                           n25553, ZN => n6365);
   U19482 : OAI22_X1 port map( A1 => n25561, A2 => n21382, B1 => n25875, B2 => 
                           n25553, ZN => n6366);
   U19483 : OAI22_X1 port map( A1 => n25561, A2 => n21381, B1 => n25878, B2 => 
                           n25553, ZN => n6367);
   U19484 : OAI22_X1 port map( A1 => n25561, A2 => n21380, B1 => n25881, B2 => 
                           n25553, ZN => n6368);
   U19485 : OAI22_X1 port map( A1 => n25561, A2 => n21379, B1 => n25884, B2 => 
                           n25553, ZN => n6369);
   U19486 : OAI22_X1 port map( A1 => n25561, A2 => n21378, B1 => n25887, B2 => 
                           n25553, ZN => n6370);
   U19487 : OAI22_X1 port map( A1 => n25561, A2 => n21377, B1 => n25890, B2 => 
                           n25554, ZN => n6371);
   U19488 : OAI22_X1 port map( A1 => n25561, A2 => n21376, B1 => n25893, B2 => 
                           n25554, ZN => n6372);
   U19489 : OAI22_X1 port map( A1 => n25562, A2 => n21375, B1 => n25896, B2 => 
                           n25554, ZN => n6373);
   U19490 : OAI22_X1 port map( A1 => n25562, A2 => n21374, B1 => n25899, B2 => 
                           n25554, ZN => n6374);
   U19491 : OAI22_X1 port map( A1 => n25562, A2 => n21373, B1 => n25902, B2 => 
                           n25554, ZN => n6375);
   U19492 : OAI22_X1 port map( A1 => n25562, A2 => n21372, B1 => n25905, B2 => 
                           n25554, ZN => n6376);
   U19493 : OAI22_X1 port map( A1 => n25562, A2 => n21371, B1 => n25908, B2 => 
                           n25554, ZN => n6377);
   U19494 : OAI22_X1 port map( A1 => n25562, A2 => n21370, B1 => n25911, B2 => 
                           n25554, ZN => n6378);
   U19495 : OAI22_X1 port map( A1 => n25562, A2 => n21369, B1 => n25914, B2 => 
                           n25554, ZN => n6379);
   U19496 : OAI22_X1 port map( A1 => n25562, A2 => n21368, B1 => n25917, B2 => 
                           n25554, ZN => n6380);
   U19497 : OAI22_X1 port map( A1 => n25562, A2 => n21367, B1 => n25920, B2 => 
                           n25554, ZN => n6381);
   U19498 : OAI22_X1 port map( A1 => n25562, A2 => n21366, B1 => n25923, B2 => 
                           n25554, ZN => n6382);
   U19499 : OAI22_X1 port map( A1 => n25562, A2 => n21365, B1 => n25926, B2 => 
                           n25555, ZN => n6383);
   U19500 : OAI22_X1 port map( A1 => n25562, A2 => n21364, B1 => n25929, B2 => 
                           n25555, ZN => n6384);
   U19501 : OAI22_X1 port map( A1 => n25562, A2 => n21363, B1 => n25932, B2 => 
                           n25555, ZN => n6385);
   U19502 : OAI22_X1 port map( A1 => n25563, A2 => n21362, B1 => n25935, B2 => 
                           n25555, ZN => n6386);
   U19503 : OAI22_X1 port map( A1 => n25563, A2 => n21361, B1 => n25938, B2 => 
                           n25555, ZN => n6387);
   U19504 : OAI22_X1 port map( A1 => n25563, A2 => n21360, B1 => n25941, B2 => 
                           n25555, ZN => n6388);
   U19505 : OAI22_X1 port map( A1 => n25563, A2 => n21359, B1 => n25944, B2 => 
                           n25555, ZN => n6389);
   U19506 : OAI22_X1 port map( A1 => n25563, A2 => n21358, B1 => n25947, B2 => 
                           n25555, ZN => n6390);
   U19507 : OAI22_X1 port map( A1 => n25563, A2 => n21357, B1 => n25950, B2 => 
                           n25555, ZN => n6391);
   U19508 : OAI22_X1 port map( A1 => n25563, A2 => n21356, B1 => n25953, B2 => 
                           n25555, ZN => n6392);
   U19509 : OAI22_X1 port map( A1 => n25563, A2 => n21355, B1 => n25956, B2 => 
                           n25555, ZN => n6393);
   U19510 : OAI22_X1 port map( A1 => n25563, A2 => n21354, B1 => n25959, B2 => 
                           n25555, ZN => n6394);
   U19511 : OAI22_X1 port map( A1 => n25636, A2 => n21285, B1 => n25781, B2 => 
                           n25628, ZN => n6719);
   U19512 : OAI22_X1 port map( A1 => n25636, A2 => n21284, B1 => n25784, B2 => 
                           n25628, ZN => n6720);
   U19513 : OAI22_X1 port map( A1 => n25636, A2 => n21283, B1 => n25787, B2 => 
                           n25628, ZN => n6721);
   U19514 : OAI22_X1 port map( A1 => n25636, A2 => n21282, B1 => n25790, B2 => 
                           n25628, ZN => n6722);
   U19515 : OAI22_X1 port map( A1 => n25636, A2 => n21281, B1 => n25793, B2 => 
                           n25628, ZN => n6723);
   U19516 : OAI22_X1 port map( A1 => n25636, A2 => n21280, B1 => n25796, B2 => 
                           n25628, ZN => n6724);
   U19517 : OAI22_X1 port map( A1 => n25636, A2 => n21279, B1 => n25799, B2 => 
                           n25628, ZN => n6725);
   U19518 : OAI22_X1 port map( A1 => n25636, A2 => n21278, B1 => n25802, B2 => 
                           n25628, ZN => n6726);
   U19519 : OAI22_X1 port map( A1 => n25636, A2 => n21277, B1 => n25805, B2 => 
                           n25628, ZN => n6727);
   U19520 : OAI22_X1 port map( A1 => n25636, A2 => n21276, B1 => n25808, B2 => 
                           n25628, ZN => n6728);
   U19521 : OAI22_X1 port map( A1 => n25636, A2 => n21275, B1 => n25811, B2 => 
                           n25628, ZN => n6729);
   U19522 : OAI22_X1 port map( A1 => n25636, A2 => n21274, B1 => n25814, B2 => 
                           n25628, ZN => n6730);
   U19523 : OAI22_X1 port map( A1 => n25637, A2 => n21273, B1 => n25817, B2 => 
                           n25629, ZN => n6731);
   U19524 : OAI22_X1 port map( A1 => n25637, A2 => n21272, B1 => n25820, B2 => 
                           n25629, ZN => n6732);
   U19525 : OAI22_X1 port map( A1 => n25637, A2 => n21271, B1 => n25823, B2 => 
                           n25629, ZN => n6733);
   U19526 : OAI22_X1 port map( A1 => n25637, A2 => n21270, B1 => n25826, B2 => 
                           n25629, ZN => n6734);
   U19527 : OAI22_X1 port map( A1 => n25637, A2 => n21269, B1 => n25829, B2 => 
                           n25629, ZN => n6735);
   U19528 : OAI22_X1 port map( A1 => n25637, A2 => n21268, B1 => n25832, B2 => 
                           n25629, ZN => n6736);
   U19529 : OAI22_X1 port map( A1 => n25637, A2 => n21267, B1 => n25835, B2 => 
                           n25629, ZN => n6737);
   U19530 : OAI22_X1 port map( A1 => n25637, A2 => n21266, B1 => n25838, B2 => 
                           n25629, ZN => n6738);
   U19531 : OAI22_X1 port map( A1 => n25637, A2 => n21265, B1 => n25841, B2 => 
                           n25629, ZN => n6739);
   U19532 : OAI22_X1 port map( A1 => n25637, A2 => n21264, B1 => n25844, B2 => 
                           n25629, ZN => n6740);
   U19533 : OAI22_X1 port map( A1 => n25637, A2 => n21263, B1 => n25847, B2 => 
                           n25629, ZN => n6741);
   U19534 : OAI22_X1 port map( A1 => n25637, A2 => n21262, B1 => n25850, B2 => 
                           n25629, ZN => n6742);
   U19535 : OAI22_X1 port map( A1 => n25637, A2 => n21261, B1 => n25853, B2 => 
                           n25630, ZN => n6743);
   U19536 : OAI22_X1 port map( A1 => n25638, A2 => n21260, B1 => n25856, B2 => 
                           n25630, ZN => n6744);
   U19537 : OAI22_X1 port map( A1 => n25638, A2 => n21259, B1 => n25859, B2 => 
                           n25630, ZN => n6745);
   U19538 : OAI22_X1 port map( A1 => n25638, A2 => n21258, B1 => n25862, B2 => 
                           n25630, ZN => n6746);
   U19539 : OAI22_X1 port map( A1 => n25638, A2 => n21257, B1 => n25865, B2 => 
                           n25630, ZN => n6747);
   U19540 : OAI22_X1 port map( A1 => n25638, A2 => n21256, B1 => n25868, B2 => 
                           n25630, ZN => n6748);
   U19541 : OAI22_X1 port map( A1 => n25638, A2 => n21255, B1 => n25871, B2 => 
                           n25630, ZN => n6749);
   U19542 : OAI22_X1 port map( A1 => n25638, A2 => n21254, B1 => n25874, B2 => 
                           n25630, ZN => n6750);
   U19543 : OAI22_X1 port map( A1 => n25638, A2 => n21253, B1 => n25877, B2 => 
                           n25630, ZN => n6751);
   U19544 : OAI22_X1 port map( A1 => n25638, A2 => n21252, B1 => n25880, B2 => 
                           n25630, ZN => n6752);
   U19545 : OAI22_X1 port map( A1 => n25638, A2 => n21251, B1 => n25883, B2 => 
                           n25630, ZN => n6753);
   U19546 : OAI22_X1 port map( A1 => n25638, A2 => n21250, B1 => n25886, B2 => 
                           n25630, ZN => n6754);
   U19547 : OAI22_X1 port map( A1 => n25638, A2 => n21249, B1 => n25889, B2 => 
                           n25631, ZN => n6755);
   U19548 : OAI22_X1 port map( A1 => n25638, A2 => n21248, B1 => n25892, B2 => 
                           n25631, ZN => n6756);
   U19549 : OAI22_X1 port map( A1 => n25639, A2 => n21247, B1 => n25895, B2 => 
                           n25631, ZN => n6757);
   U19550 : OAI22_X1 port map( A1 => n25639, A2 => n21246, B1 => n25898, B2 => 
                           n25631, ZN => n6758);
   U19551 : OAI22_X1 port map( A1 => n25639, A2 => n21245, B1 => n25901, B2 => 
                           n25631, ZN => n6759);
   U19552 : OAI22_X1 port map( A1 => n25639, A2 => n21244, B1 => n25904, B2 => 
                           n25631, ZN => n6760);
   U19553 : OAI22_X1 port map( A1 => n25639, A2 => n21243, B1 => n25907, B2 => 
                           n25631, ZN => n6761);
   U19554 : OAI22_X1 port map( A1 => n25639, A2 => n21242, B1 => n25910, B2 => 
                           n25631, ZN => n6762);
   U19555 : OAI22_X1 port map( A1 => n25639, A2 => n21241, B1 => n25913, B2 => 
                           n25631, ZN => n6763);
   U19556 : OAI22_X1 port map( A1 => n25639, A2 => n21240, B1 => n25916, B2 => 
                           n25631, ZN => n6764);
   U19557 : OAI22_X1 port map( A1 => n25639, A2 => n21239, B1 => n25919, B2 => 
                           n25631, ZN => n6765);
   U19558 : OAI22_X1 port map( A1 => n25639, A2 => n21238, B1 => n25922, B2 => 
                           n25631, ZN => n6766);
   U19559 : OAI22_X1 port map( A1 => n25639, A2 => n21237, B1 => n25925, B2 => 
                           n25632, ZN => n6767);
   U19560 : OAI22_X1 port map( A1 => n25639, A2 => n21236, B1 => n25928, B2 => 
                           n25632, ZN => n6768);
   U19561 : OAI22_X1 port map( A1 => n25639, A2 => n21235, B1 => n25931, B2 => 
                           n25632, ZN => n6769);
   U19562 : OAI22_X1 port map( A1 => n25640, A2 => n21234, B1 => n25934, B2 => 
                           n25632, ZN => n6770);
   U19563 : OAI22_X1 port map( A1 => n25640, A2 => n21233, B1 => n25937, B2 => 
                           n25632, ZN => n6771);
   U19564 : OAI22_X1 port map( A1 => n25640, A2 => n21232, B1 => n25940, B2 => 
                           n25632, ZN => n6772);
   U19565 : OAI22_X1 port map( A1 => n25640, A2 => n21231, B1 => n25943, B2 => 
                           n25632, ZN => n6773);
   U19566 : OAI22_X1 port map( A1 => n25640, A2 => n21230, B1 => n25946, B2 => 
                           n25632, ZN => n6774);
   U19567 : OAI22_X1 port map( A1 => n25640, A2 => n21229, B1 => n25949, B2 => 
                           n25632, ZN => n6775);
   U19568 : OAI22_X1 port map( A1 => n25640, A2 => n21228, B1 => n25952, B2 => 
                           n25632, ZN => n6776);
   U19569 : OAI22_X1 port map( A1 => n25640, A2 => n21227, B1 => n25955, B2 => 
                           n25632, ZN => n6777);
   U19570 : OAI22_X1 port map( A1 => n25640, A2 => n21226, B1 => n25958, B2 => 
                           n25632, ZN => n6778);
   U19571 : OAI22_X1 port map( A1 => n25764, A2 => n21029, B1 => n25781, B2 => 
                           n25756, ZN => n7359);
   U19572 : OAI22_X1 port map( A1 => n25764, A2 => n21028, B1 => n25784, B2 => 
                           n25756, ZN => n7360);
   U19573 : OAI22_X1 port map( A1 => n25764, A2 => n21027, B1 => n25787, B2 => 
                           n25756, ZN => n7361);
   U19574 : OAI22_X1 port map( A1 => n25764, A2 => n21026, B1 => n25790, B2 => 
                           n25756, ZN => n7362);
   U19575 : OAI22_X1 port map( A1 => n25764, A2 => n21025, B1 => n25793, B2 => 
                           n25756, ZN => n7363);
   U19576 : OAI22_X1 port map( A1 => n25764, A2 => n21024, B1 => n25796, B2 => 
                           n25756, ZN => n7364);
   U19577 : OAI22_X1 port map( A1 => n25764, A2 => n21023, B1 => n25799, B2 => 
                           n25756, ZN => n7365);
   U19578 : OAI22_X1 port map( A1 => n25764, A2 => n21022, B1 => n25802, B2 => 
                           n25756, ZN => n7366);
   U19579 : OAI22_X1 port map( A1 => n25764, A2 => n21021, B1 => n25805, B2 => 
                           n25756, ZN => n7367);
   U19580 : OAI22_X1 port map( A1 => n25764, A2 => n21020, B1 => n25808, B2 => 
                           n25756, ZN => n7368);
   U19581 : OAI22_X1 port map( A1 => n25764, A2 => n21019, B1 => n25811, B2 => 
                           n25756, ZN => n7369);
   U19582 : OAI22_X1 port map( A1 => n25764, A2 => n21018, B1 => n25814, B2 => 
                           n25756, ZN => n7370);
   U19583 : OAI22_X1 port map( A1 => n25765, A2 => n21017, B1 => n25817, B2 => 
                           n25757, ZN => n7371);
   U19584 : OAI22_X1 port map( A1 => n25765, A2 => n21016, B1 => n25820, B2 => 
                           n25757, ZN => n7372);
   U19585 : OAI22_X1 port map( A1 => n25765, A2 => n21015, B1 => n25823, B2 => 
                           n25757, ZN => n7373);
   U19586 : OAI22_X1 port map( A1 => n25765, A2 => n21014, B1 => n25826, B2 => 
                           n25757, ZN => n7374);
   U19587 : OAI22_X1 port map( A1 => n25765, A2 => n21013, B1 => n25829, B2 => 
                           n25757, ZN => n7375);
   U19588 : OAI22_X1 port map( A1 => n25765, A2 => n21012, B1 => n25832, B2 => 
                           n25757, ZN => n7376);
   U19589 : OAI22_X1 port map( A1 => n25765, A2 => n21011, B1 => n25835, B2 => 
                           n25757, ZN => n7377);
   U19590 : OAI22_X1 port map( A1 => n25765, A2 => n21010, B1 => n25838, B2 => 
                           n25757, ZN => n7378);
   U19591 : OAI22_X1 port map( A1 => n25765, A2 => n21009, B1 => n25841, B2 => 
                           n25757, ZN => n7379);
   U19592 : OAI22_X1 port map( A1 => n25765, A2 => n21008, B1 => n25844, B2 => 
                           n25757, ZN => n7380);
   U19593 : OAI22_X1 port map( A1 => n25765, A2 => n21007, B1 => n25847, B2 => 
                           n25757, ZN => n7381);
   U19594 : OAI22_X1 port map( A1 => n25765, A2 => n21006, B1 => n25850, B2 => 
                           n25757, ZN => n7382);
   U19595 : OAI22_X1 port map( A1 => n25765, A2 => n21005, B1 => n25853, B2 => 
                           n25758, ZN => n7383);
   U19596 : OAI22_X1 port map( A1 => n25766, A2 => n21004, B1 => n25856, B2 => 
                           n25758, ZN => n7384);
   U19597 : OAI22_X1 port map( A1 => n25766, A2 => n21003, B1 => n25859, B2 => 
                           n25758, ZN => n7385);
   U19598 : OAI22_X1 port map( A1 => n25766, A2 => n21002, B1 => n25862, B2 => 
                           n25758, ZN => n7386);
   U19599 : OAI22_X1 port map( A1 => n25766, A2 => n21001, B1 => n25865, B2 => 
                           n25758, ZN => n7387);
   U19600 : OAI22_X1 port map( A1 => n25766, A2 => n21000, B1 => n25868, B2 => 
                           n25758, ZN => n7388);
   U19601 : OAI22_X1 port map( A1 => n25766, A2 => n20999, B1 => n25871, B2 => 
                           n25758, ZN => n7389);
   U19602 : OAI22_X1 port map( A1 => n25766, A2 => n20998, B1 => n25874, B2 => 
                           n25758, ZN => n7390);
   U19603 : OAI22_X1 port map( A1 => n25766, A2 => n20997, B1 => n25877, B2 => 
                           n25758, ZN => n7391);
   U19604 : OAI22_X1 port map( A1 => n25766, A2 => n20996, B1 => n25880, B2 => 
                           n25758, ZN => n7392);
   U19605 : OAI22_X1 port map( A1 => n25766, A2 => n20995, B1 => n25883, B2 => 
                           n25758, ZN => n7393);
   U19606 : OAI22_X1 port map( A1 => n25766, A2 => n20994, B1 => n25886, B2 => 
                           n25758, ZN => n7394);
   U19607 : OAI22_X1 port map( A1 => n25766, A2 => n20993, B1 => n25889, B2 => 
                           n25759, ZN => n7395);
   U19608 : OAI22_X1 port map( A1 => n25766, A2 => n20992, B1 => n25892, B2 => 
                           n25759, ZN => n7396);
   U19609 : OAI22_X1 port map( A1 => n25767, A2 => n20991, B1 => n25895, B2 => 
                           n25759, ZN => n7397);
   U19610 : OAI22_X1 port map( A1 => n25767, A2 => n20990, B1 => n25898, B2 => 
                           n25759, ZN => n7398);
   U19611 : OAI22_X1 port map( A1 => n25767, A2 => n20989, B1 => n25901, B2 => 
                           n25759, ZN => n7399);
   U19612 : OAI22_X1 port map( A1 => n25767, A2 => n20988, B1 => n25904, B2 => 
                           n25759, ZN => n7400);
   U19613 : OAI22_X1 port map( A1 => n25767, A2 => n20987, B1 => n25907, B2 => 
                           n25759, ZN => n7401);
   U19614 : OAI22_X1 port map( A1 => n25767, A2 => n20986, B1 => n25910, B2 => 
                           n25759, ZN => n7402);
   U19615 : OAI22_X1 port map( A1 => n25767, A2 => n20985, B1 => n25913, B2 => 
                           n25759, ZN => n7403);
   U19616 : OAI22_X1 port map( A1 => n25767, A2 => n20984, B1 => n25916, B2 => 
                           n25759, ZN => n7404);
   U19617 : OAI22_X1 port map( A1 => n25767, A2 => n20983, B1 => n25919, B2 => 
                           n25759, ZN => n7405);
   U19618 : OAI22_X1 port map( A1 => n25767, A2 => n20982, B1 => n25922, B2 => 
                           n25759, ZN => n7406);
   U19619 : OAI22_X1 port map( A1 => n25767, A2 => n20981, B1 => n25925, B2 => 
                           n25760, ZN => n7407);
   U19620 : OAI22_X1 port map( A1 => n25767, A2 => n20980, B1 => n25928, B2 => 
                           n25760, ZN => n7408);
   U19621 : OAI22_X1 port map( A1 => n25767, A2 => n20979, B1 => n25931, B2 => 
                           n25760, ZN => n7409);
   U19622 : OAI22_X1 port map( A1 => n25768, A2 => n20978, B1 => n25934, B2 => 
                           n25760, ZN => n7410);
   U19623 : OAI22_X1 port map( A1 => n25768, A2 => n20977, B1 => n25937, B2 => 
                           n25760, ZN => n7411);
   U19624 : OAI22_X1 port map( A1 => n25768, A2 => n20976, B1 => n25940, B2 => 
                           n25760, ZN => n7412);
   U19625 : OAI22_X1 port map( A1 => n25768, A2 => n20975, B1 => n25943, B2 => 
                           n25760, ZN => n7413);
   U19626 : OAI22_X1 port map( A1 => n25768, A2 => n20974, B1 => n25946, B2 => 
                           n25760, ZN => n7414);
   U19627 : OAI22_X1 port map( A1 => n25768, A2 => n20973, B1 => n25949, B2 => 
                           n25760, ZN => n7415);
   U19628 : OAI22_X1 port map( A1 => n25768, A2 => n20972, B1 => n25952, B2 => 
                           n25760, ZN => n7416);
   U19629 : OAI22_X1 port map( A1 => n25768, A2 => n20971, B1 => n25955, B2 => 
                           n25760, ZN => n7417);
   U19630 : OAI22_X1 port map( A1 => n25768, A2 => n20970, B1 => n25958, B2 => 
                           n25760, ZN => n7418);
   U19631 : OAI22_X1 port map( A1 => n25533, A2 => n20773, B1 => n25782, B2 => 
                           n25525, ZN => n6207);
   U19632 : OAI22_X1 port map( A1 => n25533, A2 => n20772, B1 => n25785, B2 => 
                           n25525, ZN => n6208);
   U19633 : OAI22_X1 port map( A1 => n25533, A2 => n20771, B1 => n25788, B2 => 
                           n25525, ZN => n6209);
   U19634 : OAI22_X1 port map( A1 => n25533, A2 => n20770, B1 => n25791, B2 => 
                           n25525, ZN => n6210);
   U19635 : OAI22_X1 port map( A1 => n25533, A2 => n20769, B1 => n25794, B2 => 
                           n25525, ZN => n6211);
   U19636 : OAI22_X1 port map( A1 => n25533, A2 => n20768, B1 => n25797, B2 => 
                           n25525, ZN => n6212);
   U19637 : OAI22_X1 port map( A1 => n25533, A2 => n20767, B1 => n25800, B2 => 
                           n25525, ZN => n6213);
   U19638 : OAI22_X1 port map( A1 => n25533, A2 => n20766, B1 => n25803, B2 => 
                           n25525, ZN => n6214);
   U19639 : OAI22_X1 port map( A1 => n25533, A2 => n20765, B1 => n25806, B2 => 
                           n25525, ZN => n6215);
   U19640 : OAI22_X1 port map( A1 => n25533, A2 => n20764, B1 => n25809, B2 => 
                           n25525, ZN => n6216);
   U19641 : OAI22_X1 port map( A1 => n25533, A2 => n20763, B1 => n25812, B2 => 
                           n25525, ZN => n6217);
   U19642 : OAI22_X1 port map( A1 => n25533, A2 => n20762, B1 => n25815, B2 => 
                           n25525, ZN => n6218);
   U19643 : OAI22_X1 port map( A1 => n25534, A2 => n20761, B1 => n25818, B2 => 
                           n25526, ZN => n6219);
   U19644 : OAI22_X1 port map( A1 => n25534, A2 => n20760, B1 => n25821, B2 => 
                           n25526, ZN => n6220);
   U19645 : OAI22_X1 port map( A1 => n25534, A2 => n20759, B1 => n25824, B2 => 
                           n25526, ZN => n6221);
   U19646 : OAI22_X1 port map( A1 => n25534, A2 => n20758, B1 => n25827, B2 => 
                           n25526, ZN => n6222);
   U19647 : OAI22_X1 port map( A1 => n25534, A2 => n20757, B1 => n25830, B2 => 
                           n25526, ZN => n6223);
   U19648 : OAI22_X1 port map( A1 => n25534, A2 => n20756, B1 => n25833, B2 => 
                           n25526, ZN => n6224);
   U19649 : OAI22_X1 port map( A1 => n25534, A2 => n20755, B1 => n25836, B2 => 
                           n25526, ZN => n6225);
   U19650 : OAI22_X1 port map( A1 => n25534, A2 => n20754, B1 => n25839, B2 => 
                           n25526, ZN => n6226);
   U19651 : OAI22_X1 port map( A1 => n25534, A2 => n20753, B1 => n25842, B2 => 
                           n25526, ZN => n6227);
   U19652 : OAI22_X1 port map( A1 => n25534, A2 => n20752, B1 => n25845, B2 => 
                           n25526, ZN => n6228);
   U19653 : OAI22_X1 port map( A1 => n25534, A2 => n20751, B1 => n25848, B2 => 
                           n25526, ZN => n6229);
   U19654 : OAI22_X1 port map( A1 => n25534, A2 => n20750, B1 => n25851, B2 => 
                           n25526, ZN => n6230);
   U19655 : OAI22_X1 port map( A1 => n25534, A2 => n20749, B1 => n25854, B2 => 
                           n25527, ZN => n6231);
   U19656 : OAI22_X1 port map( A1 => n25535, A2 => n20748, B1 => n25857, B2 => 
                           n25527, ZN => n6232);
   U19657 : OAI22_X1 port map( A1 => n25535, A2 => n20747, B1 => n25860, B2 => 
                           n25527, ZN => n6233);
   U19658 : OAI22_X1 port map( A1 => n25535, A2 => n20746, B1 => n25863, B2 => 
                           n25527, ZN => n6234);
   U19659 : OAI22_X1 port map( A1 => n25535, A2 => n20745, B1 => n25866, B2 => 
                           n25527, ZN => n6235);
   U19660 : OAI22_X1 port map( A1 => n25535, A2 => n20744, B1 => n25869, B2 => 
                           n25527, ZN => n6236);
   U19661 : OAI22_X1 port map( A1 => n25535, A2 => n20743, B1 => n25872, B2 => 
                           n25527, ZN => n6237);
   U19662 : OAI22_X1 port map( A1 => n25535, A2 => n20742, B1 => n25875, B2 => 
                           n25527, ZN => n6238);
   U19663 : OAI22_X1 port map( A1 => n25535, A2 => n20741, B1 => n25878, B2 => 
                           n25527, ZN => n6239);
   U19664 : OAI22_X1 port map( A1 => n25535, A2 => n20740, B1 => n25881, B2 => 
                           n25527, ZN => n6240);
   U19665 : OAI22_X1 port map( A1 => n25535, A2 => n20739, B1 => n25884, B2 => 
                           n25527, ZN => n6241);
   U19666 : OAI22_X1 port map( A1 => n25535, A2 => n20738, B1 => n25887, B2 => 
                           n25527, ZN => n6242);
   U19667 : OAI22_X1 port map( A1 => n25535, A2 => n20737, B1 => n25890, B2 => 
                           n25528, ZN => n6243);
   U19668 : OAI22_X1 port map( A1 => n25535, A2 => n20736, B1 => n25893, B2 => 
                           n25528, ZN => n6244);
   U19669 : OAI22_X1 port map( A1 => n25536, A2 => n20735, B1 => n25896, B2 => 
                           n25528, ZN => n6245);
   U19670 : OAI22_X1 port map( A1 => n25536, A2 => n20734, B1 => n25899, B2 => 
                           n25528, ZN => n6246);
   U19671 : OAI22_X1 port map( A1 => n25536, A2 => n20733, B1 => n25902, B2 => 
                           n25528, ZN => n6247);
   U19672 : OAI22_X1 port map( A1 => n25536, A2 => n20732, B1 => n25905, B2 => 
                           n25528, ZN => n6248);
   U19673 : OAI22_X1 port map( A1 => n25536, A2 => n20731, B1 => n25908, B2 => 
                           n25528, ZN => n6249);
   U19674 : OAI22_X1 port map( A1 => n25536, A2 => n20730, B1 => n25911, B2 => 
                           n25528, ZN => n6250);
   U19675 : OAI22_X1 port map( A1 => n25536, A2 => n20729, B1 => n25914, B2 => 
                           n25528, ZN => n6251);
   U19676 : OAI22_X1 port map( A1 => n25536, A2 => n20728, B1 => n25917, B2 => 
                           n25528, ZN => n6252);
   U19677 : OAI22_X1 port map( A1 => n25536, A2 => n20727, B1 => n25920, B2 => 
                           n25528, ZN => n6253);
   U19678 : OAI22_X1 port map( A1 => n25536, A2 => n20726, B1 => n25923, B2 => 
                           n25528, ZN => n6254);
   U19679 : OAI22_X1 port map( A1 => n25536, A2 => n20725, B1 => n25926, B2 => 
                           n25529, ZN => n6255);
   U19680 : OAI22_X1 port map( A1 => n25536, A2 => n20724, B1 => n25929, B2 => 
                           n25529, ZN => n6256);
   U19681 : OAI22_X1 port map( A1 => n25536, A2 => n20723, B1 => n25932, B2 => 
                           n25529, ZN => n6257);
   U19682 : OAI22_X1 port map( A1 => n25537, A2 => n20722, B1 => n25935, B2 => 
                           n25529, ZN => n6258);
   U19683 : OAI22_X1 port map( A1 => n25537, A2 => n20721, B1 => n25938, B2 => 
                           n25529, ZN => n6259);
   U19684 : OAI22_X1 port map( A1 => n25537, A2 => n20720, B1 => n25941, B2 => 
                           n25529, ZN => n6260);
   U19685 : OAI22_X1 port map( A1 => n25537, A2 => n20719, B1 => n25944, B2 => 
                           n25529, ZN => n6261);
   U19686 : OAI22_X1 port map( A1 => n25537, A2 => n20718, B1 => n25947, B2 => 
                           n25529, ZN => n6262);
   U19687 : OAI22_X1 port map( A1 => n25537, A2 => n20717, B1 => n25950, B2 => 
                           n25529, ZN => n6263);
   U19688 : OAI22_X1 port map( A1 => n25537, A2 => n20716, B1 => n25953, B2 => 
                           n25529, ZN => n6264);
   U19689 : OAI22_X1 port map( A1 => n25537, A2 => n20715, B1 => n25956, B2 => 
                           n25529, ZN => n6265);
   U19690 : OAI22_X1 port map( A1 => n25537, A2 => n20714, B1 => n25959, B2 => 
                           n25529, ZN => n6266);
   U19691 : OAI22_X1 port map( A1 => n25726, A2 => n20709, B1 => n25781, B2 => 
                           n25718, ZN => n7167);
   U19692 : OAI22_X1 port map( A1 => n25726, A2 => n20708, B1 => n25784, B2 => 
                           n25718, ZN => n7168);
   U19693 : OAI22_X1 port map( A1 => n25726, A2 => n20707, B1 => n25787, B2 => 
                           n25718, ZN => n7169);
   U19694 : OAI22_X1 port map( A1 => n25726, A2 => n20706, B1 => n25790, B2 => 
                           n25718, ZN => n7170);
   U19695 : OAI22_X1 port map( A1 => n25726, A2 => n20705, B1 => n25793, B2 => 
                           n25718, ZN => n7171);
   U19696 : OAI22_X1 port map( A1 => n25726, A2 => n20704, B1 => n25796, B2 => 
                           n25718, ZN => n7172);
   U19697 : OAI22_X1 port map( A1 => n25726, A2 => n20703, B1 => n25799, B2 => 
                           n25718, ZN => n7173);
   U19698 : OAI22_X1 port map( A1 => n25726, A2 => n20702, B1 => n25802, B2 => 
                           n25718, ZN => n7174);
   U19699 : OAI22_X1 port map( A1 => n25726, A2 => n20701, B1 => n25805, B2 => 
                           n25718, ZN => n7175);
   U19700 : OAI22_X1 port map( A1 => n25726, A2 => n20700, B1 => n25808, B2 => 
                           n25718, ZN => n7176);
   U19701 : OAI22_X1 port map( A1 => n25726, A2 => n20699, B1 => n25811, B2 => 
                           n25718, ZN => n7177);
   U19702 : OAI22_X1 port map( A1 => n25726, A2 => n20698, B1 => n25814, B2 => 
                           n25718, ZN => n7178);
   U19703 : OAI22_X1 port map( A1 => n25727, A2 => n20697, B1 => n25817, B2 => 
                           n25719, ZN => n7179);
   U19704 : OAI22_X1 port map( A1 => n25727, A2 => n20696, B1 => n25820, B2 => 
                           n25719, ZN => n7180);
   U19705 : OAI22_X1 port map( A1 => n25727, A2 => n20695, B1 => n25823, B2 => 
                           n25719, ZN => n7181);
   U19706 : OAI22_X1 port map( A1 => n25727, A2 => n20694, B1 => n25826, B2 => 
                           n25719, ZN => n7182);
   U19707 : OAI22_X1 port map( A1 => n25727, A2 => n20693, B1 => n25829, B2 => 
                           n25719, ZN => n7183);
   U19708 : OAI22_X1 port map( A1 => n25727, A2 => n20692, B1 => n25832, B2 => 
                           n25719, ZN => n7184);
   U19709 : OAI22_X1 port map( A1 => n25727, A2 => n20691, B1 => n25835, B2 => 
                           n25719, ZN => n7185);
   U19710 : OAI22_X1 port map( A1 => n25727, A2 => n20690, B1 => n25838, B2 => 
                           n25719, ZN => n7186);
   U19711 : OAI22_X1 port map( A1 => n25727, A2 => n20689, B1 => n25841, B2 => 
                           n25719, ZN => n7187);
   U19712 : OAI22_X1 port map( A1 => n25727, A2 => n20688, B1 => n25844, B2 => 
                           n25719, ZN => n7188);
   U19713 : OAI22_X1 port map( A1 => n25727, A2 => n20687, B1 => n25847, B2 => 
                           n25719, ZN => n7189);
   U19714 : OAI22_X1 port map( A1 => n25727, A2 => n20686, B1 => n25850, B2 => 
                           n25719, ZN => n7190);
   U19715 : OAI22_X1 port map( A1 => n25727, A2 => n20685, B1 => n25853, B2 => 
                           n25720, ZN => n7191);
   U19716 : OAI22_X1 port map( A1 => n25728, A2 => n20684, B1 => n25856, B2 => 
                           n25720, ZN => n7192);
   U19717 : OAI22_X1 port map( A1 => n25728, A2 => n20683, B1 => n25859, B2 => 
                           n25720, ZN => n7193);
   U19718 : OAI22_X1 port map( A1 => n25728, A2 => n20682, B1 => n25862, B2 => 
                           n25720, ZN => n7194);
   U19719 : OAI22_X1 port map( A1 => n25728, A2 => n20681, B1 => n25865, B2 => 
                           n25720, ZN => n7195);
   U19720 : OAI22_X1 port map( A1 => n25728, A2 => n20680, B1 => n25868, B2 => 
                           n25720, ZN => n7196);
   U19721 : OAI22_X1 port map( A1 => n25728, A2 => n20679, B1 => n25871, B2 => 
                           n25720, ZN => n7197);
   U19722 : OAI22_X1 port map( A1 => n25728, A2 => n20678, B1 => n25874, B2 => 
                           n25720, ZN => n7198);
   U19723 : OAI22_X1 port map( A1 => n25728, A2 => n20677, B1 => n25877, B2 => 
                           n25720, ZN => n7199);
   U19724 : OAI22_X1 port map( A1 => n25728, A2 => n20676, B1 => n25880, B2 => 
                           n25720, ZN => n7200);
   U19725 : OAI22_X1 port map( A1 => n25728, A2 => n20675, B1 => n25883, B2 => 
                           n25720, ZN => n7201);
   U19726 : OAI22_X1 port map( A1 => n25728, A2 => n20674, B1 => n25886, B2 => 
                           n25720, ZN => n7202);
   U19727 : OAI22_X1 port map( A1 => n25728, A2 => n20673, B1 => n25889, B2 => 
                           n25721, ZN => n7203);
   U19728 : OAI22_X1 port map( A1 => n25728, A2 => n20672, B1 => n25892, B2 => 
                           n25721, ZN => n7204);
   U19729 : OAI22_X1 port map( A1 => n25729, A2 => n20671, B1 => n25895, B2 => 
                           n25721, ZN => n7205);
   U19730 : OAI22_X1 port map( A1 => n25729, A2 => n20670, B1 => n25898, B2 => 
                           n25721, ZN => n7206);
   U19731 : OAI22_X1 port map( A1 => n25729, A2 => n20669, B1 => n25901, B2 => 
                           n25721, ZN => n7207);
   U19732 : OAI22_X1 port map( A1 => n25729, A2 => n20668, B1 => n25904, B2 => 
                           n25721, ZN => n7208);
   U19733 : OAI22_X1 port map( A1 => n25729, A2 => n20667, B1 => n25907, B2 => 
                           n25721, ZN => n7209);
   U19734 : OAI22_X1 port map( A1 => n25729, A2 => n20666, B1 => n25910, B2 => 
                           n25721, ZN => n7210);
   U19735 : OAI22_X1 port map( A1 => n25729, A2 => n20665, B1 => n25913, B2 => 
                           n25721, ZN => n7211);
   U19736 : OAI22_X1 port map( A1 => n25729, A2 => n20664, B1 => n25916, B2 => 
                           n25721, ZN => n7212);
   U19737 : OAI22_X1 port map( A1 => n25729, A2 => n20663, B1 => n25919, B2 => 
                           n25721, ZN => n7213);
   U19738 : OAI22_X1 port map( A1 => n25729, A2 => n20662, B1 => n25922, B2 => 
                           n25721, ZN => n7214);
   U19739 : OAI22_X1 port map( A1 => n25729, A2 => n20661, B1 => n25925, B2 => 
                           n25722, ZN => n7215);
   U19740 : OAI22_X1 port map( A1 => n25729, A2 => n20660, B1 => n25928, B2 => 
                           n25722, ZN => n7216);
   U19741 : OAI22_X1 port map( A1 => n25729, A2 => n20659, B1 => n25931, B2 => 
                           n25722, ZN => n7217);
   U19742 : OAI22_X1 port map( A1 => n25730, A2 => n20658, B1 => n25934, B2 => 
                           n25722, ZN => n7218);
   U19743 : OAI22_X1 port map( A1 => n25730, A2 => n20657, B1 => n25937, B2 => 
                           n25722, ZN => n7219);
   U19744 : OAI22_X1 port map( A1 => n25730, A2 => n20656, B1 => n25940, B2 => 
                           n25722, ZN => n7220);
   U19745 : OAI22_X1 port map( A1 => n25730, A2 => n20655, B1 => n25943, B2 => 
                           n25722, ZN => n7221);
   U19746 : OAI22_X1 port map( A1 => n25730, A2 => n20654, B1 => n25946, B2 => 
                           n25722, ZN => n7222);
   U19747 : OAI22_X1 port map( A1 => n25730, A2 => n20653, B1 => n25949, B2 => 
                           n25722, ZN => n7223);
   U19748 : OAI22_X1 port map( A1 => n25730, A2 => n20652, B1 => n25952, B2 => 
                           n25722, ZN => n7224);
   U19749 : OAI22_X1 port map( A1 => n25730, A2 => n20651, B1 => n25955, B2 => 
                           n25722, ZN => n7225);
   U19750 : OAI22_X1 port map( A1 => n25730, A2 => n20650, B1 => n25958, B2 => 
                           n25722, ZN => n7226);
   U19751 : OAI22_X1 port map( A1 => n25623, A2 => n20461, B1 => n25782, B2 => 
                           n25615, ZN => n6655);
   U19752 : OAI22_X1 port map( A1 => n25623, A2 => n20460, B1 => n25785, B2 => 
                           n25615, ZN => n6656);
   U19753 : OAI22_X1 port map( A1 => n25623, A2 => n20459, B1 => n25788, B2 => 
                           n25615, ZN => n6657);
   U19754 : OAI22_X1 port map( A1 => n25623, A2 => n20458, B1 => n25791, B2 => 
                           n25615, ZN => n6658);
   U19755 : OAI22_X1 port map( A1 => n25623, A2 => n20457, B1 => n25794, B2 => 
                           n25615, ZN => n6659);
   U19756 : OAI22_X1 port map( A1 => n25623, A2 => n20456, B1 => n25797, B2 => 
                           n25615, ZN => n6660);
   U19757 : OAI22_X1 port map( A1 => n25623, A2 => n20455, B1 => n25800, B2 => 
                           n25615, ZN => n6661);
   U19758 : OAI22_X1 port map( A1 => n25623, A2 => n20454, B1 => n25803, B2 => 
                           n25615, ZN => n6662);
   U19759 : OAI22_X1 port map( A1 => n25623, A2 => n20453, B1 => n25806, B2 => 
                           n25615, ZN => n6663);
   U19760 : OAI22_X1 port map( A1 => n25623, A2 => n20452, B1 => n25809, B2 => 
                           n25615, ZN => n6664);
   U19761 : OAI22_X1 port map( A1 => n25623, A2 => n20451, B1 => n25812, B2 => 
                           n25615, ZN => n6665);
   U19762 : OAI22_X1 port map( A1 => n25623, A2 => n20450, B1 => n25815, B2 => 
                           n25615, ZN => n6666);
   U19763 : OAI22_X1 port map( A1 => n25624, A2 => n20449, B1 => n25818, B2 => 
                           n25616, ZN => n6667);
   U19764 : OAI22_X1 port map( A1 => n25624, A2 => n20448, B1 => n25821, B2 => 
                           n25616, ZN => n6668);
   U19765 : OAI22_X1 port map( A1 => n25624, A2 => n20447, B1 => n25824, B2 => 
                           n25616, ZN => n6669);
   U19766 : OAI22_X1 port map( A1 => n25624, A2 => n20446, B1 => n25827, B2 => 
                           n25616, ZN => n6670);
   U19767 : OAI22_X1 port map( A1 => n25624, A2 => n20445, B1 => n25830, B2 => 
                           n25616, ZN => n6671);
   U19768 : OAI22_X1 port map( A1 => n25624, A2 => n20444, B1 => n25833, B2 => 
                           n25616, ZN => n6672);
   U19769 : OAI22_X1 port map( A1 => n25624, A2 => n20443, B1 => n25836, B2 => 
                           n25616, ZN => n6673);
   U19770 : OAI22_X1 port map( A1 => n25624, A2 => n20442, B1 => n25839, B2 => 
                           n25616, ZN => n6674);
   U19771 : OAI22_X1 port map( A1 => n25624, A2 => n20441, B1 => n25842, B2 => 
                           n25616, ZN => n6675);
   U19772 : OAI22_X1 port map( A1 => n25624, A2 => n20440, B1 => n25845, B2 => 
                           n25616, ZN => n6676);
   U19773 : OAI22_X1 port map( A1 => n25624, A2 => n20439, B1 => n25848, B2 => 
                           n25616, ZN => n6677);
   U19774 : OAI22_X1 port map( A1 => n25624, A2 => n20438, B1 => n25851, B2 => 
                           n25616, ZN => n6678);
   U19775 : OAI22_X1 port map( A1 => n25624, A2 => n20437, B1 => n25854, B2 => 
                           n25617, ZN => n6679);
   U19776 : OAI22_X1 port map( A1 => n25625, A2 => n20436, B1 => n25857, B2 => 
                           n25617, ZN => n6680);
   U19777 : OAI22_X1 port map( A1 => n25625, A2 => n20435, B1 => n25860, B2 => 
                           n25617, ZN => n6681);
   U19778 : OAI22_X1 port map( A1 => n25625, A2 => n20434, B1 => n25863, B2 => 
                           n25617, ZN => n6682);
   U19779 : OAI22_X1 port map( A1 => n25625, A2 => n20433, B1 => n25866, B2 => 
                           n25617, ZN => n6683);
   U19780 : OAI22_X1 port map( A1 => n25625, A2 => n20432, B1 => n25869, B2 => 
                           n25617, ZN => n6684);
   U19781 : OAI22_X1 port map( A1 => n25625, A2 => n20431, B1 => n25872, B2 => 
                           n25617, ZN => n6685);
   U19782 : OAI22_X1 port map( A1 => n25625, A2 => n20430, B1 => n25875, B2 => 
                           n25617, ZN => n6686);
   U19783 : OAI22_X1 port map( A1 => n25625, A2 => n20429, B1 => n25878, B2 => 
                           n25617, ZN => n6687);
   U19784 : OAI22_X1 port map( A1 => n25625, A2 => n20428, B1 => n25881, B2 => 
                           n25617, ZN => n6688);
   U19785 : OAI22_X1 port map( A1 => n25625, A2 => n20427, B1 => n25884, B2 => 
                           n25617, ZN => n6689);
   U19786 : OAI22_X1 port map( A1 => n25625, A2 => n20426, B1 => n25887, B2 => 
                           n25617, ZN => n6690);
   U19787 : OAI22_X1 port map( A1 => n25625, A2 => n20425, B1 => n25890, B2 => 
                           n25618, ZN => n6691);
   U19788 : OAI22_X1 port map( A1 => n25625, A2 => n20424, B1 => n25893, B2 => 
                           n25618, ZN => n6692);
   U19789 : OAI22_X1 port map( A1 => n25626, A2 => n20423, B1 => n25896, B2 => 
                           n25618, ZN => n6693);
   U19790 : OAI22_X1 port map( A1 => n25626, A2 => n20422, B1 => n25899, B2 => 
                           n25618, ZN => n6694);
   U19791 : OAI22_X1 port map( A1 => n25626, A2 => n20421, B1 => n25902, B2 => 
                           n25618, ZN => n6695);
   U19792 : OAI22_X1 port map( A1 => n25626, A2 => n20420, B1 => n25905, B2 => 
                           n25618, ZN => n6696);
   U19793 : OAI22_X1 port map( A1 => n25626, A2 => n20419, B1 => n25908, B2 => 
                           n25618, ZN => n6697);
   U19794 : OAI22_X1 port map( A1 => n25626, A2 => n20418, B1 => n25911, B2 => 
                           n25618, ZN => n6698);
   U19795 : OAI22_X1 port map( A1 => n25626, A2 => n20417, B1 => n25914, B2 => 
                           n25618, ZN => n6699);
   U19796 : OAI22_X1 port map( A1 => n25626, A2 => n20416, B1 => n25917, B2 => 
                           n25618, ZN => n6700);
   U19797 : OAI22_X1 port map( A1 => n25626, A2 => n20415, B1 => n25920, B2 => 
                           n25618, ZN => n6701);
   U19798 : OAI22_X1 port map( A1 => n25626, A2 => n20414, B1 => n25923, B2 => 
                           n25618, ZN => n6702);
   U19799 : OAI22_X1 port map( A1 => n25626, A2 => n20413, B1 => n25926, B2 => 
                           n25619, ZN => n6703);
   U19800 : OAI22_X1 port map( A1 => n25626, A2 => n20412, B1 => n25929, B2 => 
                           n25619, ZN => n6704);
   U19801 : OAI22_X1 port map( A1 => n25626, A2 => n20411, B1 => n25932, B2 => 
                           n25619, ZN => n6705);
   U19802 : OAI22_X1 port map( A1 => n25627, A2 => n20410, B1 => n25935, B2 => 
                           n25619, ZN => n6706);
   U19803 : OAI22_X1 port map( A1 => n25627, A2 => n20409, B1 => n25938, B2 => 
                           n25619, ZN => n6707);
   U19804 : OAI22_X1 port map( A1 => n25627, A2 => n20408, B1 => n25941, B2 => 
                           n25619, ZN => n6708);
   U19805 : OAI22_X1 port map( A1 => n25627, A2 => n20407, B1 => n25944, B2 => 
                           n25619, ZN => n6709);
   U19806 : OAI22_X1 port map( A1 => n25627, A2 => n20406, B1 => n25947, B2 => 
                           n25619, ZN => n6710);
   U19807 : OAI22_X1 port map( A1 => n25627, A2 => n20405, B1 => n25950, B2 => 
                           n25619, ZN => n6711);
   U19808 : OAI22_X1 port map( A1 => n25627, A2 => n20404, B1 => n25953, B2 => 
                           n25619, ZN => n6712);
   U19809 : OAI22_X1 port map( A1 => n25627, A2 => n20403, B1 => n25956, B2 => 
                           n25619, ZN => n6713);
   U19810 : OAI22_X1 port map( A1 => n25627, A2 => n20402, B1 => n25959, B2 => 
                           n25619, ZN => n6714);
   U19811 : OAI22_X1 port map( A1 => n25546, A2 => n20397, B1 => n25782, B2 => 
                           n25538, ZN => n6271);
   U19812 : OAI22_X1 port map( A1 => n25546, A2 => n20396, B1 => n25785, B2 => 
                           n25538, ZN => n6272);
   U19813 : OAI22_X1 port map( A1 => n25546, A2 => n20395, B1 => n25788, B2 => 
                           n25538, ZN => n6273);
   U19814 : OAI22_X1 port map( A1 => n25546, A2 => n20394, B1 => n25791, B2 => 
                           n25538, ZN => n6274);
   U19815 : OAI22_X1 port map( A1 => n25546, A2 => n20393, B1 => n25794, B2 => 
                           n25538, ZN => n6275);
   U19816 : OAI22_X1 port map( A1 => n25546, A2 => n20392, B1 => n25797, B2 => 
                           n25538, ZN => n6276);
   U19817 : OAI22_X1 port map( A1 => n25546, A2 => n20391, B1 => n25800, B2 => 
                           n25538, ZN => n6277);
   U19818 : OAI22_X1 port map( A1 => n25546, A2 => n20390, B1 => n25803, B2 => 
                           n25538, ZN => n6278);
   U19819 : OAI22_X1 port map( A1 => n25546, A2 => n20389, B1 => n25806, B2 => 
                           n25538, ZN => n6279);
   U19820 : OAI22_X1 port map( A1 => n25546, A2 => n20388, B1 => n25809, B2 => 
                           n25538, ZN => n6280);
   U19821 : OAI22_X1 port map( A1 => n25546, A2 => n20387, B1 => n25812, B2 => 
                           n25538, ZN => n6281);
   U19822 : OAI22_X1 port map( A1 => n25546, A2 => n20386, B1 => n25815, B2 => 
                           n25538, ZN => n6282);
   U19823 : OAI22_X1 port map( A1 => n25547, A2 => n20385, B1 => n25818, B2 => 
                           n25539, ZN => n6283);
   U19824 : OAI22_X1 port map( A1 => n25547, A2 => n20384, B1 => n25821, B2 => 
                           n25539, ZN => n6284);
   U19825 : OAI22_X1 port map( A1 => n25547, A2 => n20383, B1 => n25824, B2 => 
                           n25539, ZN => n6285);
   U19826 : OAI22_X1 port map( A1 => n25547, A2 => n20382, B1 => n25827, B2 => 
                           n25539, ZN => n6286);
   U19827 : OAI22_X1 port map( A1 => n25547, A2 => n20381, B1 => n25830, B2 => 
                           n25539, ZN => n6287);
   U19828 : OAI22_X1 port map( A1 => n25547, A2 => n20380, B1 => n25833, B2 => 
                           n25539, ZN => n6288);
   U19829 : OAI22_X1 port map( A1 => n25547, A2 => n20379, B1 => n25836, B2 => 
                           n25539, ZN => n6289);
   U19830 : OAI22_X1 port map( A1 => n25547, A2 => n20378, B1 => n25839, B2 => 
                           n25539, ZN => n6290);
   U19831 : OAI22_X1 port map( A1 => n25547, A2 => n20377, B1 => n25842, B2 => 
                           n25539, ZN => n6291);
   U19832 : OAI22_X1 port map( A1 => n25547, A2 => n20376, B1 => n25845, B2 => 
                           n25539, ZN => n6292);
   U19833 : OAI22_X1 port map( A1 => n25547, A2 => n20375, B1 => n25848, B2 => 
                           n25539, ZN => n6293);
   U19834 : OAI22_X1 port map( A1 => n25547, A2 => n20374, B1 => n25851, B2 => 
                           n25539, ZN => n6294);
   U19835 : OAI22_X1 port map( A1 => n25547, A2 => n20373, B1 => n25854, B2 => 
                           n25540, ZN => n6295);
   U19836 : OAI22_X1 port map( A1 => n25548, A2 => n20372, B1 => n25857, B2 => 
                           n25540, ZN => n6296);
   U19837 : OAI22_X1 port map( A1 => n25548, A2 => n20371, B1 => n25860, B2 => 
                           n25540, ZN => n6297);
   U19838 : OAI22_X1 port map( A1 => n25548, A2 => n20370, B1 => n25863, B2 => 
                           n25540, ZN => n6298);
   U19839 : OAI22_X1 port map( A1 => n25548, A2 => n20369, B1 => n25866, B2 => 
                           n25540, ZN => n6299);
   U19840 : OAI22_X1 port map( A1 => n25548, A2 => n20368, B1 => n25869, B2 => 
                           n25540, ZN => n6300);
   U19841 : OAI22_X1 port map( A1 => n25548, A2 => n20367, B1 => n25872, B2 => 
                           n25540, ZN => n6301);
   U19842 : OAI22_X1 port map( A1 => n25548, A2 => n20366, B1 => n25875, B2 => 
                           n25540, ZN => n6302);
   U19843 : OAI22_X1 port map( A1 => n25548, A2 => n20365, B1 => n25878, B2 => 
                           n25540, ZN => n6303);
   U19844 : OAI22_X1 port map( A1 => n25548, A2 => n20364, B1 => n25881, B2 => 
                           n25540, ZN => n6304);
   U19845 : OAI22_X1 port map( A1 => n25548, A2 => n20363, B1 => n25884, B2 => 
                           n25540, ZN => n6305);
   U19846 : OAI22_X1 port map( A1 => n25548, A2 => n20362, B1 => n25887, B2 => 
                           n25540, ZN => n6306);
   U19847 : OAI22_X1 port map( A1 => n25548, A2 => n20361, B1 => n25890, B2 => 
                           n25541, ZN => n6307);
   U19848 : OAI22_X1 port map( A1 => n25548, A2 => n20360, B1 => n25893, B2 => 
                           n25541, ZN => n6308);
   U19849 : OAI22_X1 port map( A1 => n25549, A2 => n20359, B1 => n25896, B2 => 
                           n25541, ZN => n6309);
   U19850 : OAI22_X1 port map( A1 => n25549, A2 => n20358, B1 => n25899, B2 => 
                           n25541, ZN => n6310);
   U19851 : OAI22_X1 port map( A1 => n25549, A2 => n20357, B1 => n25902, B2 => 
                           n25541, ZN => n6311);
   U19852 : OAI22_X1 port map( A1 => n25549, A2 => n20356, B1 => n25905, B2 => 
                           n25541, ZN => n6312);
   U19853 : OAI22_X1 port map( A1 => n25549, A2 => n20355, B1 => n25908, B2 => 
                           n25541, ZN => n6313);
   U19854 : OAI22_X1 port map( A1 => n25549, A2 => n20354, B1 => n25911, B2 => 
                           n25541, ZN => n6314);
   U19855 : OAI22_X1 port map( A1 => n25549, A2 => n20353, B1 => n25914, B2 => 
                           n25541, ZN => n6315);
   U19856 : OAI22_X1 port map( A1 => n25549, A2 => n20352, B1 => n25917, B2 => 
                           n25541, ZN => n6316);
   U19857 : OAI22_X1 port map( A1 => n25549, A2 => n20351, B1 => n25920, B2 => 
                           n25541, ZN => n6317);
   U19858 : OAI22_X1 port map( A1 => n25549, A2 => n20350, B1 => n25923, B2 => 
                           n25541, ZN => n6318);
   U19859 : OAI22_X1 port map( A1 => n25549, A2 => n20349, B1 => n25926, B2 => 
                           n25542, ZN => n6319);
   U19860 : OAI22_X1 port map( A1 => n25549, A2 => n20348, B1 => n25929, B2 => 
                           n25542, ZN => n6320);
   U19861 : OAI22_X1 port map( A1 => n25549, A2 => n20347, B1 => n25932, B2 => 
                           n25542, ZN => n6321);
   U19862 : OAI22_X1 port map( A1 => n25550, A2 => n20346, B1 => n25935, B2 => 
                           n25542, ZN => n6322);
   U19863 : OAI22_X1 port map( A1 => n25550, A2 => n20345, B1 => n25938, B2 => 
                           n25542, ZN => n6323);
   U19864 : OAI22_X1 port map( A1 => n25550, A2 => n20344, B1 => n25941, B2 => 
                           n25542, ZN => n6324);
   U19865 : OAI22_X1 port map( A1 => n25550, A2 => n20343, B1 => n25944, B2 => 
                           n25542, ZN => n6325);
   U19866 : OAI22_X1 port map( A1 => n25550, A2 => n20342, B1 => n25947, B2 => 
                           n25542, ZN => n6326);
   U19867 : OAI22_X1 port map( A1 => n25550, A2 => n20341, B1 => n25950, B2 => 
                           n25542, ZN => n6327);
   U19868 : OAI22_X1 port map( A1 => n25550, A2 => n20340, B1 => n25953, B2 => 
                           n25542, ZN => n6328);
   U19869 : OAI22_X1 port map( A1 => n25550, A2 => n20339, B1 => n25956, B2 => 
                           n25542, ZN => n6329);
   U19870 : OAI22_X1 port map( A1 => n25550, A2 => n20338, B1 => n25959, B2 => 
                           n25542, ZN => n6330);
   U19871 : OAI22_X1 port map( A1 => n25520, A2 => n20333, B1 => n25782, B2 => 
                           n25512, ZN => n6143);
   U19872 : OAI22_X1 port map( A1 => n25520, A2 => n20332, B1 => n25785, B2 => 
                           n25512, ZN => n6144);
   U19873 : OAI22_X1 port map( A1 => n25520, A2 => n20331, B1 => n25788, B2 => 
                           n25512, ZN => n6145);
   U19874 : OAI22_X1 port map( A1 => n25520, A2 => n20330, B1 => n25791, B2 => 
                           n25512, ZN => n6146);
   U19875 : OAI22_X1 port map( A1 => n25520, A2 => n20329, B1 => n25794, B2 => 
                           n25512, ZN => n6147);
   U19876 : OAI22_X1 port map( A1 => n25520, A2 => n20328, B1 => n25797, B2 => 
                           n25512, ZN => n6148);
   U19877 : OAI22_X1 port map( A1 => n25520, A2 => n20327, B1 => n25800, B2 => 
                           n25512, ZN => n6149);
   U19878 : OAI22_X1 port map( A1 => n25520, A2 => n20326, B1 => n25803, B2 => 
                           n25512, ZN => n6150);
   U19879 : OAI22_X1 port map( A1 => n25520, A2 => n20325, B1 => n25806, B2 => 
                           n25512, ZN => n6151);
   U19880 : OAI22_X1 port map( A1 => n25520, A2 => n20324, B1 => n25809, B2 => 
                           n25512, ZN => n6152);
   U19881 : OAI22_X1 port map( A1 => n25520, A2 => n20323, B1 => n25812, B2 => 
                           n25512, ZN => n6153);
   U19882 : OAI22_X1 port map( A1 => n25520, A2 => n20322, B1 => n25815, B2 => 
                           n25512, ZN => n6154);
   U19883 : OAI22_X1 port map( A1 => n25521, A2 => n20321, B1 => n25818, B2 => 
                           n25513, ZN => n6155);
   U19884 : OAI22_X1 port map( A1 => n25521, A2 => n20320, B1 => n25821, B2 => 
                           n25513, ZN => n6156);
   U19885 : OAI22_X1 port map( A1 => n25521, A2 => n20319, B1 => n25824, B2 => 
                           n25513, ZN => n6157);
   U19886 : OAI22_X1 port map( A1 => n25521, A2 => n20318, B1 => n25827, B2 => 
                           n25513, ZN => n6158);
   U19887 : OAI22_X1 port map( A1 => n25521, A2 => n20317, B1 => n25830, B2 => 
                           n25513, ZN => n6159);
   U19888 : OAI22_X1 port map( A1 => n25521, A2 => n20316, B1 => n25833, B2 => 
                           n25513, ZN => n6160);
   U19889 : OAI22_X1 port map( A1 => n25521, A2 => n20315, B1 => n25836, B2 => 
                           n25513, ZN => n6161);
   U19890 : OAI22_X1 port map( A1 => n25521, A2 => n20314, B1 => n25839, B2 => 
                           n25513, ZN => n6162);
   U19891 : OAI22_X1 port map( A1 => n25521, A2 => n20313, B1 => n25842, B2 => 
                           n25513, ZN => n6163);
   U19892 : OAI22_X1 port map( A1 => n25521, A2 => n20312, B1 => n25845, B2 => 
                           n25513, ZN => n6164);
   U19893 : OAI22_X1 port map( A1 => n25521, A2 => n20311, B1 => n25848, B2 => 
                           n25513, ZN => n6165);
   U19894 : OAI22_X1 port map( A1 => n25521, A2 => n20310, B1 => n25851, B2 => 
                           n25513, ZN => n6166);
   U19895 : OAI22_X1 port map( A1 => n25521, A2 => n20309, B1 => n25854, B2 => 
                           n25514, ZN => n6167);
   U19896 : OAI22_X1 port map( A1 => n25522, A2 => n20308, B1 => n25857, B2 => 
                           n25514, ZN => n6168);
   U19897 : OAI22_X1 port map( A1 => n25522, A2 => n20307, B1 => n25860, B2 => 
                           n25514, ZN => n6169);
   U19898 : OAI22_X1 port map( A1 => n25522, A2 => n20306, B1 => n25863, B2 => 
                           n25514, ZN => n6170);
   U19899 : OAI22_X1 port map( A1 => n25522, A2 => n20305, B1 => n25866, B2 => 
                           n25514, ZN => n6171);
   U19900 : OAI22_X1 port map( A1 => n25522, A2 => n20304, B1 => n25869, B2 => 
                           n25514, ZN => n6172);
   U19901 : OAI22_X1 port map( A1 => n25522, A2 => n20303, B1 => n25872, B2 => 
                           n25514, ZN => n6173);
   U19902 : OAI22_X1 port map( A1 => n25522, A2 => n20302, B1 => n25875, B2 => 
                           n25514, ZN => n6174);
   U19903 : OAI22_X1 port map( A1 => n25522, A2 => n20301, B1 => n25878, B2 => 
                           n25514, ZN => n6175);
   U19904 : OAI22_X1 port map( A1 => n25522, A2 => n20300, B1 => n25881, B2 => 
                           n25514, ZN => n6176);
   U19905 : OAI22_X1 port map( A1 => n25522, A2 => n20299, B1 => n25884, B2 => 
                           n25514, ZN => n6177);
   U19906 : OAI22_X1 port map( A1 => n25522, A2 => n20298, B1 => n25887, B2 => 
                           n25514, ZN => n6178);
   U19907 : OAI22_X1 port map( A1 => n25522, A2 => n20297, B1 => n25890, B2 => 
                           n25515, ZN => n6179);
   U19908 : OAI22_X1 port map( A1 => n25522, A2 => n20296, B1 => n25893, B2 => 
                           n25515, ZN => n6180);
   U19909 : OAI22_X1 port map( A1 => n25523, A2 => n20295, B1 => n25896, B2 => 
                           n25515, ZN => n6181);
   U19910 : OAI22_X1 port map( A1 => n25523, A2 => n20294, B1 => n25899, B2 => 
                           n25515, ZN => n6182);
   U19911 : OAI22_X1 port map( A1 => n25523, A2 => n20293, B1 => n25902, B2 => 
                           n25515, ZN => n6183);
   U19912 : OAI22_X1 port map( A1 => n25523, A2 => n20292, B1 => n25905, B2 => 
                           n25515, ZN => n6184);
   U19913 : OAI22_X1 port map( A1 => n25523, A2 => n20291, B1 => n25908, B2 => 
                           n25515, ZN => n6185);
   U19914 : OAI22_X1 port map( A1 => n25523, A2 => n20290, B1 => n25911, B2 => 
                           n25515, ZN => n6186);
   U19915 : OAI22_X1 port map( A1 => n25523, A2 => n20289, B1 => n25914, B2 => 
                           n25515, ZN => n6187);
   U19916 : OAI22_X1 port map( A1 => n25523, A2 => n20288, B1 => n25917, B2 => 
                           n25515, ZN => n6188);
   U19917 : OAI22_X1 port map( A1 => n25523, A2 => n20287, B1 => n25920, B2 => 
                           n25515, ZN => n6189);
   U19918 : OAI22_X1 port map( A1 => n25523, A2 => n20286, B1 => n25923, B2 => 
                           n25515, ZN => n6190);
   U19919 : OAI22_X1 port map( A1 => n25523, A2 => n20285, B1 => n25926, B2 => 
                           n25516, ZN => n6191);
   U19920 : OAI22_X1 port map( A1 => n25523, A2 => n20284, B1 => n25929, B2 => 
                           n25516, ZN => n6192);
   U19921 : OAI22_X1 port map( A1 => n25523, A2 => n20283, B1 => n25932, B2 => 
                           n25516, ZN => n6193);
   U19922 : OAI22_X1 port map( A1 => n25524, A2 => n20282, B1 => n25935, B2 => 
                           n25516, ZN => n6194);
   U19923 : OAI22_X1 port map( A1 => n25524, A2 => n20281, B1 => n25938, B2 => 
                           n25516, ZN => n6195);
   U19924 : OAI22_X1 port map( A1 => n25524, A2 => n20280, B1 => n25941, B2 => 
                           n25516, ZN => n6196);
   U19925 : OAI22_X1 port map( A1 => n25524, A2 => n20279, B1 => n25944, B2 => 
                           n25516, ZN => n6197);
   U19926 : OAI22_X1 port map( A1 => n25524, A2 => n20278, B1 => n25947, B2 => 
                           n25516, ZN => n6198);
   U19927 : OAI22_X1 port map( A1 => n25524, A2 => n20277, B1 => n25950, B2 => 
                           n25516, ZN => n6199);
   U19928 : OAI22_X1 port map( A1 => n25524, A2 => n20276, B1 => n25953, B2 => 
                           n25516, ZN => n6200);
   U19929 : OAI22_X1 port map( A1 => n25524, A2 => n20275, B1 => n25956, B2 => 
                           n25516, ZN => n6201);
   U19930 : OAI22_X1 port map( A1 => n25524, A2 => n20274, B1 => n25959, B2 => 
                           n25516, ZN => n6202);
   U19931 : OAI22_X1 port map( A1 => n25610, A2 => n19876, B1 => n25782, B2 => 
                           n25602, ZN => n6591);
   U19932 : OAI22_X1 port map( A1 => n25610, A2 => n19875, B1 => n25785, B2 => 
                           n25602, ZN => n6592);
   U19933 : OAI22_X1 port map( A1 => n25610, A2 => n19874, B1 => n25788, B2 => 
                           n25602, ZN => n6593);
   U19934 : OAI22_X1 port map( A1 => n25610, A2 => n19873, B1 => n25791, B2 => 
                           n25602, ZN => n6594);
   U19935 : OAI22_X1 port map( A1 => n25610, A2 => n19872, B1 => n25794, B2 => 
                           n25602, ZN => n6595);
   U19936 : OAI22_X1 port map( A1 => n25610, A2 => n19871, B1 => n25797, B2 => 
                           n25602, ZN => n6596);
   U19937 : OAI22_X1 port map( A1 => n25610, A2 => n19870, B1 => n25800, B2 => 
                           n25602, ZN => n6597);
   U19938 : OAI22_X1 port map( A1 => n25610, A2 => n19869, B1 => n25803, B2 => 
                           n25602, ZN => n6598);
   U19939 : OAI22_X1 port map( A1 => n25610, A2 => n19868, B1 => n25806, B2 => 
                           n25602, ZN => n6599);
   U19940 : OAI22_X1 port map( A1 => n25610, A2 => n19867, B1 => n25809, B2 => 
                           n25602, ZN => n6600);
   U19941 : OAI22_X1 port map( A1 => n25610, A2 => n19866, B1 => n25812, B2 => 
                           n25602, ZN => n6601);
   U19942 : OAI22_X1 port map( A1 => n25610, A2 => n19865, B1 => n25815, B2 => 
                           n25602, ZN => n6602);
   U19943 : OAI22_X1 port map( A1 => n25611, A2 => n19864, B1 => n25818, B2 => 
                           n25603, ZN => n6603);
   U19944 : OAI22_X1 port map( A1 => n25611, A2 => n19863, B1 => n25821, B2 => 
                           n25603, ZN => n6604);
   U19945 : OAI22_X1 port map( A1 => n25611, A2 => n19862, B1 => n25824, B2 => 
                           n25603, ZN => n6605);
   U19946 : OAI22_X1 port map( A1 => n25611, A2 => n19861, B1 => n25827, B2 => 
                           n25603, ZN => n6606);
   U19947 : OAI22_X1 port map( A1 => n25611, A2 => n19860, B1 => n25830, B2 => 
                           n25603, ZN => n6607);
   U19948 : OAI22_X1 port map( A1 => n25611, A2 => n19859, B1 => n25833, B2 => 
                           n25603, ZN => n6608);
   U19949 : OAI22_X1 port map( A1 => n25611, A2 => n19858, B1 => n25836, B2 => 
                           n25603, ZN => n6609);
   U19950 : OAI22_X1 port map( A1 => n25611, A2 => n19857, B1 => n25839, B2 => 
                           n25603, ZN => n6610);
   U19951 : OAI22_X1 port map( A1 => n25611, A2 => n19856, B1 => n25842, B2 => 
                           n25603, ZN => n6611);
   U19952 : OAI22_X1 port map( A1 => n25611, A2 => n19855, B1 => n25845, B2 => 
                           n25603, ZN => n6612);
   U19953 : OAI22_X1 port map( A1 => n25611, A2 => n19854, B1 => n25848, B2 => 
                           n25603, ZN => n6613);
   U19954 : OAI22_X1 port map( A1 => n25611, A2 => n19853, B1 => n25851, B2 => 
                           n25603, ZN => n6614);
   U19955 : OAI22_X1 port map( A1 => n25611, A2 => n19852, B1 => n25854, B2 => 
                           n25604, ZN => n6615);
   U19956 : OAI22_X1 port map( A1 => n25612, A2 => n19851, B1 => n25857, B2 => 
                           n25604, ZN => n6616);
   U19957 : OAI22_X1 port map( A1 => n25612, A2 => n19850, B1 => n25860, B2 => 
                           n25604, ZN => n6617);
   U19958 : OAI22_X1 port map( A1 => n25612, A2 => n19849, B1 => n25863, B2 => 
                           n25604, ZN => n6618);
   U19959 : OAI22_X1 port map( A1 => n25612, A2 => n19848, B1 => n25866, B2 => 
                           n25604, ZN => n6619);
   U19960 : OAI22_X1 port map( A1 => n25612, A2 => n19847, B1 => n25869, B2 => 
                           n25604, ZN => n6620);
   U19961 : OAI22_X1 port map( A1 => n25612, A2 => n19846, B1 => n25872, B2 => 
                           n25604, ZN => n6621);
   U19962 : OAI22_X1 port map( A1 => n25612, A2 => n19845, B1 => n25875, B2 => 
                           n25604, ZN => n6622);
   U19963 : OAI22_X1 port map( A1 => n25612, A2 => n19844, B1 => n25878, B2 => 
                           n25604, ZN => n6623);
   U19964 : OAI22_X1 port map( A1 => n25612, A2 => n19843, B1 => n25881, B2 => 
                           n25604, ZN => n6624);
   U19965 : OAI22_X1 port map( A1 => n25612, A2 => n19842, B1 => n25884, B2 => 
                           n25604, ZN => n6625);
   U19966 : OAI22_X1 port map( A1 => n25612, A2 => n19841, B1 => n25887, B2 => 
                           n25604, ZN => n6626);
   U19967 : OAI22_X1 port map( A1 => n25612, A2 => n19840, B1 => n25890, B2 => 
                           n25605, ZN => n6627);
   U19968 : OAI22_X1 port map( A1 => n25612, A2 => n19839, B1 => n25893, B2 => 
                           n25605, ZN => n6628);
   U19969 : OAI22_X1 port map( A1 => n25613, A2 => n19838, B1 => n25896, B2 => 
                           n25605, ZN => n6629);
   U19970 : OAI22_X1 port map( A1 => n25613, A2 => n19837, B1 => n25899, B2 => 
                           n25605, ZN => n6630);
   U19971 : OAI22_X1 port map( A1 => n25613, A2 => n19836, B1 => n25902, B2 => 
                           n25605, ZN => n6631);
   U19972 : OAI22_X1 port map( A1 => n25613, A2 => n19835, B1 => n25905, B2 => 
                           n25605, ZN => n6632);
   U19973 : OAI22_X1 port map( A1 => n25613, A2 => n19834, B1 => n25908, B2 => 
                           n25605, ZN => n6633);
   U19974 : OAI22_X1 port map( A1 => n25613, A2 => n19833, B1 => n25911, B2 => 
                           n25605, ZN => n6634);
   U19975 : OAI22_X1 port map( A1 => n25613, A2 => n19832, B1 => n25914, B2 => 
                           n25605, ZN => n6635);
   U19976 : OAI22_X1 port map( A1 => n25613, A2 => n19831, B1 => n25917, B2 => 
                           n25605, ZN => n6636);
   U19977 : OAI22_X1 port map( A1 => n25613, A2 => n19830, B1 => n25920, B2 => 
                           n25605, ZN => n6637);
   U19978 : OAI22_X1 port map( A1 => n25613, A2 => n19829, B1 => n25923, B2 => 
                           n25605, ZN => n6638);
   U19979 : OAI22_X1 port map( A1 => n25613, A2 => n19828, B1 => n25926, B2 => 
                           n25606, ZN => n6639);
   U19980 : OAI22_X1 port map( A1 => n25613, A2 => n19827, B1 => n25929, B2 => 
                           n25606, ZN => n6640);
   U19981 : OAI22_X1 port map( A1 => n25613, A2 => n19826, B1 => n25932, B2 => 
                           n25606, ZN => n6641);
   U19982 : OAI22_X1 port map( A1 => n25614, A2 => n19825, B1 => n25935, B2 => 
                           n25606, ZN => n6642);
   U19983 : OAI22_X1 port map( A1 => n25614, A2 => n19824, B1 => n25938, B2 => 
                           n25606, ZN => n6643);
   U19984 : OAI22_X1 port map( A1 => n25614, A2 => n19823, B1 => n25941, B2 => 
                           n25606, ZN => n6644);
   U19985 : OAI22_X1 port map( A1 => n25614, A2 => n19822, B1 => n25944, B2 => 
                           n25606, ZN => n6645);
   U19986 : OAI22_X1 port map( A1 => n25614, A2 => n19821, B1 => n25947, B2 => 
                           n25606, ZN => n6646);
   U19987 : OAI22_X1 port map( A1 => n25614, A2 => n19820, B1 => n25950, B2 => 
                           n25606, ZN => n6647);
   U19988 : OAI22_X1 port map( A1 => n25614, A2 => n19819, B1 => n25953, B2 => 
                           n25606, ZN => n6648);
   U19989 : OAI22_X1 port map( A1 => n25614, A2 => n19818, B1 => n25956, B2 => 
                           n25606, ZN => n6649);
   U19990 : OAI22_X1 port map( A1 => n25614, A2 => n19817, B1 => n25959, B2 => 
                           n25606, ZN => n6650);
   U19991 : OAI22_X1 port map( A1 => n25662, A2 => n19812, B1 => n25781, B2 => 
                           n25654, ZN => n6847);
   U19992 : OAI22_X1 port map( A1 => n25662, A2 => n19811, B1 => n25784, B2 => 
                           n25654, ZN => n6848);
   U19993 : OAI22_X1 port map( A1 => n25662, A2 => n19810, B1 => n25787, B2 => 
                           n25654, ZN => n6849);
   U19994 : OAI22_X1 port map( A1 => n25662, A2 => n19809, B1 => n25790, B2 => 
                           n25654, ZN => n6850);
   U19995 : OAI22_X1 port map( A1 => n25662, A2 => n19808, B1 => n25793, B2 => 
                           n25654, ZN => n6851);
   U19996 : OAI22_X1 port map( A1 => n25662, A2 => n19807, B1 => n25796, B2 => 
                           n25654, ZN => n6852);
   U19997 : OAI22_X1 port map( A1 => n25662, A2 => n19806, B1 => n25799, B2 => 
                           n25654, ZN => n6853);
   U19998 : OAI22_X1 port map( A1 => n25662, A2 => n19805, B1 => n25802, B2 => 
                           n25654, ZN => n6854);
   U19999 : OAI22_X1 port map( A1 => n25662, A2 => n19804, B1 => n25805, B2 => 
                           n25654, ZN => n6855);
   U20000 : OAI22_X1 port map( A1 => n25662, A2 => n19803, B1 => n25808, B2 => 
                           n25654, ZN => n6856);
   U20001 : OAI22_X1 port map( A1 => n25662, A2 => n19802, B1 => n25811, B2 => 
                           n25654, ZN => n6857);
   U20002 : OAI22_X1 port map( A1 => n25662, A2 => n19801, B1 => n25814, B2 => 
                           n25654, ZN => n6858);
   U20003 : OAI22_X1 port map( A1 => n25663, A2 => n19800, B1 => n25817, B2 => 
                           n25655, ZN => n6859);
   U20004 : OAI22_X1 port map( A1 => n25663, A2 => n19799, B1 => n25820, B2 => 
                           n25655, ZN => n6860);
   U20005 : OAI22_X1 port map( A1 => n25663, A2 => n19798, B1 => n25823, B2 => 
                           n25655, ZN => n6861);
   U20006 : OAI22_X1 port map( A1 => n25663, A2 => n19797, B1 => n25826, B2 => 
                           n25655, ZN => n6862);
   U20007 : OAI22_X1 port map( A1 => n25663, A2 => n19796, B1 => n25829, B2 => 
                           n25655, ZN => n6863);
   U20008 : OAI22_X1 port map( A1 => n25663, A2 => n19795, B1 => n25832, B2 => 
                           n25655, ZN => n6864);
   U20009 : OAI22_X1 port map( A1 => n25663, A2 => n19794, B1 => n25835, B2 => 
                           n25655, ZN => n6865);
   U20010 : OAI22_X1 port map( A1 => n25663, A2 => n19793, B1 => n25838, B2 => 
                           n25655, ZN => n6866);
   U20011 : OAI22_X1 port map( A1 => n25663, A2 => n19792, B1 => n25841, B2 => 
                           n25655, ZN => n6867);
   U20012 : OAI22_X1 port map( A1 => n25663, A2 => n19791, B1 => n25844, B2 => 
                           n25655, ZN => n6868);
   U20013 : OAI22_X1 port map( A1 => n25663, A2 => n19790, B1 => n25847, B2 => 
                           n25655, ZN => n6869);
   U20014 : OAI22_X1 port map( A1 => n25663, A2 => n19789, B1 => n25850, B2 => 
                           n25655, ZN => n6870);
   U20015 : OAI22_X1 port map( A1 => n25663, A2 => n19788, B1 => n25853, B2 => 
                           n25656, ZN => n6871);
   U20016 : OAI22_X1 port map( A1 => n25664, A2 => n19787, B1 => n25856, B2 => 
                           n25656, ZN => n6872);
   U20017 : OAI22_X1 port map( A1 => n25664, A2 => n19786, B1 => n25859, B2 => 
                           n25656, ZN => n6873);
   U20018 : OAI22_X1 port map( A1 => n25664, A2 => n19785, B1 => n25862, B2 => 
                           n25656, ZN => n6874);
   U20019 : OAI22_X1 port map( A1 => n25664, A2 => n19784, B1 => n25865, B2 => 
                           n25656, ZN => n6875);
   U20020 : OAI22_X1 port map( A1 => n25664, A2 => n19783, B1 => n25868, B2 => 
                           n25656, ZN => n6876);
   U20021 : OAI22_X1 port map( A1 => n25664, A2 => n19782, B1 => n25871, B2 => 
                           n25656, ZN => n6877);
   U20022 : OAI22_X1 port map( A1 => n25664, A2 => n19781, B1 => n25874, B2 => 
                           n25656, ZN => n6878);
   U20023 : OAI22_X1 port map( A1 => n25664, A2 => n19780, B1 => n25877, B2 => 
                           n25656, ZN => n6879);
   U20024 : OAI22_X1 port map( A1 => n25664, A2 => n19779, B1 => n25880, B2 => 
                           n25656, ZN => n6880);
   U20025 : OAI22_X1 port map( A1 => n25664, A2 => n19778, B1 => n25883, B2 => 
                           n25656, ZN => n6881);
   U20026 : OAI22_X1 port map( A1 => n25664, A2 => n19777, B1 => n25886, B2 => 
                           n25656, ZN => n6882);
   U20027 : OAI22_X1 port map( A1 => n25664, A2 => n19776, B1 => n25889, B2 => 
                           n25657, ZN => n6883);
   U20028 : OAI22_X1 port map( A1 => n25664, A2 => n19775, B1 => n25892, B2 => 
                           n25657, ZN => n6884);
   U20029 : OAI22_X1 port map( A1 => n25665, A2 => n19774, B1 => n25895, B2 => 
                           n25657, ZN => n6885);
   U20030 : OAI22_X1 port map( A1 => n25665, A2 => n19773, B1 => n25898, B2 => 
                           n25657, ZN => n6886);
   U20031 : OAI22_X1 port map( A1 => n25665, A2 => n19772, B1 => n25901, B2 => 
                           n25657, ZN => n6887);
   U20032 : OAI22_X1 port map( A1 => n25665, A2 => n19771, B1 => n25904, B2 => 
                           n25657, ZN => n6888);
   U20033 : OAI22_X1 port map( A1 => n25665, A2 => n19770, B1 => n25907, B2 => 
                           n25657, ZN => n6889);
   U20034 : OAI22_X1 port map( A1 => n25665, A2 => n19769, B1 => n25910, B2 => 
                           n25657, ZN => n6890);
   U20035 : OAI22_X1 port map( A1 => n25665, A2 => n19768, B1 => n25913, B2 => 
                           n25657, ZN => n6891);
   U20036 : OAI22_X1 port map( A1 => n25665, A2 => n19767, B1 => n25916, B2 => 
                           n25657, ZN => n6892);
   U20037 : OAI22_X1 port map( A1 => n25665, A2 => n19766, B1 => n25919, B2 => 
                           n25657, ZN => n6893);
   U20038 : OAI22_X1 port map( A1 => n25665, A2 => n19765, B1 => n25922, B2 => 
                           n25657, ZN => n6894);
   U20039 : OAI22_X1 port map( A1 => n25665, A2 => n19764, B1 => n25925, B2 => 
                           n25658, ZN => n6895);
   U20040 : OAI22_X1 port map( A1 => n25665, A2 => n19763, B1 => n25928, B2 => 
                           n25658, ZN => n6896);
   U20041 : OAI22_X1 port map( A1 => n25665, A2 => n19762, B1 => n25931, B2 => 
                           n25658, ZN => n6897);
   U20042 : OAI22_X1 port map( A1 => n25666, A2 => n19761, B1 => n25934, B2 => 
                           n25658, ZN => n6898);
   U20043 : OAI22_X1 port map( A1 => n25666, A2 => n19760, B1 => n25937, B2 => 
                           n25658, ZN => n6899);
   U20044 : OAI22_X1 port map( A1 => n25666, A2 => n19759, B1 => n25940, B2 => 
                           n25658, ZN => n6900);
   U20045 : OAI22_X1 port map( A1 => n25666, A2 => n19758, B1 => n25943, B2 => 
                           n25658, ZN => n6901);
   U20046 : OAI22_X1 port map( A1 => n25666, A2 => n19757, B1 => n25946, B2 => 
                           n25658, ZN => n6902);
   U20047 : OAI22_X1 port map( A1 => n25666, A2 => n19756, B1 => n25949, B2 => 
                           n25658, ZN => n6903);
   U20048 : OAI22_X1 port map( A1 => n25666, A2 => n19755, B1 => n25952, B2 => 
                           n25658, ZN => n6904);
   U20049 : OAI22_X1 port map( A1 => n25666, A2 => n19754, B1 => n25955, B2 => 
                           n25658, ZN => n6905);
   U20050 : OAI22_X1 port map( A1 => n25666, A2 => n19753, B1 => n25958, B2 => 
                           n25658, ZN => n6906);
   U20051 : OAI22_X1 port map( A1 => n25713, A2 => n19621, B1 => n25781, B2 => 
                           n25705, ZN => n7103);
   U20052 : OAI22_X1 port map( A1 => n25713, A2 => n19620, B1 => n25784, B2 => 
                           n25705, ZN => n7104);
   U20053 : OAI22_X1 port map( A1 => n25713, A2 => n19619, B1 => n25787, B2 => 
                           n25705, ZN => n7105);
   U20054 : OAI22_X1 port map( A1 => n25713, A2 => n19618, B1 => n25790, B2 => 
                           n25705, ZN => n7106);
   U20055 : OAI22_X1 port map( A1 => n25713, A2 => n19617, B1 => n25793, B2 => 
                           n25705, ZN => n7107);
   U20056 : OAI22_X1 port map( A1 => n25713, A2 => n19616, B1 => n25796, B2 => 
                           n25705, ZN => n7108);
   U20057 : OAI22_X1 port map( A1 => n25713, A2 => n19615, B1 => n25799, B2 => 
                           n25705, ZN => n7109);
   U20058 : OAI22_X1 port map( A1 => n25713, A2 => n19614, B1 => n25802, B2 => 
                           n25705, ZN => n7110);
   U20059 : OAI22_X1 port map( A1 => n25713, A2 => n19613, B1 => n25805, B2 => 
                           n25705, ZN => n7111);
   U20060 : OAI22_X1 port map( A1 => n25713, A2 => n19612, B1 => n25808, B2 => 
                           n25705, ZN => n7112);
   U20061 : OAI22_X1 port map( A1 => n25713, A2 => n19611, B1 => n25811, B2 => 
                           n25705, ZN => n7113);
   U20062 : OAI22_X1 port map( A1 => n25713, A2 => n19610, B1 => n25814, B2 => 
                           n25705, ZN => n7114);
   U20063 : OAI22_X1 port map( A1 => n25714, A2 => n19609, B1 => n25817, B2 => 
                           n25706, ZN => n7115);
   U20064 : OAI22_X1 port map( A1 => n25714, A2 => n19608, B1 => n25820, B2 => 
                           n25706, ZN => n7116);
   U20065 : OAI22_X1 port map( A1 => n25714, A2 => n19607, B1 => n25823, B2 => 
                           n25706, ZN => n7117);
   U20066 : OAI22_X1 port map( A1 => n25714, A2 => n19606, B1 => n25826, B2 => 
                           n25706, ZN => n7118);
   U20067 : OAI22_X1 port map( A1 => n25714, A2 => n19605, B1 => n25829, B2 => 
                           n25706, ZN => n7119);
   U20068 : OAI22_X1 port map( A1 => n25714, A2 => n19604, B1 => n25832, B2 => 
                           n25706, ZN => n7120);
   U20069 : OAI22_X1 port map( A1 => n25714, A2 => n19603, B1 => n25835, B2 => 
                           n25706, ZN => n7121);
   U20070 : OAI22_X1 port map( A1 => n25714, A2 => n19602, B1 => n25838, B2 => 
                           n25706, ZN => n7122);
   U20071 : OAI22_X1 port map( A1 => n25714, A2 => n19601, B1 => n25841, B2 => 
                           n25706, ZN => n7123);
   U20072 : OAI22_X1 port map( A1 => n25714, A2 => n19600, B1 => n25844, B2 => 
                           n25706, ZN => n7124);
   U20073 : OAI22_X1 port map( A1 => n25714, A2 => n19599, B1 => n25847, B2 => 
                           n25706, ZN => n7125);
   U20074 : OAI22_X1 port map( A1 => n25714, A2 => n19598, B1 => n25850, B2 => 
                           n25706, ZN => n7126);
   U20075 : OAI22_X1 port map( A1 => n25714, A2 => n19597, B1 => n25853, B2 => 
                           n25707, ZN => n7127);
   U20076 : OAI22_X1 port map( A1 => n25715, A2 => n19596, B1 => n25856, B2 => 
                           n25707, ZN => n7128);
   U20077 : OAI22_X1 port map( A1 => n25715, A2 => n19595, B1 => n25859, B2 => 
                           n25707, ZN => n7129);
   U20078 : OAI22_X1 port map( A1 => n25715, A2 => n19594, B1 => n25862, B2 => 
                           n25707, ZN => n7130);
   U20079 : OAI22_X1 port map( A1 => n25715, A2 => n19593, B1 => n25865, B2 => 
                           n25707, ZN => n7131);
   U20080 : OAI22_X1 port map( A1 => n25715, A2 => n19592, B1 => n25868, B2 => 
                           n25707, ZN => n7132);
   U20081 : OAI22_X1 port map( A1 => n25715, A2 => n19591, B1 => n25871, B2 => 
                           n25707, ZN => n7133);
   U20082 : OAI22_X1 port map( A1 => n25715, A2 => n19590, B1 => n25874, B2 => 
                           n25707, ZN => n7134);
   U20083 : OAI22_X1 port map( A1 => n25715, A2 => n19589, B1 => n25877, B2 => 
                           n25707, ZN => n7135);
   U20084 : OAI22_X1 port map( A1 => n25715, A2 => n19588, B1 => n25880, B2 => 
                           n25707, ZN => n7136);
   U20085 : OAI22_X1 port map( A1 => n25715, A2 => n19587, B1 => n25883, B2 => 
                           n25707, ZN => n7137);
   U20086 : OAI22_X1 port map( A1 => n25715, A2 => n19586, B1 => n25886, B2 => 
                           n25707, ZN => n7138);
   U20087 : OAI22_X1 port map( A1 => n25715, A2 => n19585, B1 => n25889, B2 => 
                           n25708, ZN => n7139);
   U20088 : OAI22_X1 port map( A1 => n25715, A2 => n19584, B1 => n25892, B2 => 
                           n25708, ZN => n7140);
   U20089 : OAI22_X1 port map( A1 => n25716, A2 => n19583, B1 => n25895, B2 => 
                           n25708, ZN => n7141);
   U20090 : OAI22_X1 port map( A1 => n25716, A2 => n19582, B1 => n25898, B2 => 
                           n25708, ZN => n7142);
   U20091 : OAI22_X1 port map( A1 => n25716, A2 => n19581, B1 => n25901, B2 => 
                           n25708, ZN => n7143);
   U20092 : OAI22_X1 port map( A1 => n25716, A2 => n19580, B1 => n25904, B2 => 
                           n25708, ZN => n7144);
   U20093 : OAI22_X1 port map( A1 => n25716, A2 => n19579, B1 => n25907, B2 => 
                           n25708, ZN => n7145);
   U20094 : OAI22_X1 port map( A1 => n25716, A2 => n19578, B1 => n25910, B2 => 
                           n25708, ZN => n7146);
   U20095 : OAI22_X1 port map( A1 => n25716, A2 => n19577, B1 => n25913, B2 => 
                           n25708, ZN => n7147);
   U20096 : OAI22_X1 port map( A1 => n25716, A2 => n19576, B1 => n25916, B2 => 
                           n25708, ZN => n7148);
   U20097 : OAI22_X1 port map( A1 => n25716, A2 => n19575, B1 => n25919, B2 => 
                           n25708, ZN => n7149);
   U20098 : OAI22_X1 port map( A1 => n25716, A2 => n19574, B1 => n25922, B2 => 
                           n25708, ZN => n7150);
   U20099 : OAI22_X1 port map( A1 => n25716, A2 => n19573, B1 => n25925, B2 => 
                           n25709, ZN => n7151);
   U20100 : OAI22_X1 port map( A1 => n25716, A2 => n19572, B1 => n25928, B2 => 
                           n25709, ZN => n7152);
   U20101 : OAI22_X1 port map( A1 => n25716, A2 => n19571, B1 => n25931, B2 => 
                           n25709, ZN => n7153);
   U20102 : OAI22_X1 port map( A1 => n25717, A2 => n19570, B1 => n25934, B2 => 
                           n25709, ZN => n7154);
   U20103 : OAI22_X1 port map( A1 => n25717, A2 => n19569, B1 => n25937, B2 => 
                           n25709, ZN => n7155);
   U20104 : OAI22_X1 port map( A1 => n25717, A2 => n19568, B1 => n25940, B2 => 
                           n25709, ZN => n7156);
   U20105 : OAI22_X1 port map( A1 => n25717, A2 => n19567, B1 => n25943, B2 => 
                           n25709, ZN => n7157);
   U20106 : OAI22_X1 port map( A1 => n25717, A2 => n19566, B1 => n25946, B2 => 
                           n25709, ZN => n7158);
   U20107 : OAI22_X1 port map( A1 => n25717, A2 => n19565, B1 => n25949, B2 => 
                           n25709, ZN => n7159);
   U20108 : OAI22_X1 port map( A1 => n25717, A2 => n19564, B1 => n25952, B2 => 
                           n25709, ZN => n7160);
   U20109 : OAI22_X1 port map( A1 => n25717, A2 => n19563, B1 => n25955, B2 => 
                           n25709, ZN => n7161);
   U20110 : OAI22_X1 port map( A1 => n25717, A2 => n19562, B1 => n25958, B2 => 
                           n25709, ZN => n7162);
   U20111 : NOR3_X1 port map( A1 => n19492, A2 => n25046, A3 => n19491, ZN => 
                           n23928);
   U20112 : NOR3_X1 port map( A1 => n19487, A2 => n25244, A3 => n19486, ZN => 
                           n22731);
   U20113 : OAI21_X1 port map( B1 => n21490, B2 => n21512, A => n25974, ZN => 
                           n21517);
   U20114 : OAI21_X1 port map( B1 => n21484, B2 => n21531, A => n25974, ZN => 
                           n21532);
   U20115 : OAI21_X1 port map( B1 => n21490, B2 => n21494, A => n25973, ZN => 
                           n21499);
   U20116 : OAI21_X1 port map( B1 => n21480, B2 => n21487, A => n25973, ZN => 
                           n21485);
   U20117 : BUF_X1 port map( A => n22788, Z => n25046);
   U20118 : BUF_X1 port map( A => n21591, Z => n25244);
   U20119 : BUF_X1 port map( A => n22788, Z => n25049);
   U20120 : BUF_X1 port map( A => n22788, Z => n25048);
   U20121 : BUF_X1 port map( A => n22788, Z => n25047);
   U20122 : BUF_X1 port map( A => n21591, Z => n25247);
   U20123 : BUF_X1 port map( A => n21591, Z => n25245);
   U20124 : BUF_X1 port map( A => n21591, Z => n25246);
   U20125 : NOR3_X1 port map( A1 => n19489, A2 => n19493, A3 => n19490, ZN => 
                           n23946);
   U20126 : NOR3_X1 port map( A1 => n19484, A2 => n19488, A3 => n19485, ZN => 
                           n22749);
   U20127 : NAND2_X1 port map( A1 => n23930, A2 => n23937, ZN => n22770);
   U20128 : NAND2_X1 port map( A1 => n23930, A2 => n23940, ZN => n22800);
   U20129 : NAND2_X1 port map( A1 => n22733, A2 => n22740, ZN => n21573);
   U20130 : NAND2_X1 port map( A1 => n22733, A2 => n22743, ZN => n21603);
   U20131 : NAND2_X1 port map( A1 => n19482, A2 => n19483, ZN => n21481);
   U20132 : BUF_X1 port map( A => n19478, Z => n25974);
   U20133 : BUF_X1 port map( A => n19478, Z => n25973);
   U20134 : BUF_X1 port map( A => n19478, Z => n25975);
   U20135 : NAND2_X1 port map( A1 => n23930, A2 => n23935, ZN => n22774);
   U20136 : NAND2_X1 port map( A1 => n22733, A2 => n22738, ZN => n21577);
   U20137 : BUF_X1 port map( A => n19478, Z => n25976);
   U20138 : BUF_X1 port map( A => n19478, Z => n25977);
   U20139 : NAND2_X1 port map( A1 => n23929, A2 => n23930, ZN => n22760);
   U20140 : NAND2_X1 port map( A1 => n23927, A2 => n23930, ZN => n22765);
   U20141 : NAND2_X1 port map( A1 => n23933, A2 => n23930, ZN => n22795);
   U20142 : NAND2_X1 port map( A1 => n22732, A2 => n22733, ZN => n21563);
   U20143 : NAND2_X1 port map( A1 => n22730, A2 => n22733, ZN => n21568);
   U20144 : NAND2_X1 port map( A1 => n22736, A2 => n22733, ZN => n21598);
   U20145 : NAND2_X1 port map( A1 => n23934, A2 => n23939, ZN => n22784);
   U20146 : NAND2_X1 port map( A1 => n23934, A2 => n23940, ZN => n22799);
   U20147 : NAND2_X1 port map( A1 => n22737, A2 => n22742, ZN => n21587);
   U20148 : NAND2_X1 port map( A1 => n22737, A2 => n22743, ZN => n21602);
   U20149 : NAND2_X1 port map( A1 => n23931, A2 => n23940, ZN => n22794);
   U20150 : NAND2_X1 port map( A1 => n22734, A2 => n22743, ZN => n21597);
   U20151 : NAND2_X1 port map( A1 => n23933, A2 => n23934, ZN => n22790);
   U20152 : NAND2_X1 port map( A1 => n23946, A2 => n23934, ZN => n22785);
   U20153 : NAND2_X1 port map( A1 => n22736, A2 => n22737, ZN => n21593);
   U20154 : NAND2_X1 port map( A1 => n22749, A2 => n22737, ZN => n21588);
   U20155 : NAND2_X1 port map( A1 => n23937, A2 => n23931, ZN => n22775);
   U20156 : NAND2_X1 port map( A1 => n22740, A2 => n22734, ZN => n21578);
   U20157 : BUF_X1 port map( A => n19557, Z => n25782);
   U20158 : BUF_X1 port map( A => n19556, Z => n25785);
   U20159 : BUF_X1 port map( A => n19555, Z => n25788);
   U20160 : BUF_X1 port map( A => n19554, Z => n25791);
   U20161 : BUF_X1 port map( A => n19553, Z => n25794);
   U20162 : BUF_X1 port map( A => n19552, Z => n25797);
   U20163 : BUF_X1 port map( A => n19551, Z => n25800);
   U20164 : BUF_X1 port map( A => n19550, Z => n25803);
   U20165 : BUF_X1 port map( A => n19549, Z => n25806);
   U20166 : BUF_X1 port map( A => n19548, Z => n25809);
   U20167 : BUF_X1 port map( A => n19547, Z => n25812);
   U20168 : BUF_X1 port map( A => n19546, Z => n25815);
   U20169 : BUF_X1 port map( A => n19545, Z => n25818);
   U20170 : BUF_X1 port map( A => n19544, Z => n25821);
   U20171 : BUF_X1 port map( A => n19543, Z => n25824);
   U20172 : BUF_X1 port map( A => n19542, Z => n25827);
   U20173 : BUF_X1 port map( A => n19541, Z => n25830);
   U20174 : BUF_X1 port map( A => n19540, Z => n25833);
   U20175 : BUF_X1 port map( A => n19539, Z => n25836);
   U20176 : BUF_X1 port map( A => n19538, Z => n25839);
   U20177 : BUF_X1 port map( A => n19537, Z => n25842);
   U20178 : BUF_X1 port map( A => n19536, Z => n25845);
   U20179 : BUF_X1 port map( A => n19535, Z => n25848);
   U20180 : BUF_X1 port map( A => n19534, Z => n25851);
   U20181 : BUF_X1 port map( A => n19533, Z => n25854);
   U20182 : BUF_X1 port map( A => n19532, Z => n25857);
   U20183 : BUF_X1 port map( A => n19531, Z => n25860);
   U20184 : BUF_X1 port map( A => n19530, Z => n25863);
   U20185 : BUF_X1 port map( A => n19529, Z => n25866);
   U20186 : BUF_X1 port map( A => n19528, Z => n25869);
   U20187 : BUF_X1 port map( A => n19527, Z => n25872);
   U20188 : BUF_X1 port map( A => n19526, Z => n25875);
   U20189 : BUF_X1 port map( A => n19525, Z => n25878);
   U20190 : BUF_X1 port map( A => n19524, Z => n25881);
   U20191 : BUF_X1 port map( A => n19523, Z => n25884);
   U20192 : BUF_X1 port map( A => n19522, Z => n25887);
   U20193 : BUF_X1 port map( A => n19521, Z => n25890);
   U20194 : BUF_X1 port map( A => n19520, Z => n25893);
   U20195 : BUF_X1 port map( A => n19519, Z => n25896);
   U20196 : BUF_X1 port map( A => n19518, Z => n25899);
   U20197 : BUF_X1 port map( A => n19517, Z => n25902);
   U20198 : BUF_X1 port map( A => n19516, Z => n25905);
   U20199 : BUF_X1 port map( A => n19515, Z => n25908);
   U20200 : BUF_X1 port map( A => n19514, Z => n25911);
   U20201 : BUF_X1 port map( A => n19513, Z => n25914);
   U20202 : BUF_X1 port map( A => n19512, Z => n25917);
   U20203 : BUF_X1 port map( A => n19511, Z => n25920);
   U20204 : BUF_X1 port map( A => n19510, Z => n25923);
   U20205 : BUF_X1 port map( A => n19509, Z => n25926);
   U20206 : BUF_X1 port map( A => n19508, Z => n25929);
   U20207 : BUF_X1 port map( A => n19507, Z => n25932);
   U20208 : BUF_X1 port map( A => n19506, Z => n25935);
   U20209 : BUF_X1 port map( A => n19505, Z => n25938);
   U20210 : BUF_X1 port map( A => n19504, Z => n25941);
   U20211 : BUF_X1 port map( A => n19503, Z => n25944);
   U20212 : BUF_X1 port map( A => n19502, Z => n25947);
   U20213 : BUF_X1 port map( A => n19501, Z => n25950);
   U20214 : BUF_X1 port map( A => n19500, Z => n25953);
   U20215 : BUF_X1 port map( A => n19499, Z => n25956);
   U20216 : BUF_X1 port map( A => n19498, Z => n25959);
   U20217 : BUF_X1 port map( A => n19497, Z => n25962);
   U20218 : BUF_X1 port map( A => n19496, Z => n25965);
   U20219 : BUF_X1 port map( A => n19495, Z => n25968);
   U20220 : BUF_X1 port map( A => n19494, Z => n25971);
   U20221 : BUF_X1 port map( A => n22788, Z => n25050);
   U20222 : BUF_X1 port map( A => n21591, Z => n25248);
   U20223 : BUF_X1 port map( A => n19557, Z => n25781);
   U20224 : BUF_X1 port map( A => n19556, Z => n25784);
   U20225 : BUF_X1 port map( A => n19555, Z => n25787);
   U20226 : BUF_X1 port map( A => n19554, Z => n25790);
   U20227 : BUF_X1 port map( A => n19553, Z => n25793);
   U20228 : BUF_X1 port map( A => n19552, Z => n25796);
   U20229 : BUF_X1 port map( A => n19551, Z => n25799);
   U20230 : BUF_X1 port map( A => n19550, Z => n25802);
   U20231 : BUF_X1 port map( A => n19549, Z => n25805);
   U20232 : BUF_X1 port map( A => n19548, Z => n25808);
   U20233 : BUF_X1 port map( A => n19547, Z => n25811);
   U20234 : BUF_X1 port map( A => n19546, Z => n25814);
   U20235 : BUF_X1 port map( A => n19545, Z => n25817);
   U20236 : BUF_X1 port map( A => n19544, Z => n25820);
   U20237 : BUF_X1 port map( A => n19543, Z => n25823);
   U20238 : BUF_X1 port map( A => n19542, Z => n25826);
   U20239 : BUF_X1 port map( A => n19541, Z => n25829);
   U20240 : BUF_X1 port map( A => n19540, Z => n25832);
   U20241 : BUF_X1 port map( A => n19539, Z => n25835);
   U20242 : BUF_X1 port map( A => n19538, Z => n25838);
   U20243 : BUF_X1 port map( A => n19537, Z => n25841);
   U20244 : BUF_X1 port map( A => n19536, Z => n25844);
   U20245 : BUF_X1 port map( A => n19535, Z => n25847);
   U20246 : BUF_X1 port map( A => n19534, Z => n25850);
   U20247 : BUF_X1 port map( A => n19533, Z => n25853);
   U20248 : BUF_X1 port map( A => n19532, Z => n25856);
   U20249 : BUF_X1 port map( A => n19531, Z => n25859);
   U20250 : BUF_X1 port map( A => n19530, Z => n25862);
   U20251 : BUF_X1 port map( A => n19529, Z => n25865);
   U20252 : BUF_X1 port map( A => n19528, Z => n25868);
   U20253 : BUF_X1 port map( A => n19527, Z => n25871);
   U20254 : BUF_X1 port map( A => n19526, Z => n25874);
   U20255 : BUF_X1 port map( A => n19525, Z => n25877);
   U20256 : BUF_X1 port map( A => n19524, Z => n25880);
   U20257 : BUF_X1 port map( A => n19523, Z => n25883);
   U20258 : BUF_X1 port map( A => n19522, Z => n25886);
   U20259 : BUF_X1 port map( A => n19521, Z => n25889);
   U20260 : BUF_X1 port map( A => n19520, Z => n25892);
   U20261 : BUF_X1 port map( A => n19519, Z => n25895);
   U20262 : BUF_X1 port map( A => n19518, Z => n25898);
   U20263 : BUF_X1 port map( A => n19517, Z => n25901);
   U20264 : BUF_X1 port map( A => n19516, Z => n25904);
   U20265 : BUF_X1 port map( A => n19515, Z => n25907);
   U20266 : BUF_X1 port map( A => n19514, Z => n25910);
   U20267 : BUF_X1 port map( A => n19513, Z => n25913);
   U20268 : BUF_X1 port map( A => n19512, Z => n25916);
   U20269 : BUF_X1 port map( A => n19511, Z => n25919);
   U20270 : BUF_X1 port map( A => n19510, Z => n25922);
   U20271 : BUF_X1 port map( A => n19509, Z => n25925);
   U20272 : BUF_X1 port map( A => n19508, Z => n25928);
   U20273 : BUF_X1 port map( A => n19507, Z => n25931);
   U20274 : BUF_X1 port map( A => n19506, Z => n25934);
   U20275 : BUF_X1 port map( A => n19505, Z => n25937);
   U20276 : BUF_X1 port map( A => n19504, Z => n25940);
   U20277 : BUF_X1 port map( A => n19503, Z => n25943);
   U20278 : BUF_X1 port map( A => n19502, Z => n25946);
   U20279 : BUF_X1 port map( A => n19501, Z => n25949);
   U20280 : BUF_X1 port map( A => n19500, Z => n25952);
   U20281 : BUF_X1 port map( A => n19499, Z => n25955);
   U20282 : BUF_X1 port map( A => n19498, Z => n25958);
   U20283 : BUF_X1 port map( A => n19497, Z => n25961);
   U20284 : BUF_X1 port map( A => n19496, Z => n25964);
   U20285 : BUF_X1 port map( A => n19495, Z => n25967);
   U20286 : BUF_X1 port map( A => n19494, Z => n25970);
   U20287 : NAND2_X1 port map( A1 => n23946, A2 => n23930, ZN => n22789);
   U20288 : NAND2_X1 port map( A1 => n22749, A2 => n22733, ZN => n21592);
   U20289 : NAND2_X1 port map( A1 => n23929, A2 => n23934, ZN => n22769);
   U20290 : NAND2_X1 port map( A1 => n22732, A2 => n22737, ZN => n21572);
   U20291 : NAND2_X1 port map( A1 => n23929, A2 => n23931, ZN => n22759);
   U20292 : NAND2_X1 port map( A1 => n23935, A2 => n23931, ZN => n22764);
   U20293 : NAND2_X1 port map( A1 => n22732, A2 => n22734, ZN => n21562);
   U20294 : NAND2_X1 port map( A1 => n22738, A2 => n22734, ZN => n21567);
   U20295 : OAI21_X1 port map( B1 => n21480, B2 => n21484, A => n25973, ZN => 
                           n21482);
   U20296 : OAI21_X1 port map( B1 => n21480, B2 => n21490, A => n25973, ZN => 
                           n21488);
   U20297 : BUF_X1 port map( A => n19557, Z => n25783);
   U20298 : BUF_X1 port map( A => n19556, Z => n25786);
   U20299 : BUF_X1 port map( A => n19555, Z => n25789);
   U20300 : BUF_X1 port map( A => n19554, Z => n25792);
   U20301 : BUF_X1 port map( A => n19553, Z => n25795);
   U20302 : BUF_X1 port map( A => n19552, Z => n25798);
   U20303 : BUF_X1 port map( A => n19551, Z => n25801);
   U20304 : BUF_X1 port map( A => n19550, Z => n25804);
   U20305 : BUF_X1 port map( A => n19549, Z => n25807);
   U20306 : BUF_X1 port map( A => n19548, Z => n25810);
   U20307 : BUF_X1 port map( A => n19547, Z => n25813);
   U20308 : BUF_X1 port map( A => n19546, Z => n25816);
   U20309 : BUF_X1 port map( A => n19545, Z => n25819);
   U20310 : BUF_X1 port map( A => n19544, Z => n25822);
   U20311 : BUF_X1 port map( A => n19543, Z => n25825);
   U20312 : BUF_X1 port map( A => n19542, Z => n25828);
   U20313 : BUF_X1 port map( A => n19541, Z => n25831);
   U20314 : BUF_X1 port map( A => n19540, Z => n25834);
   U20315 : BUF_X1 port map( A => n19539, Z => n25837);
   U20316 : BUF_X1 port map( A => n19538, Z => n25840);
   U20317 : BUF_X1 port map( A => n19537, Z => n25843);
   U20318 : BUF_X1 port map( A => n19536, Z => n25846);
   U20319 : BUF_X1 port map( A => n19535, Z => n25849);
   U20320 : BUF_X1 port map( A => n19534, Z => n25852);
   U20321 : BUF_X1 port map( A => n19533, Z => n25855);
   U20322 : BUF_X1 port map( A => n19532, Z => n25858);
   U20323 : BUF_X1 port map( A => n19531, Z => n25861);
   U20324 : BUF_X1 port map( A => n19530, Z => n25864);
   U20325 : BUF_X1 port map( A => n19529, Z => n25867);
   U20326 : BUF_X1 port map( A => n19528, Z => n25870);
   U20327 : BUF_X1 port map( A => n19527, Z => n25873);
   U20328 : BUF_X1 port map( A => n19526, Z => n25876);
   U20329 : BUF_X1 port map( A => n19525, Z => n25879);
   U20330 : BUF_X1 port map( A => n19524, Z => n25882);
   U20331 : BUF_X1 port map( A => n19523, Z => n25885);
   U20332 : BUF_X1 port map( A => n19522, Z => n25888);
   U20333 : BUF_X1 port map( A => n19521, Z => n25891);
   U20334 : BUF_X1 port map( A => n19520, Z => n25894);
   U20335 : BUF_X1 port map( A => n19519, Z => n25897);
   U20336 : BUF_X1 port map( A => n19518, Z => n25900);
   U20337 : BUF_X1 port map( A => n19517, Z => n25903);
   U20338 : BUF_X1 port map( A => n19516, Z => n25906);
   U20339 : BUF_X1 port map( A => n19515, Z => n25909);
   U20340 : BUF_X1 port map( A => n19514, Z => n25912);
   U20341 : BUF_X1 port map( A => n19513, Z => n25915);
   U20342 : BUF_X1 port map( A => n19512, Z => n25918);
   U20343 : BUF_X1 port map( A => n19511, Z => n25921);
   U20344 : BUF_X1 port map( A => n19510, Z => n25924);
   U20345 : BUF_X1 port map( A => n19509, Z => n25927);
   U20346 : BUF_X1 port map( A => n19508, Z => n25930);
   U20347 : BUF_X1 port map( A => n19507, Z => n25933);
   U20348 : BUF_X1 port map( A => n19506, Z => n25936);
   U20349 : BUF_X1 port map( A => n19505, Z => n25939);
   U20350 : BUF_X1 port map( A => n19504, Z => n25942);
   U20351 : BUF_X1 port map( A => n19503, Z => n25945);
   U20352 : BUF_X1 port map( A => n19502, Z => n25948);
   U20353 : BUF_X1 port map( A => n19501, Z => n25951);
   U20354 : BUF_X1 port map( A => n19500, Z => n25954);
   U20355 : BUF_X1 port map( A => n19499, Z => n25957);
   U20356 : BUF_X1 port map( A => n19498, Z => n25960);
   U20357 : BUF_X1 port map( A => n19497, Z => n25963);
   U20358 : BUF_X1 port map( A => n19496, Z => n25966);
   U20359 : BUF_X1 port map( A => n19495, Z => n25969);
   U20360 : BUF_X1 port map( A => n19494, Z => n25972);
   U20361 : OAI21_X1 port map( B1 => n21484, B2 => n21521, A => n25974, ZN => 
                           n21522);
   U20362 : OAI21_X1 port map( B1 => n21490, B2 => n21503, A => n25973, ZN => 
                           n21508);
   U20363 : OAI21_X1 port map( B1 => n21484, B2 => n21549, A => n25974, ZN => 
                           n21550);
   U20364 : OAI21_X1 port map( B1 => n21490, B2 => n21549, A => n25974, ZN => 
                           n21554);
   U20365 : OAI21_X1 port map( B1 => n21490, B2 => n21521, A => n25974, ZN => 
                           n21526);
   U20366 : OAI21_X1 port map( B1 => n21481, B2 => n21494, A => n25973, ZN => 
                           n21492);
   U20367 : OAI21_X1 port map( B1 => n21487, B2 => n21503, A => n25973, ZN => 
                           n21506);
   U20368 : OAI21_X1 port map( B1 => n21487, B2 => n21521, A => n25974, ZN => 
                           n21524);
   U20369 : OAI21_X1 port map( B1 => n21481, B2 => n21549, A => n25975, ZN => 
                           n21547);
   U20370 : OAI21_X1 port map( B1 => n21487, B2 => n21549, A => n25975, ZN => 
                           n21552);
   U20371 : OAI21_X1 port map( B1 => n21487, B2 => n21512, A => n25974, ZN => 
                           n21515);
   U20372 : OAI21_X1 port map( B1 => n21481, B2 => n21503, A => n25973, ZN => 
                           n21501);
   U20373 : OAI21_X1 port map( B1 => n21487, B2 => n21494, A => n25973, ZN => 
                           n21497);
   U20374 : OAI21_X1 port map( B1 => n21484, B2 => n21494, A => n25973, ZN => 
                           n21495);
   U20375 : OAI21_X1 port map( B1 => n21481, B2 => n21540, A => n25975, ZN => 
                           n21538);
   U20376 : OAI21_X1 port map( B1 => n21487, B2 => n21540, A => n25975, ZN => 
                           n21543);
   U20377 : OAI21_X1 port map( B1 => n21490, B2 => n21531, A => n25975, ZN => 
                           n21536);
   U20378 : OAI21_X1 port map( B1 => n21484, B2 => n21540, A => n25975, ZN => 
                           n21541);
   U20379 : OAI21_X1 port map( B1 => n21481, B2 => n21512, A => n25974, ZN => 
                           n21510);
   U20380 : OAI21_X1 port map( B1 => n21481, B2 => n21531, A => n25974, ZN => 
                           n21529);
   U20381 : OAI21_X1 port map( B1 => n21490, B2 => n21540, A => n25975, ZN => 
                           n21545);
   U20382 : OAI21_X1 port map( B1 => n21487, B2 => n21531, A => n25975, ZN => 
                           n21534);
   U20383 : OAI21_X1 port map( B1 => n21484, B2 => n21512, A => n25974, ZN => 
                           n21513);
   U20384 : OAI21_X1 port map( B1 => n21484, B2 => n21503, A => n25973, ZN => 
                           n21504);
   U20385 : AND2_X1 port map( A1 => n23930, A2 => n23939, ZN => n22787);
   U20386 : AND2_X1 port map( A1 => n22733, A2 => n22742, ZN => n21590);
   U20387 : AND2_X1 port map( A1 => n23934, A2 => n23937, ZN => n22777);
   U20388 : AND2_X1 port map( A1 => n22737, A2 => n22740, ZN => n21580);
   U20389 : AND2_X1 port map( A1 => n23935, A2 => n23934, ZN => n22773);
   U20390 : AND2_X1 port map( A1 => n23927, A2 => n23934, ZN => n22767);
   U20391 : AND2_X1 port map( A1 => n22738, A2 => n22737, ZN => n21576);
   U20392 : AND2_X1 port map( A1 => n22730, A2 => n22737, ZN => n21570);
   U20393 : AND2_X1 port map( A1 => n23939, A2 => n23931, ZN => n22779);
   U20394 : AND2_X1 port map( A1 => n23933, A2 => n23931, ZN => n22768);
   U20395 : AND2_X1 port map( A1 => n23946, A2 => n23931, ZN => n22793);
   U20396 : AND2_X1 port map( A1 => n23927, A2 => n23931, ZN => n22803);
   U20397 : AND2_X1 port map( A1 => n22742, A2 => n22734, ZN => n21582);
   U20398 : AND2_X1 port map( A1 => n22736, A2 => n22734, ZN => n21571);
   U20399 : AND2_X1 port map( A1 => n22749, A2 => n22734, ZN => n21596);
   U20400 : AND2_X1 port map( A1 => n22730, A2 => n22734, ZN => n21606);
   U20401 : AND2_X1 port map( A1 => n23928, A2 => n23940, ZN => n22778);
   U20402 : AND2_X1 port map( A1 => n22731, A2 => n22743, ZN => n21581);
   U20403 : AND2_X1 port map( A1 => n23929, A2 => n23928, ZN => n22762);
   U20404 : AND2_X1 port map( A1 => n23927, A2 => n23928, ZN => n22763);
   U20405 : AND2_X1 port map( A1 => n23935, A2 => n23928, ZN => n22772);
   U20406 : AND2_X1 port map( A1 => n23939, A2 => n23928, ZN => n22792);
   U20407 : AND2_X1 port map( A1 => n23933, A2 => n23928, ZN => n22797);
   U20408 : AND2_X1 port map( A1 => n23937, A2 => n23928, ZN => n22802);
   U20409 : AND2_X1 port map( A1 => n22732, A2 => n22731, ZN => n21565);
   U20410 : AND2_X1 port map( A1 => n22730, A2 => n22731, ZN => n21566);
   U20411 : AND2_X1 port map( A1 => n22738, A2 => n22731, ZN => n21575);
   U20412 : AND2_X1 port map( A1 => n22742, A2 => n22731, ZN => n21595);
   U20413 : AND2_X1 port map( A1 => n22736, A2 => n22731, ZN => n21600);
   U20414 : AND2_X1 port map( A1 => n22740, A2 => n22731, ZN => n21605);
   U20415 : OAI221_X1 port map( B1 => n19800, B2 => n25167, C1 => n19864, C2 =>
                           n25161, A => n23710, ZN => n23709);
   U20416 : AOI22_X1 port map( A1 => n25155, A2 => n20120, B1 => n25149, B2 => 
                           n18220, ZN => n23710);
   U20417 : OAI221_X1 port map( B1 => n19799, B2 => n25167, C1 => n19863, C2 =>
                           n25161, A => n23692, ZN => n23691);
   U20418 : AOI22_X1 port map( A1 => n25155, A2 => n20119, B1 => n25149, B2 => 
                           n18199, ZN => n23692);
   U20419 : OAI221_X1 port map( B1 => n19798, B2 => n25167, C1 => n19862, C2 =>
                           n25161, A => n23674, ZN => n23673);
   U20420 : AOI22_X1 port map( A1 => n25155, A2 => n20118, B1 => n25149, B2 => 
                           n18178, ZN => n23674);
   U20421 : OAI221_X1 port map( B1 => n19797, B2 => n25167, C1 => n19861, C2 =>
                           n25161, A => n23656, ZN => n23655);
   U20422 : AOI22_X1 port map( A1 => n25155, A2 => n20117, B1 => n25149, B2 => 
                           n18157, ZN => n23656);
   U20423 : OAI221_X1 port map( B1 => n19796, B2 => n25167, C1 => n19860, C2 =>
                           n25161, A => n23638, ZN => n23637);
   U20424 : AOI22_X1 port map( A1 => n25155, A2 => n20116, B1 => n25149, B2 => 
                           n18136, ZN => n23638);
   U20425 : OAI221_X1 port map( B1 => n19795, B2 => n25167, C1 => n19859, C2 =>
                           n25161, A => n23620, ZN => n23619);
   U20426 : AOI22_X1 port map( A1 => n25155, A2 => n20115, B1 => n25149, B2 => 
                           n18115, ZN => n23620);
   U20427 : OAI221_X1 port map( B1 => n19794, B2 => n25167, C1 => n19858, C2 =>
                           n25161, A => n23602, ZN => n23601);
   U20428 : AOI22_X1 port map( A1 => n25155, A2 => n20114, B1 => n25149, B2 => 
                           n18094, ZN => n23602);
   U20429 : OAI221_X1 port map( B1 => n19793, B2 => n25167, C1 => n19857, C2 =>
                           n25161, A => n23584, ZN => n23583);
   U20430 : AOI22_X1 port map( A1 => n25155, A2 => n20113, B1 => n25149, B2 => 
                           n18073, ZN => n23584);
   U20431 : OAI221_X1 port map( B1 => n19792, B2 => n25167, C1 => n19856, C2 =>
                           n25161, A => n23566, ZN => n23565);
   U20432 : AOI22_X1 port map( A1 => n25155, A2 => n20112, B1 => n25149, B2 => 
                           n18052, ZN => n23566);
   U20433 : OAI221_X1 port map( B1 => n19791, B2 => n25167, C1 => n19855, C2 =>
                           n25161, A => n23548, ZN => n23547);
   U20434 : AOI22_X1 port map( A1 => n25155, A2 => n20111, B1 => n25149, B2 => 
                           n18031, ZN => n23548);
   U20435 : OAI221_X1 port map( B1 => n19790, B2 => n25167, C1 => n19854, C2 =>
                           n25161, A => n23530, ZN => n23529);
   U20436 : AOI22_X1 port map( A1 => n25155, A2 => n20110, B1 => n25149, B2 => 
                           n18010, ZN => n23530);
   U20437 : OAI221_X1 port map( B1 => n19789, B2 => n25167, C1 => n19853, C2 =>
                           n25161, A => n23512, ZN => n23511);
   U20438 : AOI22_X1 port map( A1 => n25155, A2 => n20109, B1 => n25149, B2 => 
                           n17989, ZN => n23512);
   U20439 : OAI221_X1 port map( B1 => n19788, B2 => n25168, C1 => n19852, C2 =>
                           n25162, A => n23494, ZN => n23493);
   U20440 : AOI22_X1 port map( A1 => n25156, A2 => n20108, B1 => n25150, B2 => 
                           n17968, ZN => n23494);
   U20441 : OAI221_X1 port map( B1 => n19787, B2 => n25168, C1 => n19851, C2 =>
                           n25162, A => n23476, ZN => n23475);
   U20442 : AOI22_X1 port map( A1 => n25156, A2 => n20107, B1 => n25150, B2 => 
                           n17947, ZN => n23476);
   U20443 : OAI221_X1 port map( B1 => n19786, B2 => n25168, C1 => n19850, C2 =>
                           n25162, A => n23458, ZN => n23457);
   U20444 : AOI22_X1 port map( A1 => n25156, A2 => n20106, B1 => n25150, B2 => 
                           n17926, ZN => n23458);
   U20445 : OAI221_X1 port map( B1 => n19785, B2 => n25168, C1 => n19849, C2 =>
                           n25162, A => n23440, ZN => n23439);
   U20446 : AOI22_X1 port map( A1 => n25156, A2 => n20105, B1 => n25150, B2 => 
                           n17905, ZN => n23440);
   U20447 : OAI221_X1 port map( B1 => n19784, B2 => n25168, C1 => n19848, C2 =>
                           n25162, A => n23422, ZN => n23421);
   U20448 : AOI22_X1 port map( A1 => n25156, A2 => n20104, B1 => n25150, B2 => 
                           n17884, ZN => n23422);
   U20449 : OAI221_X1 port map( B1 => n19783, B2 => n25168, C1 => n19847, C2 =>
                           n25162, A => n23404, ZN => n23403);
   U20450 : AOI22_X1 port map( A1 => n25156, A2 => n20103, B1 => n25150, B2 => 
                           n17863, ZN => n23404);
   U20451 : OAI221_X1 port map( B1 => n19782, B2 => n25168, C1 => n19846, C2 =>
                           n25162, A => n23386, ZN => n23385);
   U20452 : AOI22_X1 port map( A1 => n25156, A2 => n20102, B1 => n25150, B2 => 
                           n17842, ZN => n23386);
   U20453 : OAI221_X1 port map( B1 => n19781, B2 => n25168, C1 => n19845, C2 =>
                           n25162, A => n23368, ZN => n23367);
   U20454 : AOI22_X1 port map( A1 => n25156, A2 => n20101, B1 => n25150, B2 => 
                           n17821, ZN => n23368);
   U20455 : OAI221_X1 port map( B1 => n19780, B2 => n25168, C1 => n19844, C2 =>
                           n25162, A => n23350, ZN => n23349);
   U20456 : AOI22_X1 port map( A1 => n25156, A2 => n20100, B1 => n25150, B2 => 
                           n17800, ZN => n23350);
   U20457 : OAI221_X1 port map( B1 => n19779, B2 => n25168, C1 => n19843, C2 =>
                           n25162, A => n23332, ZN => n23331);
   U20458 : AOI22_X1 port map( A1 => n25156, A2 => n20099, B1 => n25150, B2 => 
                           n17779, ZN => n23332);
   U20459 : OAI221_X1 port map( B1 => n19778, B2 => n25168, C1 => n19842, C2 =>
                           n25162, A => n23314, ZN => n23313);
   U20460 : AOI22_X1 port map( A1 => n25156, A2 => n20098, B1 => n25150, B2 => 
                           n17758, ZN => n23314);
   U20461 : OAI221_X1 port map( B1 => n19777, B2 => n25168, C1 => n19841, C2 =>
                           n25162, A => n23296, ZN => n23295);
   U20462 : AOI22_X1 port map( A1 => n25156, A2 => n20097, B1 => n25150, B2 => 
                           n17737, ZN => n23296);
   U20463 : OAI221_X1 port map( B1 => n19776, B2 => n25169, C1 => n19840, C2 =>
                           n25163, A => n23278, ZN => n23277);
   U20464 : AOI22_X1 port map( A1 => n25157, A2 => n20096, B1 => n25151, B2 => 
                           n17716, ZN => n23278);
   U20465 : OAI221_X1 port map( B1 => n19775, B2 => n25169, C1 => n19839, C2 =>
                           n25163, A => n23260, ZN => n23259);
   U20466 : AOI22_X1 port map( A1 => n25157, A2 => n20095, B1 => n25151, B2 => 
                           n17695, ZN => n23260);
   U20467 : OAI221_X1 port map( B1 => n19774, B2 => n25169, C1 => n19838, C2 =>
                           n25163, A => n23242, ZN => n23241);
   U20468 : AOI22_X1 port map( A1 => n25157, A2 => n20094, B1 => n25151, B2 => 
                           n17674, ZN => n23242);
   U20469 : OAI221_X1 port map( B1 => n19773, B2 => n25169, C1 => n19837, C2 =>
                           n25163, A => n23224, ZN => n23223);
   U20470 : AOI22_X1 port map( A1 => n25157, A2 => n20093, B1 => n25151, B2 => 
                           n17653, ZN => n23224);
   U20471 : OAI221_X1 port map( B1 => n19772, B2 => n25169, C1 => n19836, C2 =>
                           n25163, A => n23206, ZN => n23205);
   U20472 : AOI22_X1 port map( A1 => n25157, A2 => n20092, B1 => n25151, B2 => 
                           n17632, ZN => n23206);
   U20473 : OAI221_X1 port map( B1 => n19771, B2 => n25169, C1 => n19835, C2 =>
                           n25163, A => n23188, ZN => n23187);
   U20474 : AOI22_X1 port map( A1 => n25157, A2 => n20091, B1 => n25151, B2 => 
                           n17611, ZN => n23188);
   U20475 : OAI221_X1 port map( B1 => n19770, B2 => n25169, C1 => n19834, C2 =>
                           n25163, A => n23170, ZN => n23169);
   U20476 : AOI22_X1 port map( A1 => n25157, A2 => n20090, B1 => n25151, B2 => 
                           n17590, ZN => n23170);
   U20477 : OAI221_X1 port map( B1 => n19769, B2 => n25169, C1 => n19833, C2 =>
                           n25163, A => n23152, ZN => n23151);
   U20478 : AOI22_X1 port map( A1 => n25157, A2 => n20089, B1 => n25151, B2 => 
                           n17569, ZN => n23152);
   U20479 : OAI221_X1 port map( B1 => n19768, B2 => n25169, C1 => n19832, C2 =>
                           n25163, A => n23134, ZN => n23133);
   U20480 : AOI22_X1 port map( A1 => n25157, A2 => n20088, B1 => n25151, B2 => 
                           n17548, ZN => n23134);
   U20481 : OAI221_X1 port map( B1 => n19767, B2 => n25169, C1 => n19831, C2 =>
                           n25163, A => n23116, ZN => n23115);
   U20482 : AOI22_X1 port map( A1 => n25157, A2 => n20087, B1 => n25151, B2 => 
                           n17527, ZN => n23116);
   U20483 : OAI221_X1 port map( B1 => n19766, B2 => n25169, C1 => n19830, C2 =>
                           n25163, A => n23098, ZN => n23097);
   U20484 : AOI22_X1 port map( A1 => n25157, A2 => n20086, B1 => n25151, B2 => 
                           n17506, ZN => n23098);
   U20485 : OAI221_X1 port map( B1 => n19765, B2 => n25169, C1 => n19829, C2 =>
                           n25163, A => n23080, ZN => n23079);
   U20486 : AOI22_X1 port map( A1 => n25157, A2 => n20085, B1 => n25151, B2 => 
                           n17485, ZN => n23080);
   U20487 : OAI221_X1 port map( B1 => n19764, B2 => n25170, C1 => n19828, C2 =>
                           n25164, A => n23062, ZN => n23061);
   U20488 : AOI22_X1 port map( A1 => n25158, A2 => n20084, B1 => n25152, B2 => 
                           n17464, ZN => n23062);
   U20489 : OAI221_X1 port map( B1 => n19763, B2 => n25170, C1 => n19827, C2 =>
                           n25164, A => n23044, ZN => n23043);
   U20490 : AOI22_X1 port map( A1 => n25158, A2 => n20083, B1 => n25152, B2 => 
                           n17443, ZN => n23044);
   U20491 : OAI221_X1 port map( B1 => n19762, B2 => n25170, C1 => n19826, C2 =>
                           n25164, A => n23026, ZN => n23025);
   U20492 : AOI22_X1 port map( A1 => n25158, A2 => n20082, B1 => n25152, B2 => 
                           n17422, ZN => n23026);
   U20493 : OAI221_X1 port map( B1 => n19761, B2 => n25170, C1 => n19825, C2 =>
                           n25164, A => n23008, ZN => n23007);
   U20494 : AOI22_X1 port map( A1 => n25158, A2 => n20081, B1 => n25152, B2 => 
                           n17401, ZN => n23008);
   U20495 : OAI221_X1 port map( B1 => n19760, B2 => n25170, C1 => n19824, C2 =>
                           n25164, A => n22990, ZN => n22989);
   U20496 : AOI22_X1 port map( A1 => n25158, A2 => n20080, B1 => n25152, B2 => 
                           n17380, ZN => n22990);
   U20497 : OAI221_X1 port map( B1 => n19759, B2 => n25170, C1 => n19823, C2 =>
                           n25164, A => n22972, ZN => n22971);
   U20498 : AOI22_X1 port map( A1 => n25158, A2 => n20079, B1 => n25152, B2 => 
                           n17359, ZN => n22972);
   U20499 : OAI221_X1 port map( B1 => n19758, B2 => n25170, C1 => n19822, C2 =>
                           n25164, A => n22954, ZN => n22953);
   U20500 : AOI22_X1 port map( A1 => n25158, A2 => n20078, B1 => n25152, B2 => 
                           n17338, ZN => n22954);
   U20501 : OAI221_X1 port map( B1 => n19757, B2 => n25170, C1 => n19821, C2 =>
                           n25164, A => n22936, ZN => n22935);
   U20502 : AOI22_X1 port map( A1 => n25158, A2 => n20077, B1 => n25152, B2 => 
                           n17317, ZN => n22936);
   U20503 : OAI221_X1 port map( B1 => n19756, B2 => n25170, C1 => n19820, C2 =>
                           n25164, A => n22918, ZN => n22917);
   U20504 : AOI22_X1 port map( A1 => n25158, A2 => n20076, B1 => n25152, B2 => 
                           n17296, ZN => n22918);
   U20505 : OAI221_X1 port map( B1 => n19755, B2 => n25170, C1 => n19819, C2 =>
                           n25164, A => n22900, ZN => n22899);
   U20506 : AOI22_X1 port map( A1 => n25158, A2 => n20075, B1 => n25152, B2 => 
                           n17275, ZN => n22900);
   U20507 : OAI221_X1 port map( B1 => n19754, B2 => n25170, C1 => n19818, C2 =>
                           n25164, A => n22882, ZN => n22881);
   U20508 : AOI22_X1 port map( A1 => n25158, A2 => n20074, B1 => n25152, B2 => 
                           n17254, ZN => n22882);
   U20509 : OAI221_X1 port map( B1 => n19753, B2 => n25170, C1 => n19817, C2 =>
                           n25164, A => n22864, ZN => n22863);
   U20510 : AOI22_X1 port map( A1 => n25158, A2 => n20073, B1 => n25152, B2 => 
                           n17233, ZN => n22864);
   U20511 : OAI221_X1 port map( B1 => n19800, B2 => n25365, C1 => n19864, C2 =>
                           n25359, A => n22513, ZN => n22512);
   U20512 : AOI22_X1 port map( A1 => n25353, A2 => n20120, B1 => n25347, B2 => 
                           n18220, ZN => n22513);
   U20513 : OAI221_X1 port map( B1 => n19799, B2 => n25365, C1 => n19863, C2 =>
                           n25359, A => n22495, ZN => n22494);
   U20514 : AOI22_X1 port map( A1 => n25353, A2 => n20119, B1 => n25347, B2 => 
                           n18199, ZN => n22495);
   U20515 : OAI221_X1 port map( B1 => n19798, B2 => n25365, C1 => n19862, C2 =>
                           n25359, A => n22477, ZN => n22476);
   U20516 : AOI22_X1 port map( A1 => n25353, A2 => n20118, B1 => n25347, B2 => 
                           n18178, ZN => n22477);
   U20517 : OAI221_X1 port map( B1 => n19797, B2 => n25365, C1 => n19861, C2 =>
                           n25359, A => n22459, ZN => n22458);
   U20518 : AOI22_X1 port map( A1 => n25353, A2 => n20117, B1 => n25347, B2 => 
                           n18157, ZN => n22459);
   U20519 : OAI221_X1 port map( B1 => n19796, B2 => n25365, C1 => n19860, C2 =>
                           n25359, A => n22441, ZN => n22440);
   U20520 : AOI22_X1 port map( A1 => n25353, A2 => n20116, B1 => n25347, B2 => 
                           n18136, ZN => n22441);
   U20521 : OAI221_X1 port map( B1 => n19795, B2 => n25365, C1 => n19859, C2 =>
                           n25359, A => n22423, ZN => n22422);
   U20522 : AOI22_X1 port map( A1 => n25353, A2 => n20115, B1 => n25347, B2 => 
                           n18115, ZN => n22423);
   U20523 : OAI221_X1 port map( B1 => n19794, B2 => n25365, C1 => n19858, C2 =>
                           n25359, A => n22405, ZN => n22404);
   U20524 : AOI22_X1 port map( A1 => n25353, A2 => n20114, B1 => n25347, B2 => 
                           n18094, ZN => n22405);
   U20525 : OAI221_X1 port map( B1 => n19793, B2 => n25365, C1 => n19857, C2 =>
                           n25359, A => n22387, ZN => n22386);
   U20526 : AOI22_X1 port map( A1 => n25353, A2 => n20113, B1 => n25347, B2 => 
                           n18073, ZN => n22387);
   U20527 : OAI221_X1 port map( B1 => n19792, B2 => n25365, C1 => n19856, C2 =>
                           n25359, A => n22369, ZN => n22368);
   U20528 : AOI22_X1 port map( A1 => n25353, A2 => n20112, B1 => n25347, B2 => 
                           n18052, ZN => n22369);
   U20529 : OAI221_X1 port map( B1 => n19791, B2 => n25365, C1 => n19855, C2 =>
                           n25359, A => n22351, ZN => n22350);
   U20530 : AOI22_X1 port map( A1 => n25353, A2 => n20111, B1 => n25347, B2 => 
                           n18031, ZN => n22351);
   U20531 : OAI221_X1 port map( B1 => n19790, B2 => n25365, C1 => n19854, C2 =>
                           n25359, A => n22333, ZN => n22332);
   U20532 : AOI22_X1 port map( A1 => n25353, A2 => n20110, B1 => n25347, B2 => 
                           n18010, ZN => n22333);
   U20533 : OAI221_X1 port map( B1 => n19789, B2 => n25365, C1 => n19853, C2 =>
                           n25359, A => n22315, ZN => n22314);
   U20534 : AOI22_X1 port map( A1 => n25353, A2 => n20109, B1 => n25347, B2 => 
                           n17989, ZN => n22315);
   U20535 : OAI221_X1 port map( B1 => n19788, B2 => n25366, C1 => n19852, C2 =>
                           n25360, A => n22297, ZN => n22296);
   U20536 : AOI22_X1 port map( A1 => n25354, A2 => n20108, B1 => n25348, B2 => 
                           n17968, ZN => n22297);
   U20537 : OAI221_X1 port map( B1 => n19787, B2 => n25366, C1 => n19851, C2 =>
                           n25360, A => n22279, ZN => n22278);
   U20538 : AOI22_X1 port map( A1 => n25354, A2 => n20107, B1 => n25348, B2 => 
                           n17947, ZN => n22279);
   U20539 : OAI221_X1 port map( B1 => n19786, B2 => n25366, C1 => n19850, C2 =>
                           n25360, A => n22261, ZN => n22260);
   U20540 : AOI22_X1 port map( A1 => n25354, A2 => n20106, B1 => n25348, B2 => 
                           n17926, ZN => n22261);
   U20541 : OAI221_X1 port map( B1 => n19785, B2 => n25366, C1 => n19849, C2 =>
                           n25360, A => n22243, ZN => n22242);
   U20542 : AOI22_X1 port map( A1 => n25354, A2 => n20105, B1 => n25348, B2 => 
                           n17905, ZN => n22243);
   U20543 : OAI221_X1 port map( B1 => n19784, B2 => n25366, C1 => n19848, C2 =>
                           n25360, A => n22225, ZN => n22224);
   U20544 : AOI22_X1 port map( A1 => n25354, A2 => n20104, B1 => n25348, B2 => 
                           n17884, ZN => n22225);
   U20545 : OAI221_X1 port map( B1 => n19783, B2 => n25366, C1 => n19847, C2 =>
                           n25360, A => n22207, ZN => n22206);
   U20546 : AOI22_X1 port map( A1 => n25354, A2 => n20103, B1 => n25348, B2 => 
                           n17863, ZN => n22207);
   U20547 : OAI221_X1 port map( B1 => n19782, B2 => n25366, C1 => n19846, C2 =>
                           n25360, A => n22189, ZN => n22188);
   U20548 : AOI22_X1 port map( A1 => n25354, A2 => n20102, B1 => n25348, B2 => 
                           n17842, ZN => n22189);
   U20549 : OAI221_X1 port map( B1 => n19781, B2 => n25366, C1 => n19845, C2 =>
                           n25360, A => n22171, ZN => n22170);
   U20550 : AOI22_X1 port map( A1 => n25354, A2 => n20101, B1 => n25348, B2 => 
                           n17821, ZN => n22171);
   U20551 : OAI221_X1 port map( B1 => n19780, B2 => n25366, C1 => n19844, C2 =>
                           n25360, A => n22153, ZN => n22152);
   U20552 : AOI22_X1 port map( A1 => n25354, A2 => n20100, B1 => n25348, B2 => 
                           n17800, ZN => n22153);
   U20553 : OAI221_X1 port map( B1 => n19779, B2 => n25366, C1 => n19843, C2 =>
                           n25360, A => n22135, ZN => n22134);
   U20554 : AOI22_X1 port map( A1 => n25354, A2 => n20099, B1 => n25348, B2 => 
                           n17779, ZN => n22135);
   U20555 : OAI221_X1 port map( B1 => n19778, B2 => n25366, C1 => n19842, C2 =>
                           n25360, A => n22117, ZN => n22116);
   U20556 : AOI22_X1 port map( A1 => n25354, A2 => n20098, B1 => n25348, B2 => 
                           n17758, ZN => n22117);
   U20557 : OAI221_X1 port map( B1 => n19777, B2 => n25366, C1 => n19841, C2 =>
                           n25360, A => n22099, ZN => n22098);
   U20558 : AOI22_X1 port map( A1 => n25354, A2 => n20097, B1 => n25348, B2 => 
                           n17737, ZN => n22099);
   U20559 : OAI221_X1 port map( B1 => n19776, B2 => n25367, C1 => n19840, C2 =>
                           n25361, A => n22081, ZN => n22080);
   U20560 : AOI22_X1 port map( A1 => n25355, A2 => n20096, B1 => n25349, B2 => 
                           n17716, ZN => n22081);
   U20561 : OAI221_X1 port map( B1 => n19775, B2 => n25367, C1 => n19839, C2 =>
                           n25361, A => n22063, ZN => n22062);
   U20562 : AOI22_X1 port map( A1 => n25355, A2 => n20095, B1 => n25349, B2 => 
                           n17695, ZN => n22063);
   U20563 : OAI221_X1 port map( B1 => n19774, B2 => n25367, C1 => n19838, C2 =>
                           n25361, A => n22045, ZN => n22044);
   U20564 : AOI22_X1 port map( A1 => n25355, A2 => n20094, B1 => n25349, B2 => 
                           n17674, ZN => n22045);
   U20565 : OAI221_X1 port map( B1 => n19773, B2 => n25367, C1 => n19837, C2 =>
                           n25361, A => n22027, ZN => n22026);
   U20566 : AOI22_X1 port map( A1 => n25355, A2 => n20093, B1 => n25349, B2 => 
                           n17653, ZN => n22027);
   U20567 : OAI221_X1 port map( B1 => n19772, B2 => n25367, C1 => n19836, C2 =>
                           n25361, A => n22009, ZN => n22008);
   U20568 : AOI22_X1 port map( A1 => n25355, A2 => n20092, B1 => n25349, B2 => 
                           n17632, ZN => n22009);
   U20569 : OAI221_X1 port map( B1 => n19771, B2 => n25367, C1 => n19835, C2 =>
                           n25361, A => n21991, ZN => n21990);
   U20570 : AOI22_X1 port map( A1 => n25355, A2 => n20091, B1 => n25349, B2 => 
                           n17611, ZN => n21991);
   U20571 : OAI221_X1 port map( B1 => n19770, B2 => n25367, C1 => n19834, C2 =>
                           n25361, A => n21973, ZN => n21972);
   U20572 : AOI22_X1 port map( A1 => n25355, A2 => n20090, B1 => n25349, B2 => 
                           n17590, ZN => n21973);
   U20573 : OAI221_X1 port map( B1 => n19769, B2 => n25367, C1 => n19833, C2 =>
                           n25361, A => n21955, ZN => n21954);
   U20574 : AOI22_X1 port map( A1 => n25355, A2 => n20089, B1 => n25349, B2 => 
                           n17569, ZN => n21955);
   U20575 : OAI221_X1 port map( B1 => n19768, B2 => n25367, C1 => n19832, C2 =>
                           n25361, A => n21937, ZN => n21936);
   U20576 : AOI22_X1 port map( A1 => n25355, A2 => n20088, B1 => n25349, B2 => 
                           n17548, ZN => n21937);
   U20577 : OAI221_X1 port map( B1 => n19767, B2 => n25367, C1 => n19831, C2 =>
                           n25361, A => n21919, ZN => n21918);
   U20578 : AOI22_X1 port map( A1 => n25355, A2 => n20087, B1 => n25349, B2 => 
                           n17527, ZN => n21919);
   U20579 : OAI221_X1 port map( B1 => n19766, B2 => n25367, C1 => n19830, C2 =>
                           n25361, A => n21901, ZN => n21900);
   U20580 : AOI22_X1 port map( A1 => n25355, A2 => n20086, B1 => n25349, B2 => 
                           n17506, ZN => n21901);
   U20581 : OAI221_X1 port map( B1 => n19765, B2 => n25367, C1 => n19829, C2 =>
                           n25361, A => n21883, ZN => n21882);
   U20582 : AOI22_X1 port map( A1 => n25355, A2 => n20085, B1 => n25349, B2 => 
                           n17485, ZN => n21883);
   U20583 : OAI221_X1 port map( B1 => n19764, B2 => n25368, C1 => n19828, C2 =>
                           n25362, A => n21865, ZN => n21864);
   U20584 : AOI22_X1 port map( A1 => n25356, A2 => n20084, B1 => n25350, B2 => 
                           n17464, ZN => n21865);
   U20585 : OAI221_X1 port map( B1 => n19763, B2 => n25368, C1 => n19827, C2 =>
                           n25362, A => n21847, ZN => n21846);
   U20586 : AOI22_X1 port map( A1 => n25356, A2 => n20083, B1 => n25350, B2 => 
                           n17443, ZN => n21847);
   U20587 : OAI221_X1 port map( B1 => n19762, B2 => n25368, C1 => n19826, C2 =>
                           n25362, A => n21829, ZN => n21828);
   U20588 : AOI22_X1 port map( A1 => n25356, A2 => n20082, B1 => n25350, B2 => 
                           n17422, ZN => n21829);
   U20589 : OAI221_X1 port map( B1 => n19761, B2 => n25368, C1 => n19825, C2 =>
                           n25362, A => n21811, ZN => n21810);
   U20590 : AOI22_X1 port map( A1 => n25356, A2 => n20081, B1 => n25350, B2 => 
                           n17401, ZN => n21811);
   U20591 : OAI221_X1 port map( B1 => n19760, B2 => n25368, C1 => n19824, C2 =>
                           n25362, A => n21793, ZN => n21792);
   U20592 : AOI22_X1 port map( A1 => n25356, A2 => n20080, B1 => n25350, B2 => 
                           n17380, ZN => n21793);
   U20593 : OAI221_X1 port map( B1 => n19759, B2 => n25368, C1 => n19823, C2 =>
                           n25362, A => n21775, ZN => n21774);
   U20594 : AOI22_X1 port map( A1 => n25356, A2 => n20079, B1 => n25350, B2 => 
                           n17359, ZN => n21775);
   U20595 : OAI221_X1 port map( B1 => n19758, B2 => n25368, C1 => n19822, C2 =>
                           n25362, A => n21757, ZN => n21756);
   U20596 : AOI22_X1 port map( A1 => n25356, A2 => n20078, B1 => n25350, B2 => 
                           n17338, ZN => n21757);
   U20597 : OAI221_X1 port map( B1 => n19757, B2 => n25368, C1 => n19821, C2 =>
                           n25362, A => n21739, ZN => n21738);
   U20598 : AOI22_X1 port map( A1 => n25356, A2 => n20077, B1 => n25350, B2 => 
                           n17317, ZN => n21739);
   U20599 : OAI221_X1 port map( B1 => n19756, B2 => n25368, C1 => n19820, C2 =>
                           n25362, A => n21721, ZN => n21720);
   U20600 : AOI22_X1 port map( A1 => n25356, A2 => n20076, B1 => n25350, B2 => 
                           n17296, ZN => n21721);
   U20601 : OAI221_X1 port map( B1 => n19755, B2 => n25368, C1 => n19819, C2 =>
                           n25362, A => n21703, ZN => n21702);
   U20602 : AOI22_X1 port map( A1 => n25356, A2 => n20075, B1 => n25350, B2 => 
                           n17275, ZN => n21703);
   U20603 : OAI221_X1 port map( B1 => n19754, B2 => n25368, C1 => n19818, C2 =>
                           n25362, A => n21685, ZN => n21684);
   U20604 : AOI22_X1 port map( A1 => n25356, A2 => n20074, B1 => n25350, B2 => 
                           n17254, ZN => n21685);
   U20605 : OAI221_X1 port map( B1 => n19753, B2 => n25368, C1 => n19817, C2 =>
                           n25362, A => n21667, ZN => n21666);
   U20606 : AOI22_X1 port map( A1 => n25356, A2 => n20073, B1 => n25350, B2 => 
                           n17233, ZN => n21667);
   U20607 : OAI221_X1 port map( B1 => n20133, B2 => n25171, C1 => n19813, C2 =>
                           n25165, A => n22761, ZN => n22758);
   U20608 : AOI22_X1 port map( A1 => n25159, A2 => n20069, B1 => n25153, B2 => 
                           n17149, ZN => n22761);
   U20609 : OAI221_X1 port map( B1 => n21098, B2 => n25069, C1 => n20134, C2 =>
                           n25063, A => n22786, ZN => n22783);
   U20610 : AOI22_X1 port map( A1 => n25057, A2 => n24085, B1 => n25048, B2 => 
                           OUT2_63_port, ZN => n22786);
   U20611 : OAI221_X1 port map( B1 => n19752, B2 => n25171, C1 => n19816, C2 =>
                           n25165, A => n22846, ZN => n22845);
   U20612 : AOI22_X1 port map( A1 => n25159, A2 => n20072, B1 => n25153, B2 => 
                           n17212, ZN => n22846);
   U20613 : OAI221_X1 port map( B1 => n21101, B2 => n25069, C1 => n20137, C2 =>
                           n25063, A => n22854, ZN => n22853);
   U20614 : AOI22_X1 port map( A1 => n25057, A2 => n24079, B1 => n25046, B2 => 
                           OUT2_60_port, ZN => n22854);
   U20615 : OAI221_X1 port map( B1 => n19751, B2 => n25171, C1 => n19815, C2 =>
                           n25165, A => n22828, ZN => n22827);
   U20616 : AOI22_X1 port map( A1 => n25159, A2 => n20071, B1 => n25153, B2 => 
                           n17191, ZN => n22828);
   U20617 : OAI221_X1 port map( B1 => n21100, B2 => n25069, C1 => n20136, C2 =>
                           n25063, A => n22836, ZN => n22835);
   U20618 : AOI22_X1 port map( A1 => n25057, A2 => n24081, B1 => n25046, B2 => 
                           OUT2_61_port, ZN => n22836);
   U20619 : OAI221_X1 port map( B1 => n19750, B2 => n25171, C1 => n19814, C2 =>
                           n25165, A => n22810, ZN => n22809);
   U20620 : AOI22_X1 port map( A1 => n25159, A2 => n20070, B1 => n25153, B2 => 
                           n17170, ZN => n22810);
   U20621 : OAI221_X1 port map( B1 => n21099, B2 => n25069, C1 => n20135, C2 =>
                           n25063, A => n22818, ZN => n22817);
   U20622 : AOI22_X1 port map( A1 => n25057, A2 => n24083, B1 => n25046, B2 => 
                           OUT2_62_port, ZN => n22818);
   U20623 : OAI221_X1 port map( B1 => n19752, B2 => n25369, C1 => n19816, C2 =>
                           n25363, A => n21649, ZN => n21648);
   U20624 : AOI22_X1 port map( A1 => n25357, A2 => n20072, B1 => n25351, B2 => 
                           n17212, ZN => n21649);
   U20625 : OAI221_X1 port map( B1 => n21101, B2 => n25267, C1 => n20137, C2 =>
                           n25261, A => n21657, ZN => n21656);
   U20626 : AOI22_X1 port map( A1 => n25255, A2 => n24079, B1 => n25244, B2 => 
                           OUT1_60_port, ZN => n21657);
   U20627 : OAI221_X1 port map( B1 => n19751, B2 => n25369, C1 => n19815, C2 =>
                           n25363, A => n21631, ZN => n21630);
   U20628 : AOI22_X1 port map( A1 => n25357, A2 => n20071, B1 => n25351, B2 => 
                           n17191, ZN => n21631);
   U20629 : OAI221_X1 port map( B1 => n21100, B2 => n25267, C1 => n20136, C2 =>
                           n25261, A => n21639, ZN => n21638);
   U20630 : AOI22_X1 port map( A1 => n25255, A2 => n24081, B1 => n25244, B2 => 
                           OUT1_61_port, ZN => n21639);
   U20631 : OAI221_X1 port map( B1 => n19750, B2 => n25369, C1 => n19814, C2 =>
                           n25363, A => n21613, ZN => n21612);
   U20632 : AOI22_X1 port map( A1 => n25357, A2 => n20070, B1 => n25351, B2 => 
                           n17170, ZN => n21613);
   U20633 : OAI221_X1 port map( B1 => n21099, B2 => n25267, C1 => n20135, C2 =>
                           n25261, A => n21621, ZN => n21620);
   U20634 : AOI22_X1 port map( A1 => n25255, A2 => n24083, B1 => n25244, B2 => 
                           OUT1_62_port, ZN => n21621);
   U20635 : OAI221_X1 port map( B1 => n20133, B2 => n25369, C1 => n19813, C2 =>
                           n25363, A => n21564, ZN => n21561);
   U20636 : AOI22_X1 port map( A1 => n25357, A2 => n20069, B1 => n25351, B2 => 
                           n17149, ZN => n21564);
   U20637 : OAI221_X1 port map( B1 => n21098, B2 => n25267, C1 => n20134, C2 =>
                           n25261, A => n21589, ZN => n21586);
   U20638 : AOI22_X1 port map( A1 => n25255, A2 => n24085, B1 => n25246, B2 => 
                           OUT1_63_port, ZN => n21589);
   U20639 : OAI221_X1 port map( B1 => n19812, B2 => n25166, C1 => n19876, C2 =>
                           n25160, A => n23926, ZN => n23925);
   U20640 : AOI22_X1 port map( A1 => n25154, A2 => n20132, B1 => n25148, B2 => 
                           n18472, ZN => n23926);
   U20641 : OAI221_X1 port map( B1 => n19811, B2 => n25166, C1 => n19875, C2 =>
                           n25160, A => n23908, ZN => n23907);
   U20642 : AOI22_X1 port map( A1 => n25154, A2 => n20131, B1 => n25148, B2 => 
                           n18451, ZN => n23908);
   U20643 : OAI221_X1 port map( B1 => n19810, B2 => n25166, C1 => n19874, C2 =>
                           n25160, A => n23890, ZN => n23889);
   U20644 : AOI22_X1 port map( A1 => n25154, A2 => n20130, B1 => n25148, B2 => 
                           n18430, ZN => n23890);
   U20645 : OAI221_X1 port map( B1 => n19809, B2 => n25166, C1 => n19873, C2 =>
                           n25160, A => n23872, ZN => n23871);
   U20646 : AOI22_X1 port map( A1 => n25154, A2 => n20129, B1 => n25148, B2 => 
                           n18409, ZN => n23872);
   U20647 : OAI221_X1 port map( B1 => n19808, B2 => n25166, C1 => n19872, C2 =>
                           n25160, A => n23854, ZN => n23853);
   U20648 : AOI22_X1 port map( A1 => n25154, A2 => n20128, B1 => n25148, B2 => 
                           n18388, ZN => n23854);
   U20649 : OAI221_X1 port map( B1 => n19807, B2 => n25166, C1 => n19871, C2 =>
                           n25160, A => n23836, ZN => n23835);
   U20650 : AOI22_X1 port map( A1 => n25154, A2 => n20127, B1 => n25148, B2 => 
                           n18367, ZN => n23836);
   U20651 : OAI221_X1 port map( B1 => n19806, B2 => n25166, C1 => n19870, C2 =>
                           n25160, A => n23818, ZN => n23817);
   U20652 : AOI22_X1 port map( A1 => n25154, A2 => n20126, B1 => n25148, B2 => 
                           n18346, ZN => n23818);
   U20653 : OAI221_X1 port map( B1 => n19805, B2 => n25166, C1 => n19869, C2 =>
                           n25160, A => n23800, ZN => n23799);
   U20654 : AOI22_X1 port map( A1 => n25154, A2 => n20125, B1 => n25148, B2 => 
                           n18325, ZN => n23800);
   U20655 : OAI221_X1 port map( B1 => n19804, B2 => n25166, C1 => n19868, C2 =>
                           n25160, A => n23782, ZN => n23781);
   U20656 : AOI22_X1 port map( A1 => n25154, A2 => n20124, B1 => n25148, B2 => 
                           n18304, ZN => n23782);
   U20657 : OAI221_X1 port map( B1 => n19803, B2 => n25166, C1 => n19867, C2 =>
                           n25160, A => n23764, ZN => n23763);
   U20658 : AOI22_X1 port map( A1 => n25154, A2 => n20123, B1 => n25148, B2 => 
                           n18283, ZN => n23764);
   U20659 : OAI221_X1 port map( B1 => n19802, B2 => n25166, C1 => n19866, C2 =>
                           n25160, A => n23746, ZN => n23745);
   U20660 : AOI22_X1 port map( A1 => n25154, A2 => n20122, B1 => n25148, B2 => 
                           n18262, ZN => n23746);
   U20661 : OAI221_X1 port map( B1 => n19801, B2 => n25166, C1 => n19865, C2 =>
                           n25160, A => n23728, ZN => n23727);
   U20662 : AOI22_X1 port map( A1 => n25154, A2 => n20121, B1 => n25148, B2 => 
                           n18241, ZN => n23728);
   U20663 : OAI221_X1 port map( B1 => n19812, B2 => n25364, C1 => n19876, C2 =>
                           n25358, A => n22729, ZN => n22728);
   U20664 : AOI22_X1 port map( A1 => n25352, A2 => n20132, B1 => n25346, B2 => 
                           n18472, ZN => n22729);
   U20665 : OAI221_X1 port map( B1 => n19811, B2 => n25364, C1 => n19875, C2 =>
                           n25358, A => n22711, ZN => n22710);
   U20666 : AOI22_X1 port map( A1 => n25352, A2 => n20131, B1 => n25346, B2 => 
                           n18451, ZN => n22711);
   U20667 : OAI221_X1 port map( B1 => n19810, B2 => n25364, C1 => n19874, C2 =>
                           n25358, A => n22693, ZN => n22692);
   U20668 : AOI22_X1 port map( A1 => n25352, A2 => n20130, B1 => n25346, B2 => 
                           n18430, ZN => n22693);
   U20669 : OAI221_X1 port map( B1 => n19809, B2 => n25364, C1 => n19873, C2 =>
                           n25358, A => n22675, ZN => n22674);
   U20670 : AOI22_X1 port map( A1 => n25352, A2 => n20129, B1 => n25346, B2 => 
                           n18409, ZN => n22675);
   U20671 : OAI221_X1 port map( B1 => n19808, B2 => n25364, C1 => n19872, C2 =>
                           n25358, A => n22657, ZN => n22656);
   U20672 : AOI22_X1 port map( A1 => n25352, A2 => n20128, B1 => n25346, B2 => 
                           n18388, ZN => n22657);
   U20673 : OAI221_X1 port map( B1 => n19807, B2 => n25364, C1 => n19871, C2 =>
                           n25358, A => n22639, ZN => n22638);
   U20674 : AOI22_X1 port map( A1 => n25352, A2 => n20127, B1 => n25346, B2 => 
                           n18367, ZN => n22639);
   U20675 : OAI221_X1 port map( B1 => n19806, B2 => n25364, C1 => n19870, C2 =>
                           n25358, A => n22621, ZN => n22620);
   U20676 : AOI22_X1 port map( A1 => n25352, A2 => n20126, B1 => n25346, B2 => 
                           n18346, ZN => n22621);
   U20677 : OAI221_X1 port map( B1 => n19805, B2 => n25364, C1 => n19869, C2 =>
                           n25358, A => n22603, ZN => n22602);
   U20678 : AOI22_X1 port map( A1 => n25352, A2 => n20125, B1 => n25346, B2 => 
                           n18325, ZN => n22603);
   U20679 : OAI221_X1 port map( B1 => n19804, B2 => n25364, C1 => n19868, C2 =>
                           n25358, A => n22585, ZN => n22584);
   U20680 : AOI22_X1 port map( A1 => n25352, A2 => n20124, B1 => n25346, B2 => 
                           n18304, ZN => n22585);
   U20681 : OAI221_X1 port map( B1 => n19803, B2 => n25364, C1 => n19867, C2 =>
                           n25358, A => n22567, ZN => n22566);
   U20682 : AOI22_X1 port map( A1 => n25352, A2 => n20123, B1 => n25346, B2 => 
                           n18283, ZN => n22567);
   U20683 : OAI221_X1 port map( B1 => n19802, B2 => n25364, C1 => n19866, C2 =>
                           n25358, A => n22549, ZN => n22548);
   U20684 : AOI22_X1 port map( A1 => n25352, A2 => n20122, B1 => n25346, B2 => 
                           n18262, ZN => n22549);
   U20685 : OAI221_X1 port map( B1 => n19801, B2 => n25364, C1 => n19865, C2 =>
                           n25358, A => n22531, ZN => n22530);
   U20686 : AOI22_X1 port map( A1 => n25352, A2 => n20121, B1 => n25346, B2 => 
                           n18241, ZN => n22531);
   U20687 : OAI221_X1 port map( B1 => n9466, B2 => n25143, C1 => n20449, C2 => 
                           n25137, A => n23711, ZN => n23708);
   U20688 : AOI22_X1 port map( A1 => n25131, A2 => n24030, B1 => n25125, B2 => 
                           n18219, ZN => n23711);
   U20689 : OAI221_X1 port map( B1 => n21149, B2 => n25041, C1 => n20385, C2 =>
                           n25035, A => n23719, ZN => n23716);
   U20690 : AOI22_X1 port map( A1 => n25029, A2 => n24339, B1 => n25023, B2 => 
                           n18232, ZN => n23719);
   U20691 : OAI221_X1 port map( B1 => n9465, B2 => n25143, C1 => n20448, C2 => 
                           n25137, A => n23693, ZN => n23690);
   U20692 : AOI22_X1 port map( A1 => n25131, A2 => n24031, B1 => n25125, B2 => 
                           n18198, ZN => n23693);
   U20693 : OAI221_X1 port map( B1 => n21148, B2 => n25041, C1 => n20384, C2 =>
                           n25035, A => n23701, ZN => n23698);
   U20694 : AOI22_X1 port map( A1 => n25029, A2 => n24341, B1 => n25023, B2 => 
                           n18211, ZN => n23701);
   U20695 : OAI221_X1 port map( B1 => n9464, B2 => n25143, C1 => n20447, C2 => 
                           n25137, A => n23675, ZN => n23672);
   U20696 : AOI22_X1 port map( A1 => n25131, A2 => n24032, B1 => n25125, B2 => 
                           n18177, ZN => n23675);
   U20697 : OAI221_X1 port map( B1 => n21147, B2 => n25041, C1 => n20383, C2 =>
                           n25035, A => n23683, ZN => n23680);
   U20698 : AOI22_X1 port map( A1 => n25029, A2 => n24343, B1 => n25023, B2 => 
                           n18190, ZN => n23683);
   U20699 : OAI221_X1 port map( B1 => n9463, B2 => n25143, C1 => n20446, C2 => 
                           n25137, A => n23657, ZN => n23654);
   U20700 : AOI22_X1 port map( A1 => n25131, A2 => n24033, B1 => n25125, B2 => 
                           n18156, ZN => n23657);
   U20701 : OAI221_X1 port map( B1 => n21146, B2 => n25041, C1 => n20382, C2 =>
                           n25035, A => n23665, ZN => n23662);
   U20702 : AOI22_X1 port map( A1 => n25029, A2 => n24345, B1 => n25023, B2 => 
                           n18169, ZN => n23665);
   U20703 : OAI221_X1 port map( B1 => n9462, B2 => n25143, C1 => n20445, C2 => 
                           n25137, A => n23639, ZN => n23636);
   U20704 : AOI22_X1 port map( A1 => n25131, A2 => n24034, B1 => n25125, B2 => 
                           n18135, ZN => n23639);
   U20705 : OAI221_X1 port map( B1 => n21145, B2 => n25041, C1 => n20381, C2 =>
                           n25035, A => n23647, ZN => n23644);
   U20706 : AOI22_X1 port map( A1 => n25029, A2 => n24347, B1 => n25023, B2 => 
                           n18148, ZN => n23647);
   U20707 : OAI221_X1 port map( B1 => n9461, B2 => n25143, C1 => n20444, C2 => 
                           n25137, A => n23621, ZN => n23618);
   U20708 : AOI22_X1 port map( A1 => n25131, A2 => n24035, B1 => n25125, B2 => 
                           n18114, ZN => n23621);
   U20709 : OAI221_X1 port map( B1 => n21144, B2 => n25041, C1 => n20380, C2 =>
                           n25035, A => n23629, ZN => n23626);
   U20710 : AOI22_X1 port map( A1 => n25029, A2 => n24349, B1 => n25023, B2 => 
                           n18127, ZN => n23629);
   U20711 : OAI221_X1 port map( B1 => n9460, B2 => n25143, C1 => n20443, C2 => 
                           n25137, A => n23603, ZN => n23600);
   U20712 : AOI22_X1 port map( A1 => n25131, A2 => n24036, B1 => n25125, B2 => 
                           n18093, ZN => n23603);
   U20713 : OAI221_X1 port map( B1 => n21143, B2 => n25041, C1 => n20379, C2 =>
                           n25035, A => n23611, ZN => n23608);
   U20714 : AOI22_X1 port map( A1 => n25029, A2 => n24351, B1 => n25023, B2 => 
                           n18106, ZN => n23611);
   U20715 : OAI221_X1 port map( B1 => n9459, B2 => n25143, C1 => n20442, C2 => 
                           n25137, A => n23585, ZN => n23582);
   U20716 : AOI22_X1 port map( A1 => n25131, A2 => n24037, B1 => n25125, B2 => 
                           n18072, ZN => n23585);
   U20717 : OAI221_X1 port map( B1 => n21142, B2 => n25041, C1 => n20378, C2 =>
                           n25035, A => n23593, ZN => n23590);
   U20718 : AOI22_X1 port map( A1 => n25029, A2 => n24353, B1 => n25023, B2 => 
                           n18085, ZN => n23593);
   U20719 : OAI221_X1 port map( B1 => n9458, B2 => n25143, C1 => n20441, C2 => 
                           n25137, A => n23567, ZN => n23564);
   U20720 : AOI22_X1 port map( A1 => n25131, A2 => n24038, B1 => n25125, B2 => 
                           n18051, ZN => n23567);
   U20721 : OAI221_X1 port map( B1 => n21141, B2 => n25041, C1 => n20377, C2 =>
                           n25035, A => n23575, ZN => n23572);
   U20722 : AOI22_X1 port map( A1 => n25029, A2 => n24355, B1 => n25023, B2 => 
                           n18064, ZN => n23575);
   U20723 : OAI221_X1 port map( B1 => n9457, B2 => n25143, C1 => n20440, C2 => 
                           n25137, A => n23549, ZN => n23546);
   U20724 : AOI22_X1 port map( A1 => n25131, A2 => n24039, B1 => n25125, B2 => 
                           n18030, ZN => n23549);
   U20725 : OAI221_X1 port map( B1 => n21140, B2 => n25041, C1 => n20376, C2 =>
                           n25035, A => n23557, ZN => n23554);
   U20726 : AOI22_X1 port map( A1 => n25029, A2 => n24357, B1 => n25023, B2 => 
                           n18043, ZN => n23557);
   U20727 : OAI221_X1 port map( B1 => n9456, B2 => n25143, C1 => n20439, C2 => 
                           n25137, A => n23531, ZN => n23528);
   U20728 : AOI22_X1 port map( A1 => n25131, A2 => n24040, B1 => n25125, B2 => 
                           n18009, ZN => n23531);
   U20729 : OAI221_X1 port map( B1 => n21139, B2 => n25041, C1 => n20375, C2 =>
                           n25035, A => n23539, ZN => n23536);
   U20730 : AOI22_X1 port map( A1 => n25029, A2 => n24359, B1 => n25023, B2 => 
                           n18022, ZN => n23539);
   U20731 : OAI221_X1 port map( B1 => n9455, B2 => n25143, C1 => n20438, C2 => 
                           n25137, A => n23513, ZN => n23510);
   U20732 : AOI22_X1 port map( A1 => n25131, A2 => n24041, B1 => n25125, B2 => 
                           n17988, ZN => n23513);
   U20733 : OAI221_X1 port map( B1 => n21138, B2 => n25041, C1 => n20374, C2 =>
                           n25035, A => n23521, ZN => n23518);
   U20734 : AOI22_X1 port map( A1 => n25029, A2 => n24361, B1 => n25023, B2 => 
                           n18001, ZN => n23521);
   U20735 : OAI221_X1 port map( B1 => n9454, B2 => n25144, C1 => n20437, C2 => 
                           n25138, A => n23495, ZN => n23492);
   U20736 : AOI22_X1 port map( A1 => n25132, A2 => n24042, B1 => n25126, B2 => 
                           n17967, ZN => n23495);
   U20737 : OAI221_X1 port map( B1 => n21137, B2 => n25042, C1 => n20373, C2 =>
                           n25036, A => n23503, ZN => n23500);
   U20738 : AOI22_X1 port map( A1 => n25030, A2 => n24363, B1 => n25024, B2 => 
                           n17980, ZN => n23503);
   U20739 : OAI221_X1 port map( B1 => n9453, B2 => n25144, C1 => n20436, C2 => 
                           n25138, A => n23477, ZN => n23474);
   U20740 : AOI22_X1 port map( A1 => n25132, A2 => n24043, B1 => n25126, B2 => 
                           n17946, ZN => n23477);
   U20741 : OAI221_X1 port map( B1 => n21136, B2 => n25042, C1 => n20372, C2 =>
                           n25036, A => n23485, ZN => n23482);
   U20742 : AOI22_X1 port map( A1 => n25030, A2 => n24365, B1 => n25024, B2 => 
                           n17959, ZN => n23485);
   U20743 : OAI221_X1 port map( B1 => n9452, B2 => n25144, C1 => n20435, C2 => 
                           n25138, A => n23459, ZN => n23456);
   U20744 : AOI22_X1 port map( A1 => n25132, A2 => n24044, B1 => n25126, B2 => 
                           n17925, ZN => n23459);
   U20745 : OAI221_X1 port map( B1 => n21135, B2 => n25042, C1 => n20371, C2 =>
                           n25036, A => n23467, ZN => n23464);
   U20746 : AOI22_X1 port map( A1 => n25030, A2 => n24367, B1 => n25024, B2 => 
                           n17938, ZN => n23467);
   U20747 : OAI221_X1 port map( B1 => n9451, B2 => n25144, C1 => n20434, C2 => 
                           n25138, A => n23441, ZN => n23438);
   U20748 : AOI22_X1 port map( A1 => n25132, A2 => n24045, B1 => n25126, B2 => 
                           n17904, ZN => n23441);
   U20749 : OAI221_X1 port map( B1 => n21134, B2 => n25042, C1 => n20370, C2 =>
                           n25036, A => n23449, ZN => n23446);
   U20750 : AOI22_X1 port map( A1 => n25030, A2 => n24369, B1 => n25024, B2 => 
                           n17917, ZN => n23449);
   U20751 : OAI221_X1 port map( B1 => n9450, B2 => n25144, C1 => n20433, C2 => 
                           n25138, A => n23423, ZN => n23420);
   U20752 : AOI22_X1 port map( A1 => n25132, A2 => n24046, B1 => n25126, B2 => 
                           n17883, ZN => n23423);
   U20753 : OAI221_X1 port map( B1 => n21133, B2 => n25042, C1 => n20369, C2 =>
                           n25036, A => n23431, ZN => n23428);
   U20754 : AOI22_X1 port map( A1 => n25030, A2 => n24371, B1 => n25024, B2 => 
                           n17896, ZN => n23431);
   U20755 : OAI221_X1 port map( B1 => n9449, B2 => n25144, C1 => n20432, C2 => 
                           n25138, A => n23405, ZN => n23402);
   U20756 : AOI22_X1 port map( A1 => n25132, A2 => n24047, B1 => n25126, B2 => 
                           n17862, ZN => n23405);
   U20757 : OAI221_X1 port map( B1 => n21132, B2 => n25042, C1 => n20368, C2 =>
                           n25036, A => n23413, ZN => n23410);
   U20758 : AOI22_X1 port map( A1 => n25030, A2 => n24373, B1 => n25024, B2 => 
                           n17875, ZN => n23413);
   U20759 : OAI221_X1 port map( B1 => n9448, B2 => n25144, C1 => n20431, C2 => 
                           n25138, A => n23387, ZN => n23384);
   U20760 : AOI22_X1 port map( A1 => n25132, A2 => n24048, B1 => n25126, B2 => 
                           n17841, ZN => n23387);
   U20761 : OAI221_X1 port map( B1 => n21131, B2 => n25042, C1 => n20367, C2 =>
                           n25036, A => n23395, ZN => n23392);
   U20762 : AOI22_X1 port map( A1 => n25030, A2 => n24375, B1 => n25024, B2 => 
                           n17854, ZN => n23395);
   U20763 : OAI221_X1 port map( B1 => n9447, B2 => n25144, C1 => n20430, C2 => 
                           n25138, A => n23369, ZN => n23366);
   U20764 : AOI22_X1 port map( A1 => n25132, A2 => n24049, B1 => n25126, B2 => 
                           n17820, ZN => n23369);
   U20765 : OAI221_X1 port map( B1 => n21130, B2 => n25042, C1 => n20366, C2 =>
                           n25036, A => n23377, ZN => n23374);
   U20766 : AOI22_X1 port map( A1 => n25030, A2 => n24377, B1 => n25024, B2 => 
                           n17833, ZN => n23377);
   U20767 : OAI221_X1 port map( B1 => n9446, B2 => n25144, C1 => n20429, C2 => 
                           n25138, A => n23351, ZN => n23348);
   U20768 : AOI22_X1 port map( A1 => n25132, A2 => n24050, B1 => n25126, B2 => 
                           n17799, ZN => n23351);
   U20769 : OAI221_X1 port map( B1 => n21129, B2 => n25042, C1 => n20365, C2 =>
                           n25036, A => n23359, ZN => n23356);
   U20770 : AOI22_X1 port map( A1 => n25030, A2 => n24379, B1 => n25024, B2 => 
                           n17812, ZN => n23359);
   U20771 : OAI221_X1 port map( B1 => n9445, B2 => n25144, C1 => n20428, C2 => 
                           n25138, A => n23333, ZN => n23330);
   U20772 : AOI22_X1 port map( A1 => n25132, A2 => n24051, B1 => n25126, B2 => 
                           n17778, ZN => n23333);
   U20773 : OAI221_X1 port map( B1 => n21128, B2 => n25042, C1 => n20364, C2 =>
                           n25036, A => n23341, ZN => n23338);
   U20774 : AOI22_X1 port map( A1 => n25030, A2 => n24381, B1 => n25024, B2 => 
                           n17791, ZN => n23341);
   U20775 : OAI221_X1 port map( B1 => n9444, B2 => n25144, C1 => n20427, C2 => 
                           n25138, A => n23315, ZN => n23312);
   U20776 : AOI22_X1 port map( A1 => n25132, A2 => n24052, B1 => n25126, B2 => 
                           n17757, ZN => n23315);
   U20777 : OAI221_X1 port map( B1 => n21127, B2 => n25042, C1 => n20363, C2 =>
                           n25036, A => n23323, ZN => n23320);
   U20778 : AOI22_X1 port map( A1 => n25030, A2 => n24383, B1 => n25024, B2 => 
                           n17770, ZN => n23323);
   U20779 : OAI221_X1 port map( B1 => n9443, B2 => n25144, C1 => n20426, C2 => 
                           n25138, A => n23297, ZN => n23294);
   U20780 : AOI22_X1 port map( A1 => n25132, A2 => n24053, B1 => n25126, B2 => 
                           n17736, ZN => n23297);
   U20781 : OAI221_X1 port map( B1 => n21126, B2 => n25042, C1 => n20362, C2 =>
                           n25036, A => n23305, ZN => n23302);
   U20782 : AOI22_X1 port map( A1 => n25030, A2 => n24385, B1 => n25024, B2 => 
                           n17749, ZN => n23305);
   U20783 : OAI221_X1 port map( B1 => n9442, B2 => n25145, C1 => n20425, C2 => 
                           n25139, A => n23279, ZN => n23276);
   U20784 : AOI22_X1 port map( A1 => n25133, A2 => n24054, B1 => n25127, B2 => 
                           n17715, ZN => n23279);
   U20785 : OAI221_X1 port map( B1 => n21125, B2 => n25043, C1 => n20361, C2 =>
                           n25037, A => n23287, ZN => n23284);
   U20786 : AOI22_X1 port map( A1 => n25031, A2 => n24387, B1 => n25025, B2 => 
                           n17728, ZN => n23287);
   U20787 : OAI221_X1 port map( B1 => n9441, B2 => n25145, C1 => n20424, C2 => 
                           n25139, A => n23261, ZN => n23258);
   U20788 : AOI22_X1 port map( A1 => n25133, A2 => n24055, B1 => n25127, B2 => 
                           n17694, ZN => n23261);
   U20789 : OAI221_X1 port map( B1 => n21124, B2 => n25043, C1 => n20360, C2 =>
                           n25037, A => n23269, ZN => n23266);
   U20790 : AOI22_X1 port map( A1 => n25031, A2 => n24389, B1 => n25025, B2 => 
                           n17707, ZN => n23269);
   U20791 : OAI221_X1 port map( B1 => n9440, B2 => n25145, C1 => n20423, C2 => 
                           n25139, A => n23243, ZN => n23240);
   U20792 : AOI22_X1 port map( A1 => n25133, A2 => n24056, B1 => n25127, B2 => 
                           n17673, ZN => n23243);
   U20793 : OAI221_X1 port map( B1 => n21123, B2 => n25043, C1 => n20359, C2 =>
                           n25037, A => n23251, ZN => n23248);
   U20794 : AOI22_X1 port map( A1 => n25031, A2 => n24391, B1 => n25025, B2 => 
                           n17686, ZN => n23251);
   U20795 : OAI221_X1 port map( B1 => n9439, B2 => n25145, C1 => n20422, C2 => 
                           n25139, A => n23225, ZN => n23222);
   U20796 : AOI22_X1 port map( A1 => n25133, A2 => n24057, B1 => n25127, B2 => 
                           n17652, ZN => n23225);
   U20797 : OAI221_X1 port map( B1 => n21122, B2 => n25043, C1 => n20358, C2 =>
                           n25037, A => n23233, ZN => n23230);
   U20798 : AOI22_X1 port map( A1 => n25031, A2 => n24393, B1 => n25025, B2 => 
                           n17665, ZN => n23233);
   U20799 : OAI221_X1 port map( B1 => n9438, B2 => n25145, C1 => n20421, C2 => 
                           n25139, A => n23207, ZN => n23204);
   U20800 : AOI22_X1 port map( A1 => n25133, A2 => n24058, B1 => n25127, B2 => 
                           n17631, ZN => n23207);
   U20801 : OAI221_X1 port map( B1 => n21121, B2 => n25043, C1 => n20357, C2 =>
                           n25037, A => n23215, ZN => n23212);
   U20802 : AOI22_X1 port map( A1 => n25031, A2 => n24395, B1 => n25025, B2 => 
                           n17644, ZN => n23215);
   U20803 : OAI221_X1 port map( B1 => n9437, B2 => n25145, C1 => n20420, C2 => 
                           n25139, A => n23189, ZN => n23186);
   U20804 : AOI22_X1 port map( A1 => n25133, A2 => n24059, B1 => n25127, B2 => 
                           n17610, ZN => n23189);
   U20805 : OAI221_X1 port map( B1 => n21120, B2 => n25043, C1 => n20356, C2 =>
                           n25037, A => n23197, ZN => n23194);
   U20806 : AOI22_X1 port map( A1 => n25031, A2 => n24397, B1 => n25025, B2 => 
                           n17623, ZN => n23197);
   U20807 : OAI221_X1 port map( B1 => n9436, B2 => n25145, C1 => n20419, C2 => 
                           n25139, A => n23171, ZN => n23168);
   U20808 : AOI22_X1 port map( A1 => n25133, A2 => n24060, B1 => n25127, B2 => 
                           n17589, ZN => n23171);
   U20809 : OAI221_X1 port map( B1 => n21119, B2 => n25043, C1 => n20355, C2 =>
                           n25037, A => n23179, ZN => n23176);
   U20810 : AOI22_X1 port map( A1 => n25031, A2 => n24399, B1 => n25025, B2 => 
                           n17602, ZN => n23179);
   U20811 : OAI221_X1 port map( B1 => n9435, B2 => n25145, C1 => n20418, C2 => 
                           n25139, A => n23153, ZN => n23150);
   U20812 : AOI22_X1 port map( A1 => n25133, A2 => n24061, B1 => n25127, B2 => 
                           n17568, ZN => n23153);
   U20813 : OAI221_X1 port map( B1 => n21118, B2 => n25043, C1 => n20354, C2 =>
                           n25037, A => n23161, ZN => n23158);
   U20814 : AOI22_X1 port map( A1 => n25031, A2 => n24401, B1 => n25025, B2 => 
                           n17581, ZN => n23161);
   U20815 : OAI221_X1 port map( B1 => n9434, B2 => n25145, C1 => n20417, C2 => 
                           n25139, A => n23135, ZN => n23132);
   U20816 : AOI22_X1 port map( A1 => n25133, A2 => n24062, B1 => n25127, B2 => 
                           n17547, ZN => n23135);
   U20817 : OAI221_X1 port map( B1 => n21117, B2 => n25043, C1 => n20353, C2 =>
                           n25037, A => n23143, ZN => n23140);
   U20818 : AOI22_X1 port map( A1 => n25031, A2 => n24403, B1 => n25025, B2 => 
                           n17560, ZN => n23143);
   U20819 : OAI221_X1 port map( B1 => n9433, B2 => n25145, C1 => n20416, C2 => 
                           n25139, A => n23117, ZN => n23114);
   U20820 : AOI22_X1 port map( A1 => n25133, A2 => n24063, B1 => n25127, B2 => 
                           n17526, ZN => n23117);
   U20821 : OAI221_X1 port map( B1 => n21116, B2 => n25043, C1 => n20352, C2 =>
                           n25037, A => n23125, ZN => n23122);
   U20822 : AOI22_X1 port map( A1 => n25031, A2 => n24405, B1 => n25025, B2 => 
                           n17539, ZN => n23125);
   U20823 : OAI221_X1 port map( B1 => n9432, B2 => n25145, C1 => n20415, C2 => 
                           n25139, A => n23099, ZN => n23096);
   U20824 : AOI22_X1 port map( A1 => n25133, A2 => n24064, B1 => n25127, B2 => 
                           n17505, ZN => n23099);
   U20825 : OAI221_X1 port map( B1 => n21115, B2 => n25043, C1 => n20351, C2 =>
                           n25037, A => n23107, ZN => n23104);
   U20826 : AOI22_X1 port map( A1 => n25031, A2 => n24407, B1 => n25025, B2 => 
                           n17518, ZN => n23107);
   U20827 : OAI221_X1 port map( B1 => n9431, B2 => n25145, C1 => n20414, C2 => 
                           n25139, A => n23081, ZN => n23078);
   U20828 : AOI22_X1 port map( A1 => n25133, A2 => n24065, B1 => n25127, B2 => 
                           n17484, ZN => n23081);
   U20829 : OAI221_X1 port map( B1 => n21114, B2 => n25043, C1 => n20350, C2 =>
                           n25037, A => n23089, ZN => n23086);
   U20830 : AOI22_X1 port map( A1 => n25031, A2 => n24409, B1 => n25025, B2 => 
                           n17497, ZN => n23089);
   U20831 : OAI221_X1 port map( B1 => n9430, B2 => n25146, C1 => n20413, C2 => 
                           n25140, A => n23063, ZN => n23060);
   U20832 : AOI22_X1 port map( A1 => n25134, A2 => n24066, B1 => n25128, B2 => 
                           n17463, ZN => n23063);
   U20833 : OAI221_X1 port map( B1 => n21113, B2 => n25044, C1 => n20349, C2 =>
                           n25038, A => n23071, ZN => n23068);
   U20834 : AOI22_X1 port map( A1 => n25032, A2 => n24411, B1 => n25026, B2 => 
                           n17476, ZN => n23071);
   U20835 : OAI221_X1 port map( B1 => n9429, B2 => n25146, C1 => n20412, C2 => 
                           n25140, A => n23045, ZN => n23042);
   U20836 : AOI22_X1 port map( A1 => n25134, A2 => n24067, B1 => n25128, B2 => 
                           n17442, ZN => n23045);
   U20837 : OAI221_X1 port map( B1 => n21112, B2 => n25044, C1 => n20348, C2 =>
                           n25038, A => n23053, ZN => n23050);
   U20838 : AOI22_X1 port map( A1 => n25032, A2 => n24413, B1 => n25026, B2 => 
                           n17455, ZN => n23053);
   U20839 : OAI221_X1 port map( B1 => n9428, B2 => n25146, C1 => n20411, C2 => 
                           n25140, A => n23027, ZN => n23024);
   U20840 : AOI22_X1 port map( A1 => n25134, A2 => n24068, B1 => n25128, B2 => 
                           n17421, ZN => n23027);
   U20841 : OAI221_X1 port map( B1 => n21111, B2 => n25044, C1 => n20347, C2 =>
                           n25038, A => n23035, ZN => n23032);
   U20842 : AOI22_X1 port map( A1 => n25032, A2 => n24415, B1 => n25026, B2 => 
                           n17434, ZN => n23035);
   U20843 : OAI221_X1 port map( B1 => n9427, B2 => n25146, C1 => n20410, C2 => 
                           n25140, A => n23009, ZN => n23006);
   U20844 : AOI22_X1 port map( A1 => n25134, A2 => n24069, B1 => n25128, B2 => 
                           n17400, ZN => n23009);
   U20845 : OAI221_X1 port map( B1 => n21110, B2 => n25044, C1 => n20346, C2 =>
                           n25038, A => n23017, ZN => n23014);
   U20846 : AOI22_X1 port map( A1 => n25032, A2 => n24417, B1 => n25026, B2 => 
                           n17413, ZN => n23017);
   U20847 : OAI221_X1 port map( B1 => n9426, B2 => n25146, C1 => n20409, C2 => 
                           n25140, A => n22991, ZN => n22988);
   U20848 : AOI22_X1 port map( A1 => n25134, A2 => n24070, B1 => n25128, B2 => 
                           n17379, ZN => n22991);
   U20849 : OAI221_X1 port map( B1 => n21109, B2 => n25044, C1 => n20345, C2 =>
                           n25038, A => n22999, ZN => n22996);
   U20850 : AOI22_X1 port map( A1 => n25032, A2 => n24419, B1 => n25026, B2 => 
                           n17392, ZN => n22999);
   U20851 : OAI221_X1 port map( B1 => n9425, B2 => n25146, C1 => n20408, C2 => 
                           n25140, A => n22973, ZN => n22970);
   U20852 : AOI22_X1 port map( A1 => n25134, A2 => n24071, B1 => n25128, B2 => 
                           n17358, ZN => n22973);
   U20853 : OAI221_X1 port map( B1 => n21108, B2 => n25044, C1 => n20344, C2 =>
                           n25038, A => n22981, ZN => n22978);
   U20854 : AOI22_X1 port map( A1 => n25032, A2 => n24421, B1 => n25026, B2 => 
                           n17371, ZN => n22981);
   U20855 : OAI221_X1 port map( B1 => n9424, B2 => n25146, C1 => n20407, C2 => 
                           n25140, A => n22955, ZN => n22952);
   U20856 : AOI22_X1 port map( A1 => n25134, A2 => n24072, B1 => n25128, B2 => 
                           n17337, ZN => n22955);
   U20857 : OAI221_X1 port map( B1 => n21107, B2 => n25044, C1 => n20343, C2 =>
                           n25038, A => n22963, ZN => n22960);
   U20858 : AOI22_X1 port map( A1 => n25032, A2 => n24423, B1 => n25026, B2 => 
                           n17350, ZN => n22963);
   U20859 : OAI221_X1 port map( B1 => n9423, B2 => n25146, C1 => n20406, C2 => 
                           n25140, A => n22937, ZN => n22934);
   U20860 : AOI22_X1 port map( A1 => n25134, A2 => n24073, B1 => n25128, B2 => 
                           n17316, ZN => n22937);
   U20861 : OAI221_X1 port map( B1 => n21106, B2 => n25044, C1 => n20342, C2 =>
                           n25038, A => n22945, ZN => n22942);
   U20862 : AOI22_X1 port map( A1 => n25032, A2 => n24425, B1 => n25026, B2 => 
                           n17329, ZN => n22945);
   U20863 : OAI221_X1 port map( B1 => n9422, B2 => n25146, C1 => n20405, C2 => 
                           n25140, A => n22919, ZN => n22916);
   U20864 : AOI22_X1 port map( A1 => n25134, A2 => n24074, B1 => n25128, B2 => 
                           n17295, ZN => n22919);
   U20865 : OAI221_X1 port map( B1 => n21105, B2 => n25044, C1 => n20341, C2 =>
                           n25038, A => n22927, ZN => n22924);
   U20866 : AOI22_X1 port map( A1 => n25032, A2 => n24427, B1 => n25026, B2 => 
                           n17308, ZN => n22927);
   U20867 : OAI221_X1 port map( B1 => n9421, B2 => n25146, C1 => n20404, C2 => 
                           n25140, A => n22901, ZN => n22898);
   U20868 : AOI22_X1 port map( A1 => n25134, A2 => n24075, B1 => n25128, B2 => 
                           n17274, ZN => n22901);
   U20869 : OAI221_X1 port map( B1 => n21104, B2 => n25044, C1 => n20340, C2 =>
                           n25038, A => n22909, ZN => n22906);
   U20870 : AOI22_X1 port map( A1 => n25032, A2 => n24429, B1 => n25026, B2 => 
                           n17287, ZN => n22909);
   U20871 : OAI221_X1 port map( B1 => n9420, B2 => n25146, C1 => n20403, C2 => 
                           n25140, A => n22883, ZN => n22880);
   U20872 : AOI22_X1 port map( A1 => n25134, A2 => n24076, B1 => n25128, B2 => 
                           n17253, ZN => n22883);
   U20873 : OAI221_X1 port map( B1 => n21103, B2 => n25044, C1 => n20339, C2 =>
                           n25038, A => n22891, ZN => n22888);
   U20874 : AOI22_X1 port map( A1 => n25032, A2 => n24431, B1 => n25026, B2 => 
                           n17266, ZN => n22891);
   U20875 : OAI221_X1 port map( B1 => n9419, B2 => n25146, C1 => n20402, C2 => 
                           n25140, A => n22865, ZN => n22862);
   U20876 : AOI22_X1 port map( A1 => n25134, A2 => n24077, B1 => n25128, B2 => 
                           n17232, ZN => n22865);
   U20877 : OAI221_X1 port map( B1 => n21102, B2 => n25044, C1 => n20338, C2 =>
                           n25038, A => n22873, ZN => n22870);
   U20878 : AOI22_X1 port map( A1 => n25032, A2 => n24433, B1 => n25026, B2 => 
                           n17245, ZN => n22873);
   U20879 : OAI221_X1 port map( B1 => n9466, B2 => n25341, C1 => n20449, C2 => 
                           n25335, A => n22514, ZN => n22511);
   U20880 : AOI22_X1 port map( A1 => n25329, A2 => n24030, B1 => n25323, B2 => 
                           n18219, ZN => n22514);
   U20881 : OAI221_X1 port map( B1 => n21149, B2 => n25239, C1 => n20385, C2 =>
                           n25233, A => n22522, ZN => n22519);
   U20882 : AOI22_X1 port map( A1 => n25227, A2 => n24339, B1 => n25221, B2 => 
                           n18232, ZN => n22522);
   U20883 : OAI221_X1 port map( B1 => n9465, B2 => n25341, C1 => n20448, C2 => 
                           n25335, A => n22496, ZN => n22493);
   U20884 : AOI22_X1 port map( A1 => n25329, A2 => n24031, B1 => n25323, B2 => 
                           n18198, ZN => n22496);
   U20885 : OAI221_X1 port map( B1 => n21148, B2 => n25239, C1 => n20384, C2 =>
                           n25233, A => n22504, ZN => n22501);
   U20886 : AOI22_X1 port map( A1 => n25227, A2 => n24341, B1 => n25221, B2 => 
                           n18211, ZN => n22504);
   U20887 : OAI221_X1 port map( B1 => n9464, B2 => n25341, C1 => n20447, C2 => 
                           n25335, A => n22478, ZN => n22475);
   U20888 : AOI22_X1 port map( A1 => n25329, A2 => n24032, B1 => n25323, B2 => 
                           n18177, ZN => n22478);
   U20889 : OAI221_X1 port map( B1 => n21147, B2 => n25239, C1 => n20383, C2 =>
                           n25233, A => n22486, ZN => n22483);
   U20890 : AOI22_X1 port map( A1 => n25227, A2 => n24343, B1 => n25221, B2 => 
                           n18190, ZN => n22486);
   U20891 : OAI221_X1 port map( B1 => n9463, B2 => n25341, C1 => n20446, C2 => 
                           n25335, A => n22460, ZN => n22457);
   U20892 : AOI22_X1 port map( A1 => n25329, A2 => n24033, B1 => n25323, B2 => 
                           n18156, ZN => n22460);
   U20893 : OAI221_X1 port map( B1 => n21146, B2 => n25239, C1 => n20382, C2 =>
                           n25233, A => n22468, ZN => n22465);
   U20894 : AOI22_X1 port map( A1 => n25227, A2 => n24345, B1 => n25221, B2 => 
                           n18169, ZN => n22468);
   U20895 : OAI221_X1 port map( B1 => n9462, B2 => n25341, C1 => n20445, C2 => 
                           n25335, A => n22442, ZN => n22439);
   U20896 : AOI22_X1 port map( A1 => n25329, A2 => n24034, B1 => n25323, B2 => 
                           n18135, ZN => n22442);
   U20897 : OAI221_X1 port map( B1 => n21145, B2 => n25239, C1 => n20381, C2 =>
                           n25233, A => n22450, ZN => n22447);
   U20898 : AOI22_X1 port map( A1 => n25227, A2 => n24347, B1 => n25221, B2 => 
                           n18148, ZN => n22450);
   U20899 : OAI221_X1 port map( B1 => n9461, B2 => n25341, C1 => n20444, C2 => 
                           n25335, A => n22424, ZN => n22421);
   U20900 : AOI22_X1 port map( A1 => n25329, A2 => n24035, B1 => n25323, B2 => 
                           n18114, ZN => n22424);
   U20901 : OAI221_X1 port map( B1 => n21144, B2 => n25239, C1 => n20380, C2 =>
                           n25233, A => n22432, ZN => n22429);
   U20902 : AOI22_X1 port map( A1 => n25227, A2 => n24349, B1 => n25221, B2 => 
                           n18127, ZN => n22432);
   U20903 : OAI221_X1 port map( B1 => n9460, B2 => n25341, C1 => n20443, C2 => 
                           n25335, A => n22406, ZN => n22403);
   U20904 : AOI22_X1 port map( A1 => n25329, A2 => n24036, B1 => n25323, B2 => 
                           n18093, ZN => n22406);
   U20905 : OAI221_X1 port map( B1 => n21143, B2 => n25239, C1 => n20379, C2 =>
                           n25233, A => n22414, ZN => n22411);
   U20906 : AOI22_X1 port map( A1 => n25227, A2 => n24351, B1 => n25221, B2 => 
                           n18106, ZN => n22414);
   U20907 : OAI221_X1 port map( B1 => n9459, B2 => n25341, C1 => n20442, C2 => 
                           n25335, A => n22388, ZN => n22385);
   U20908 : AOI22_X1 port map( A1 => n25329, A2 => n24037, B1 => n25323, B2 => 
                           n18072, ZN => n22388);
   U20909 : OAI221_X1 port map( B1 => n21142, B2 => n25239, C1 => n20378, C2 =>
                           n25233, A => n22396, ZN => n22393);
   U20910 : AOI22_X1 port map( A1 => n25227, A2 => n24353, B1 => n25221, B2 => 
                           n18085, ZN => n22396);
   U20911 : OAI221_X1 port map( B1 => n9458, B2 => n25341, C1 => n20441, C2 => 
                           n25335, A => n22370, ZN => n22367);
   U20912 : AOI22_X1 port map( A1 => n25329, A2 => n24038, B1 => n25323, B2 => 
                           n18051, ZN => n22370);
   U20913 : OAI221_X1 port map( B1 => n21141, B2 => n25239, C1 => n20377, C2 =>
                           n25233, A => n22378, ZN => n22375);
   U20914 : AOI22_X1 port map( A1 => n25227, A2 => n24355, B1 => n25221, B2 => 
                           n18064, ZN => n22378);
   U20915 : OAI221_X1 port map( B1 => n9457, B2 => n25341, C1 => n20440, C2 => 
                           n25335, A => n22352, ZN => n22349);
   U20916 : AOI22_X1 port map( A1 => n25329, A2 => n24039, B1 => n25323, B2 => 
                           n18030, ZN => n22352);
   U20917 : OAI221_X1 port map( B1 => n21140, B2 => n25239, C1 => n20376, C2 =>
                           n25233, A => n22360, ZN => n22357);
   U20918 : AOI22_X1 port map( A1 => n25227, A2 => n24357, B1 => n25221, B2 => 
                           n18043, ZN => n22360);
   U20919 : OAI221_X1 port map( B1 => n9456, B2 => n25341, C1 => n20439, C2 => 
                           n25335, A => n22334, ZN => n22331);
   U20920 : AOI22_X1 port map( A1 => n25329, A2 => n24040, B1 => n25323, B2 => 
                           n18009, ZN => n22334);
   U20921 : OAI221_X1 port map( B1 => n21139, B2 => n25239, C1 => n20375, C2 =>
                           n25233, A => n22342, ZN => n22339);
   U20922 : AOI22_X1 port map( A1 => n25227, A2 => n24359, B1 => n25221, B2 => 
                           n18022, ZN => n22342);
   U20923 : OAI221_X1 port map( B1 => n9455, B2 => n25341, C1 => n20438, C2 => 
                           n25335, A => n22316, ZN => n22313);
   U20924 : AOI22_X1 port map( A1 => n25329, A2 => n24041, B1 => n25323, B2 => 
                           n17988, ZN => n22316);
   U20925 : OAI221_X1 port map( B1 => n21138, B2 => n25239, C1 => n20374, C2 =>
                           n25233, A => n22324, ZN => n22321);
   U20926 : AOI22_X1 port map( A1 => n25227, A2 => n24361, B1 => n25221, B2 => 
                           n18001, ZN => n22324);
   U20927 : OAI221_X1 port map( B1 => n9454, B2 => n25342, C1 => n20437, C2 => 
                           n25336, A => n22298, ZN => n22295);
   U20928 : AOI22_X1 port map( A1 => n25330, A2 => n24042, B1 => n25324, B2 => 
                           n17967, ZN => n22298);
   U20929 : OAI221_X1 port map( B1 => n21137, B2 => n25240, C1 => n20373, C2 =>
                           n25234, A => n22306, ZN => n22303);
   U20930 : AOI22_X1 port map( A1 => n25228, A2 => n24363, B1 => n25222, B2 => 
                           n17980, ZN => n22306);
   U20931 : OAI221_X1 port map( B1 => n9453, B2 => n25342, C1 => n20436, C2 => 
                           n25336, A => n22280, ZN => n22277);
   U20932 : AOI22_X1 port map( A1 => n25330, A2 => n24043, B1 => n25324, B2 => 
                           n17946, ZN => n22280);
   U20933 : OAI221_X1 port map( B1 => n21136, B2 => n25240, C1 => n20372, C2 =>
                           n25234, A => n22288, ZN => n22285);
   U20934 : AOI22_X1 port map( A1 => n25228, A2 => n24365, B1 => n25222, B2 => 
                           n17959, ZN => n22288);
   U20935 : OAI221_X1 port map( B1 => n9452, B2 => n25342, C1 => n20435, C2 => 
                           n25336, A => n22262, ZN => n22259);
   U20936 : AOI22_X1 port map( A1 => n25330, A2 => n24044, B1 => n25324, B2 => 
                           n17925, ZN => n22262);
   U20937 : OAI221_X1 port map( B1 => n21135, B2 => n25240, C1 => n20371, C2 =>
                           n25234, A => n22270, ZN => n22267);
   U20938 : AOI22_X1 port map( A1 => n25228, A2 => n24367, B1 => n25222, B2 => 
                           n17938, ZN => n22270);
   U20939 : OAI221_X1 port map( B1 => n9451, B2 => n25342, C1 => n20434, C2 => 
                           n25336, A => n22244, ZN => n22241);
   U20940 : AOI22_X1 port map( A1 => n25330, A2 => n24045, B1 => n25324, B2 => 
                           n17904, ZN => n22244);
   U20941 : OAI221_X1 port map( B1 => n21134, B2 => n25240, C1 => n20370, C2 =>
                           n25234, A => n22252, ZN => n22249);
   U20942 : AOI22_X1 port map( A1 => n25228, A2 => n24369, B1 => n25222, B2 => 
                           n17917, ZN => n22252);
   U20943 : OAI221_X1 port map( B1 => n9450, B2 => n25342, C1 => n20433, C2 => 
                           n25336, A => n22226, ZN => n22223);
   U20944 : AOI22_X1 port map( A1 => n25330, A2 => n24046, B1 => n25324, B2 => 
                           n17883, ZN => n22226);
   U20945 : OAI221_X1 port map( B1 => n21133, B2 => n25240, C1 => n20369, C2 =>
                           n25234, A => n22234, ZN => n22231);
   U20946 : AOI22_X1 port map( A1 => n25228, A2 => n24371, B1 => n25222, B2 => 
                           n17896, ZN => n22234);
   U20947 : OAI221_X1 port map( B1 => n9449, B2 => n25342, C1 => n20432, C2 => 
                           n25336, A => n22208, ZN => n22205);
   U20948 : AOI22_X1 port map( A1 => n25330, A2 => n24047, B1 => n25324, B2 => 
                           n17862, ZN => n22208);
   U20949 : OAI221_X1 port map( B1 => n21132, B2 => n25240, C1 => n20368, C2 =>
                           n25234, A => n22216, ZN => n22213);
   U20950 : AOI22_X1 port map( A1 => n25228, A2 => n24373, B1 => n25222, B2 => 
                           n17875, ZN => n22216);
   U20951 : OAI221_X1 port map( B1 => n9448, B2 => n25342, C1 => n20431, C2 => 
                           n25336, A => n22190, ZN => n22187);
   U20952 : AOI22_X1 port map( A1 => n25330, A2 => n24048, B1 => n25324, B2 => 
                           n17841, ZN => n22190);
   U20953 : OAI221_X1 port map( B1 => n21131, B2 => n25240, C1 => n20367, C2 =>
                           n25234, A => n22198, ZN => n22195);
   U20954 : AOI22_X1 port map( A1 => n25228, A2 => n24375, B1 => n25222, B2 => 
                           n17854, ZN => n22198);
   U20955 : OAI221_X1 port map( B1 => n9447, B2 => n25342, C1 => n20430, C2 => 
                           n25336, A => n22172, ZN => n22169);
   U20956 : AOI22_X1 port map( A1 => n25330, A2 => n24049, B1 => n25324, B2 => 
                           n17820, ZN => n22172);
   U20957 : OAI221_X1 port map( B1 => n21130, B2 => n25240, C1 => n20366, C2 =>
                           n25234, A => n22180, ZN => n22177);
   U20958 : AOI22_X1 port map( A1 => n25228, A2 => n24377, B1 => n25222, B2 => 
                           n17833, ZN => n22180);
   U20959 : OAI221_X1 port map( B1 => n9446, B2 => n25342, C1 => n20429, C2 => 
                           n25336, A => n22154, ZN => n22151);
   U20960 : AOI22_X1 port map( A1 => n25330, A2 => n24050, B1 => n25324, B2 => 
                           n17799, ZN => n22154);
   U20961 : OAI221_X1 port map( B1 => n21129, B2 => n25240, C1 => n20365, C2 =>
                           n25234, A => n22162, ZN => n22159);
   U20962 : AOI22_X1 port map( A1 => n25228, A2 => n24379, B1 => n25222, B2 => 
                           n17812, ZN => n22162);
   U20963 : OAI221_X1 port map( B1 => n9445, B2 => n25342, C1 => n20428, C2 => 
                           n25336, A => n22136, ZN => n22133);
   U20964 : AOI22_X1 port map( A1 => n25330, A2 => n24051, B1 => n25324, B2 => 
                           n17778, ZN => n22136);
   U20965 : OAI221_X1 port map( B1 => n21128, B2 => n25240, C1 => n20364, C2 =>
                           n25234, A => n22144, ZN => n22141);
   U20966 : AOI22_X1 port map( A1 => n25228, A2 => n24381, B1 => n25222, B2 => 
                           n17791, ZN => n22144);
   U20967 : OAI221_X1 port map( B1 => n9444, B2 => n25342, C1 => n20427, C2 => 
                           n25336, A => n22118, ZN => n22115);
   U20968 : AOI22_X1 port map( A1 => n25330, A2 => n24052, B1 => n25324, B2 => 
                           n17757, ZN => n22118);
   U20969 : OAI221_X1 port map( B1 => n21127, B2 => n25240, C1 => n20363, C2 =>
                           n25234, A => n22126, ZN => n22123);
   U20970 : AOI22_X1 port map( A1 => n25228, A2 => n24383, B1 => n25222, B2 => 
                           n17770, ZN => n22126);
   U20971 : OAI221_X1 port map( B1 => n9443, B2 => n25342, C1 => n20426, C2 => 
                           n25336, A => n22100, ZN => n22097);
   U20972 : AOI22_X1 port map( A1 => n25330, A2 => n24053, B1 => n25324, B2 => 
                           n17736, ZN => n22100);
   U20973 : OAI221_X1 port map( B1 => n21126, B2 => n25240, C1 => n20362, C2 =>
                           n25234, A => n22108, ZN => n22105);
   U20974 : AOI22_X1 port map( A1 => n25228, A2 => n24385, B1 => n25222, B2 => 
                           n17749, ZN => n22108);
   U20975 : OAI221_X1 port map( B1 => n9442, B2 => n25343, C1 => n20425, C2 => 
                           n25337, A => n22082, ZN => n22079);
   U20976 : AOI22_X1 port map( A1 => n25331, A2 => n24054, B1 => n25325, B2 => 
                           n17715, ZN => n22082);
   U20977 : OAI221_X1 port map( B1 => n21125, B2 => n25241, C1 => n20361, C2 =>
                           n25235, A => n22090, ZN => n22087);
   U20978 : AOI22_X1 port map( A1 => n25229, A2 => n24387, B1 => n25223, B2 => 
                           n17728, ZN => n22090);
   U20979 : OAI221_X1 port map( B1 => n9441, B2 => n25343, C1 => n20424, C2 => 
                           n25337, A => n22064, ZN => n22061);
   U20980 : AOI22_X1 port map( A1 => n25331, A2 => n24055, B1 => n25325, B2 => 
                           n17694, ZN => n22064);
   U20981 : OAI221_X1 port map( B1 => n21124, B2 => n25241, C1 => n20360, C2 =>
                           n25235, A => n22072, ZN => n22069);
   U20982 : AOI22_X1 port map( A1 => n25229, A2 => n24389, B1 => n25223, B2 => 
                           n17707, ZN => n22072);
   U20983 : OAI221_X1 port map( B1 => n9440, B2 => n25343, C1 => n20423, C2 => 
                           n25337, A => n22046, ZN => n22043);
   U20984 : AOI22_X1 port map( A1 => n25331, A2 => n24056, B1 => n25325, B2 => 
                           n17673, ZN => n22046);
   U20985 : OAI221_X1 port map( B1 => n21123, B2 => n25241, C1 => n20359, C2 =>
                           n25235, A => n22054, ZN => n22051);
   U20986 : AOI22_X1 port map( A1 => n25229, A2 => n24391, B1 => n25223, B2 => 
                           n17686, ZN => n22054);
   U20987 : OAI221_X1 port map( B1 => n9439, B2 => n25343, C1 => n20422, C2 => 
                           n25337, A => n22028, ZN => n22025);
   U20988 : AOI22_X1 port map( A1 => n25331, A2 => n24057, B1 => n25325, B2 => 
                           n17652, ZN => n22028);
   U20989 : OAI221_X1 port map( B1 => n21122, B2 => n25241, C1 => n20358, C2 =>
                           n25235, A => n22036, ZN => n22033);
   U20990 : AOI22_X1 port map( A1 => n25229, A2 => n24393, B1 => n25223, B2 => 
                           n17665, ZN => n22036);
   U20991 : OAI221_X1 port map( B1 => n9438, B2 => n25343, C1 => n20421, C2 => 
                           n25337, A => n22010, ZN => n22007);
   U20992 : AOI22_X1 port map( A1 => n25331, A2 => n24058, B1 => n25325, B2 => 
                           n17631, ZN => n22010);
   U20993 : OAI221_X1 port map( B1 => n21121, B2 => n25241, C1 => n20357, C2 =>
                           n25235, A => n22018, ZN => n22015);
   U20994 : AOI22_X1 port map( A1 => n25229, A2 => n24395, B1 => n25223, B2 => 
                           n17644, ZN => n22018);
   U20995 : OAI221_X1 port map( B1 => n9437, B2 => n25343, C1 => n20420, C2 => 
                           n25337, A => n21992, ZN => n21989);
   U20996 : AOI22_X1 port map( A1 => n25331, A2 => n24059, B1 => n25325, B2 => 
                           n17610, ZN => n21992);
   U20997 : OAI221_X1 port map( B1 => n21120, B2 => n25241, C1 => n20356, C2 =>
                           n25235, A => n22000, ZN => n21997);
   U20998 : AOI22_X1 port map( A1 => n25229, A2 => n24397, B1 => n25223, B2 => 
                           n17623, ZN => n22000);
   U20999 : OAI221_X1 port map( B1 => n9436, B2 => n25343, C1 => n20419, C2 => 
                           n25337, A => n21974, ZN => n21971);
   U21000 : AOI22_X1 port map( A1 => n25331, A2 => n24060, B1 => n25325, B2 => 
                           n17589, ZN => n21974);
   U21001 : OAI221_X1 port map( B1 => n21119, B2 => n25241, C1 => n20355, C2 =>
                           n25235, A => n21982, ZN => n21979);
   U21002 : AOI22_X1 port map( A1 => n25229, A2 => n24399, B1 => n25223, B2 => 
                           n17602, ZN => n21982);
   U21003 : OAI221_X1 port map( B1 => n9435, B2 => n25343, C1 => n20418, C2 => 
                           n25337, A => n21956, ZN => n21953);
   U21004 : AOI22_X1 port map( A1 => n25331, A2 => n24061, B1 => n25325, B2 => 
                           n17568, ZN => n21956);
   U21005 : OAI221_X1 port map( B1 => n21118, B2 => n25241, C1 => n20354, C2 =>
                           n25235, A => n21964, ZN => n21961);
   U21006 : AOI22_X1 port map( A1 => n25229, A2 => n24401, B1 => n25223, B2 => 
                           n17581, ZN => n21964);
   U21007 : OAI221_X1 port map( B1 => n9434, B2 => n25343, C1 => n20417, C2 => 
                           n25337, A => n21938, ZN => n21935);
   U21008 : AOI22_X1 port map( A1 => n25331, A2 => n24062, B1 => n25325, B2 => 
                           n17547, ZN => n21938);
   U21009 : OAI221_X1 port map( B1 => n21117, B2 => n25241, C1 => n20353, C2 =>
                           n25235, A => n21946, ZN => n21943);
   U21010 : AOI22_X1 port map( A1 => n25229, A2 => n24403, B1 => n25223, B2 => 
                           n17560, ZN => n21946);
   U21011 : OAI221_X1 port map( B1 => n9433, B2 => n25343, C1 => n20416, C2 => 
                           n25337, A => n21920, ZN => n21917);
   U21012 : AOI22_X1 port map( A1 => n25331, A2 => n24063, B1 => n25325, B2 => 
                           n17526, ZN => n21920);
   U21013 : OAI221_X1 port map( B1 => n21116, B2 => n25241, C1 => n20352, C2 =>
                           n25235, A => n21928, ZN => n21925);
   U21014 : AOI22_X1 port map( A1 => n25229, A2 => n24405, B1 => n25223, B2 => 
                           n17539, ZN => n21928);
   U21015 : OAI221_X1 port map( B1 => n9432, B2 => n25343, C1 => n20415, C2 => 
                           n25337, A => n21902, ZN => n21899);
   U21016 : AOI22_X1 port map( A1 => n25331, A2 => n24064, B1 => n25325, B2 => 
                           n17505, ZN => n21902);
   U21017 : OAI221_X1 port map( B1 => n21115, B2 => n25241, C1 => n20351, C2 =>
                           n25235, A => n21910, ZN => n21907);
   U21018 : AOI22_X1 port map( A1 => n25229, A2 => n24407, B1 => n25223, B2 => 
                           n17518, ZN => n21910);
   U21019 : OAI221_X1 port map( B1 => n9431, B2 => n25343, C1 => n20414, C2 => 
                           n25337, A => n21884, ZN => n21881);
   U21020 : AOI22_X1 port map( A1 => n25331, A2 => n24065, B1 => n25325, B2 => 
                           n17484, ZN => n21884);
   U21021 : OAI221_X1 port map( B1 => n21114, B2 => n25241, C1 => n20350, C2 =>
                           n25235, A => n21892, ZN => n21889);
   U21022 : AOI22_X1 port map( A1 => n25229, A2 => n24409, B1 => n25223, B2 => 
                           n17497, ZN => n21892);
   U21023 : OAI221_X1 port map( B1 => n9430, B2 => n25344, C1 => n20413, C2 => 
                           n25338, A => n21866, ZN => n21863);
   U21024 : AOI22_X1 port map( A1 => n25332, A2 => n24066, B1 => n25326, B2 => 
                           n17463, ZN => n21866);
   U21025 : OAI221_X1 port map( B1 => n21113, B2 => n25242, C1 => n20349, C2 =>
                           n25236, A => n21874, ZN => n21871);
   U21026 : AOI22_X1 port map( A1 => n25230, A2 => n24411, B1 => n25224, B2 => 
                           n17476, ZN => n21874);
   U21027 : OAI221_X1 port map( B1 => n9429, B2 => n25344, C1 => n20412, C2 => 
                           n25338, A => n21848, ZN => n21845);
   U21028 : AOI22_X1 port map( A1 => n25332, A2 => n24067, B1 => n25326, B2 => 
                           n17442, ZN => n21848);
   U21029 : OAI221_X1 port map( B1 => n21112, B2 => n25242, C1 => n20348, C2 =>
                           n25236, A => n21856, ZN => n21853);
   U21030 : AOI22_X1 port map( A1 => n25230, A2 => n24413, B1 => n25224, B2 => 
                           n17455, ZN => n21856);
   U21031 : OAI221_X1 port map( B1 => n9428, B2 => n25344, C1 => n20411, C2 => 
                           n25338, A => n21830, ZN => n21827);
   U21032 : AOI22_X1 port map( A1 => n25332, A2 => n24068, B1 => n25326, B2 => 
                           n17421, ZN => n21830);
   U21033 : OAI221_X1 port map( B1 => n21111, B2 => n25242, C1 => n20347, C2 =>
                           n25236, A => n21838, ZN => n21835);
   U21034 : AOI22_X1 port map( A1 => n25230, A2 => n24415, B1 => n25224, B2 => 
                           n17434, ZN => n21838);
   U21035 : OAI221_X1 port map( B1 => n9427, B2 => n25344, C1 => n20410, C2 => 
                           n25338, A => n21812, ZN => n21809);
   U21036 : AOI22_X1 port map( A1 => n25332, A2 => n24069, B1 => n25326, B2 => 
                           n17400, ZN => n21812);
   U21037 : OAI221_X1 port map( B1 => n21110, B2 => n25242, C1 => n20346, C2 =>
                           n25236, A => n21820, ZN => n21817);
   U21038 : AOI22_X1 port map( A1 => n25230, A2 => n24417, B1 => n25224, B2 => 
                           n17413, ZN => n21820);
   U21039 : OAI221_X1 port map( B1 => n9426, B2 => n25344, C1 => n20409, C2 => 
                           n25338, A => n21794, ZN => n21791);
   U21040 : AOI22_X1 port map( A1 => n25332, A2 => n24070, B1 => n25326, B2 => 
                           n17379, ZN => n21794);
   U21041 : OAI221_X1 port map( B1 => n21109, B2 => n25242, C1 => n20345, C2 =>
                           n25236, A => n21802, ZN => n21799);
   U21042 : AOI22_X1 port map( A1 => n25230, A2 => n24419, B1 => n25224, B2 => 
                           n17392, ZN => n21802);
   U21043 : OAI221_X1 port map( B1 => n9425, B2 => n25344, C1 => n20408, C2 => 
                           n25338, A => n21776, ZN => n21773);
   U21044 : AOI22_X1 port map( A1 => n25332, A2 => n24071, B1 => n25326, B2 => 
                           n17358, ZN => n21776);
   U21045 : OAI221_X1 port map( B1 => n21108, B2 => n25242, C1 => n20344, C2 =>
                           n25236, A => n21784, ZN => n21781);
   U21046 : AOI22_X1 port map( A1 => n25230, A2 => n24421, B1 => n25224, B2 => 
                           n17371, ZN => n21784);
   U21047 : OAI221_X1 port map( B1 => n9424, B2 => n25344, C1 => n20407, C2 => 
                           n25338, A => n21758, ZN => n21755);
   U21048 : AOI22_X1 port map( A1 => n25332, A2 => n24072, B1 => n25326, B2 => 
                           n17337, ZN => n21758);
   U21049 : OAI221_X1 port map( B1 => n21107, B2 => n25242, C1 => n20343, C2 =>
                           n25236, A => n21766, ZN => n21763);
   U21050 : AOI22_X1 port map( A1 => n25230, A2 => n24423, B1 => n25224, B2 => 
                           n17350, ZN => n21766);
   U21051 : OAI221_X1 port map( B1 => n9423, B2 => n25344, C1 => n20406, C2 => 
                           n25338, A => n21740, ZN => n21737);
   U21052 : AOI22_X1 port map( A1 => n25332, A2 => n24073, B1 => n25326, B2 => 
                           n17316, ZN => n21740);
   U21053 : OAI221_X1 port map( B1 => n21106, B2 => n25242, C1 => n20342, C2 =>
                           n25236, A => n21748, ZN => n21745);
   U21054 : AOI22_X1 port map( A1 => n25230, A2 => n24425, B1 => n25224, B2 => 
                           n17329, ZN => n21748);
   U21055 : OAI221_X1 port map( B1 => n9422, B2 => n25344, C1 => n20405, C2 => 
                           n25338, A => n21722, ZN => n21719);
   U21056 : AOI22_X1 port map( A1 => n25332, A2 => n24074, B1 => n25326, B2 => 
                           n17295, ZN => n21722);
   U21057 : OAI221_X1 port map( B1 => n21105, B2 => n25242, C1 => n20341, C2 =>
                           n25236, A => n21730, ZN => n21727);
   U21058 : AOI22_X1 port map( A1 => n25230, A2 => n24427, B1 => n25224, B2 => 
                           n17308, ZN => n21730);
   U21059 : OAI221_X1 port map( B1 => n9421, B2 => n25344, C1 => n20404, C2 => 
                           n25338, A => n21704, ZN => n21701);
   U21060 : AOI22_X1 port map( A1 => n25332, A2 => n24075, B1 => n25326, B2 => 
                           n17274, ZN => n21704);
   U21061 : OAI221_X1 port map( B1 => n21104, B2 => n25242, C1 => n20340, C2 =>
                           n25236, A => n21712, ZN => n21709);
   U21062 : AOI22_X1 port map( A1 => n25230, A2 => n24429, B1 => n25224, B2 => 
                           n17287, ZN => n21712);
   U21063 : OAI221_X1 port map( B1 => n9420, B2 => n25344, C1 => n20403, C2 => 
                           n25338, A => n21686, ZN => n21683);
   U21064 : AOI22_X1 port map( A1 => n25332, A2 => n24076, B1 => n25326, B2 => 
                           n17253, ZN => n21686);
   U21065 : OAI221_X1 port map( B1 => n21103, B2 => n25242, C1 => n20339, C2 =>
                           n25236, A => n21694, ZN => n21691);
   U21066 : AOI22_X1 port map( A1 => n25230, A2 => n24431, B1 => n25224, B2 => 
                           n17266, ZN => n21694);
   U21067 : OAI221_X1 port map( B1 => n9419, B2 => n25344, C1 => n20402, C2 => 
                           n25338, A => n21668, ZN => n21665);
   U21068 : AOI22_X1 port map( A1 => n25332, A2 => n24077, B1 => n25326, B2 => 
                           n17232, ZN => n21668);
   U21069 : OAI221_X1 port map( B1 => n21102, B2 => n25242, C1 => n20338, C2 =>
                           n25236, A => n21676, ZN => n21673);
   U21070 : AOI22_X1 port map( A1 => n25230, A2 => n24433, B1 => n25224, B2 => 
                           n17245, ZN => n21676);
   U21071 : OAI221_X1 port map( B1 => n9415, B2 => n25147, C1 => n20398, C2 => 
                           n25141, A => n22766, ZN => n22757);
   U21072 : AOI22_X1 port map( A1 => n25135, A2 => n23957, B1 => n25129, B2 => 
                           n17148, ZN => n22766);
   U21073 : OAI221_X1 port map( B1 => n21094, B2 => n25045, C1 => n20334, C2 =>
                           n25039, A => n22791, ZN => n22782);
   U21074 : AOI22_X1 port map( A1 => n25033, A2 => n24441, B1 => n25027, B2 => 
                           n17161, ZN => n22791);
   U21075 : OAI221_X1 port map( B1 => n9418, B2 => n25147, C1 => n20401, C2 => 
                           n25141, A => n22847, ZN => n22844);
   U21076 : AOI22_X1 port map( A1 => n25135, A2 => n23954, B1 => n25129, B2 => 
                           n17211, ZN => n22847);
   U21077 : OAI221_X1 port map( B1 => n21097, B2 => n25045, C1 => n20337, C2 =>
                           n25039, A => n22855, ZN => n22852);
   U21078 : AOI22_X1 port map( A1 => n25033, A2 => n24435, B1 => n25027, B2 => 
                           n17224, ZN => n22855);
   U21079 : OAI221_X1 port map( B1 => n9417, B2 => n25147, C1 => n20400, C2 => 
                           n25141, A => n22829, ZN => n22826);
   U21080 : AOI22_X1 port map( A1 => n25135, A2 => n23955, B1 => n25129, B2 => 
                           n17190, ZN => n22829);
   U21081 : OAI221_X1 port map( B1 => n21096, B2 => n25045, C1 => n20336, C2 =>
                           n25039, A => n22837, ZN => n22834);
   U21082 : AOI22_X1 port map( A1 => n25033, A2 => n24437, B1 => n25027, B2 => 
                           n17203, ZN => n22837);
   U21083 : OAI221_X1 port map( B1 => n9416, B2 => n25147, C1 => n20399, C2 => 
                           n25141, A => n22811, ZN => n22808);
   U21084 : AOI22_X1 port map( A1 => n25135, A2 => n23956, B1 => n25129, B2 => 
                           n17169, ZN => n22811);
   U21085 : OAI221_X1 port map( B1 => n21095, B2 => n25045, C1 => n20335, C2 =>
                           n25039, A => n22819, ZN => n22816);
   U21086 : AOI22_X1 port map( A1 => n25033, A2 => n24439, B1 => n25027, B2 => 
                           n17182, ZN => n22819);
   U21087 : OAI221_X1 port map( B1 => n9418, B2 => n25345, C1 => n20401, C2 => 
                           n25339, A => n21650, ZN => n21647);
   U21088 : AOI22_X1 port map( A1 => n25333, A2 => n23954, B1 => n25327, B2 => 
                           n17211, ZN => n21650);
   U21089 : OAI221_X1 port map( B1 => n21097, B2 => n25243, C1 => n20337, C2 =>
                           n25237, A => n21658, ZN => n21655);
   U21090 : AOI22_X1 port map( A1 => n25231, A2 => n24435, B1 => n25225, B2 => 
                           n17224, ZN => n21658);
   U21091 : OAI221_X1 port map( B1 => n9417, B2 => n25345, C1 => n20400, C2 => 
                           n25339, A => n21632, ZN => n21629);
   U21092 : AOI22_X1 port map( A1 => n25333, A2 => n23955, B1 => n25327, B2 => 
                           n17190, ZN => n21632);
   U21093 : OAI221_X1 port map( B1 => n21096, B2 => n25243, C1 => n20336, C2 =>
                           n25237, A => n21640, ZN => n21637);
   U21094 : AOI22_X1 port map( A1 => n25231, A2 => n24437, B1 => n25225, B2 => 
                           n17203, ZN => n21640);
   U21095 : OAI221_X1 port map( B1 => n9416, B2 => n25345, C1 => n20399, C2 => 
                           n25339, A => n21614, ZN => n21611);
   U21096 : AOI22_X1 port map( A1 => n25333, A2 => n23956, B1 => n25327, B2 => 
                           n17169, ZN => n21614);
   U21097 : OAI221_X1 port map( B1 => n21095, B2 => n25243, C1 => n20335, C2 =>
                           n25237, A => n21622, ZN => n21619);
   U21098 : AOI22_X1 port map( A1 => n25231, A2 => n24439, B1 => n25225, B2 => 
                           n17182, ZN => n21622);
   U21099 : OAI221_X1 port map( B1 => n9415, B2 => n25345, C1 => n20398, C2 => 
                           n25339, A => n21569, ZN => n21560);
   U21100 : AOI22_X1 port map( A1 => n25333, A2 => n23957, B1 => n25327, B2 => 
                           n17148, ZN => n21569);
   U21101 : OAI221_X1 port map( B1 => n21094, B2 => n25243, C1 => n20334, C2 =>
                           n25237, A => n21594, ZN => n21585);
   U21102 : AOI22_X1 port map( A1 => n25231, A2 => n24441, B1 => n25225, B2 => 
                           n17161, ZN => n21594);
   U21103 : OAI221_X1 port map( B1 => n9478, B2 => n25142, C1 => n20461, C2 => 
                           n25136, A => n23932, ZN => n23924);
   U21104 : AOI22_X1 port map( A1 => n25130, A2 => n24018, B1 => n25124, B2 => 
                           n18471, ZN => n23932);
   U21105 : OAI221_X1 port map( B1 => n9477, B2 => n25142, C1 => n20460, C2 => 
                           n25136, A => n23909, ZN => n23906);
   U21106 : AOI22_X1 port map( A1 => n25130, A2 => n24019, B1 => n25124, B2 => 
                           n18450, ZN => n23909);
   U21107 : OAI221_X1 port map( B1 => n9476, B2 => n25142, C1 => n20459, C2 => 
                           n25136, A => n23891, ZN => n23888);
   U21108 : AOI22_X1 port map( A1 => n25130, A2 => n24020, B1 => n25124, B2 => 
                           n18429, ZN => n23891);
   U21109 : OAI221_X1 port map( B1 => n9475, B2 => n25142, C1 => n20458, C2 => 
                           n25136, A => n23873, ZN => n23870);
   U21110 : AOI22_X1 port map( A1 => n25130, A2 => n24021, B1 => n25124, B2 => 
                           n18408, ZN => n23873);
   U21111 : OAI221_X1 port map( B1 => n9474, B2 => n25142, C1 => n20457, C2 => 
                           n25136, A => n23855, ZN => n23852);
   U21112 : AOI22_X1 port map( A1 => n25130, A2 => n24022, B1 => n25124, B2 => 
                           n18387, ZN => n23855);
   U21113 : OAI221_X1 port map( B1 => n9473, B2 => n25142, C1 => n20456, C2 => 
                           n25136, A => n23837, ZN => n23834);
   U21114 : AOI22_X1 port map( A1 => n25130, A2 => n24023, B1 => n25124, B2 => 
                           n18366, ZN => n23837);
   U21115 : OAI221_X1 port map( B1 => n9472, B2 => n25142, C1 => n20455, C2 => 
                           n25136, A => n23819, ZN => n23816);
   U21116 : AOI22_X1 port map( A1 => n25130, A2 => n24024, B1 => n25124, B2 => 
                           n18345, ZN => n23819);
   U21117 : OAI221_X1 port map( B1 => n9471, B2 => n25142, C1 => n20454, C2 => 
                           n25136, A => n23801, ZN => n23798);
   U21118 : AOI22_X1 port map( A1 => n25130, A2 => n24025, B1 => n25124, B2 => 
                           n18324, ZN => n23801);
   U21119 : OAI221_X1 port map( B1 => n9470, B2 => n25142, C1 => n20453, C2 => 
                           n25136, A => n23783, ZN => n23780);
   U21120 : AOI22_X1 port map( A1 => n25130, A2 => n24026, B1 => n25124, B2 => 
                           n18303, ZN => n23783);
   U21121 : OAI221_X1 port map( B1 => n9469, B2 => n25142, C1 => n20452, C2 => 
                           n25136, A => n23765, ZN => n23762);
   U21122 : AOI22_X1 port map( A1 => n25130, A2 => n24027, B1 => n25124, B2 => 
                           n18282, ZN => n23765);
   U21123 : OAI221_X1 port map( B1 => n9468, B2 => n25142, C1 => n20451, C2 => 
                           n25136, A => n23747, ZN => n23744);
   U21124 : AOI22_X1 port map( A1 => n25130, A2 => n24028, B1 => n25124, B2 => 
                           n18261, ZN => n23747);
   U21125 : OAI221_X1 port map( B1 => n9467, B2 => n25142, C1 => n20450, C2 => 
                           n25136, A => n23729, ZN => n23726);
   U21126 : AOI22_X1 port map( A1 => n25130, A2 => n24029, B1 => n25124, B2 => 
                           n18240, ZN => n23729);
   U21127 : OAI221_X1 port map( B1 => n9478, B2 => n25340, C1 => n20461, C2 => 
                           n25334, A => n22735, ZN => n22727);
   U21128 : AOI22_X1 port map( A1 => n25328, A2 => n24018, B1 => n25322, B2 => 
                           n18471, ZN => n22735);
   U21129 : OAI221_X1 port map( B1 => n9477, B2 => n25340, C1 => n20460, C2 => 
                           n25334, A => n22712, ZN => n22709);
   U21130 : AOI22_X1 port map( A1 => n25328, A2 => n24019, B1 => n25322, B2 => 
                           n18450, ZN => n22712);
   U21131 : OAI221_X1 port map( B1 => n9476, B2 => n25340, C1 => n20459, C2 => 
                           n25334, A => n22694, ZN => n22691);
   U21132 : AOI22_X1 port map( A1 => n25328, A2 => n24020, B1 => n25322, B2 => 
                           n18429, ZN => n22694);
   U21133 : OAI221_X1 port map( B1 => n9475, B2 => n25340, C1 => n20458, C2 => 
                           n25334, A => n22676, ZN => n22673);
   U21134 : AOI22_X1 port map( A1 => n25328, A2 => n24021, B1 => n25322, B2 => 
                           n18408, ZN => n22676);
   U21135 : OAI221_X1 port map( B1 => n9474, B2 => n25340, C1 => n20457, C2 => 
                           n25334, A => n22658, ZN => n22655);
   U21136 : AOI22_X1 port map( A1 => n25328, A2 => n24022, B1 => n25322, B2 => 
                           n18387, ZN => n22658);
   U21137 : OAI221_X1 port map( B1 => n9473, B2 => n25340, C1 => n20456, C2 => 
                           n25334, A => n22640, ZN => n22637);
   U21138 : AOI22_X1 port map( A1 => n25328, A2 => n24023, B1 => n25322, B2 => 
                           n18366, ZN => n22640);
   U21139 : OAI221_X1 port map( B1 => n9472, B2 => n25340, C1 => n20455, C2 => 
                           n25334, A => n22622, ZN => n22619);
   U21140 : AOI22_X1 port map( A1 => n25328, A2 => n24024, B1 => n25322, B2 => 
                           n18345, ZN => n22622);
   U21141 : OAI221_X1 port map( B1 => n9471, B2 => n25340, C1 => n20454, C2 => 
                           n25334, A => n22604, ZN => n22601);
   U21142 : AOI22_X1 port map( A1 => n25328, A2 => n24025, B1 => n25322, B2 => 
                           n18324, ZN => n22604);
   U21143 : OAI221_X1 port map( B1 => n9470, B2 => n25340, C1 => n20453, C2 => 
                           n25334, A => n22586, ZN => n22583);
   U21144 : AOI22_X1 port map( A1 => n25328, A2 => n24026, B1 => n25322, B2 => 
                           n18303, ZN => n22586);
   U21145 : OAI221_X1 port map( B1 => n9469, B2 => n25340, C1 => n20452, C2 => 
                           n25334, A => n22568, ZN => n22565);
   U21146 : AOI22_X1 port map( A1 => n25328, A2 => n24027, B1 => n25322, B2 => 
                           n18282, ZN => n22568);
   U21147 : OAI221_X1 port map( B1 => n9468, B2 => n25340, C1 => n20451, C2 => 
                           n25334, A => n22550, ZN => n22547);
   U21148 : AOI22_X1 port map( A1 => n25328, A2 => n24028, B1 => n25322, B2 => 
                           n18261, ZN => n22550);
   U21149 : OAI221_X1 port map( B1 => n9467, B2 => n25340, C1 => n20450, C2 => 
                           n25334, A => n22532, ZN => n22529);
   U21150 : AOI22_X1 port map( A1 => n25328, A2 => n24029, B1 => n25322, B2 => 
                           n18240, ZN => n22532);
   U21151 : OAI221_X1 port map( B1 => n21161, B2 => n25040, C1 => n20397, C2 =>
                           n25034, A => n23947, ZN => n23943);
   U21152 : AOI22_X1 port map( A1 => n25028, A2 => n24443, B1 => n25022, B2 => 
                           n18484, ZN => n23947);
   U21153 : OAI221_X1 port map( B1 => n21160, B2 => n25040, C1 => n20396, C2 =>
                           n25034, A => n23917, ZN => n23914);
   U21154 : AOI22_X1 port map( A1 => n25028, A2 => n24445, B1 => n25022, B2 => 
                           n18463, ZN => n23917);
   U21155 : OAI221_X1 port map( B1 => n21159, B2 => n25040, C1 => n20395, C2 =>
                           n25034, A => n23899, ZN => n23896);
   U21156 : AOI22_X1 port map( A1 => n25028, A2 => n24447, B1 => n25022, B2 => 
                           n18442, ZN => n23899);
   U21157 : OAI221_X1 port map( B1 => n21158, B2 => n25040, C1 => n20394, C2 =>
                           n25034, A => n23881, ZN => n23878);
   U21158 : AOI22_X1 port map( A1 => n25028, A2 => n24449, B1 => n25022, B2 => 
                           n18421, ZN => n23881);
   U21159 : OAI221_X1 port map( B1 => n21157, B2 => n25040, C1 => n20393, C2 =>
                           n25034, A => n23863, ZN => n23860);
   U21160 : AOI22_X1 port map( A1 => n25028, A2 => n24451, B1 => n25022, B2 => 
                           n18400, ZN => n23863);
   U21161 : OAI221_X1 port map( B1 => n21156, B2 => n25040, C1 => n20392, C2 =>
                           n25034, A => n23845, ZN => n23842);
   U21162 : AOI22_X1 port map( A1 => n25028, A2 => n24453, B1 => n25022, B2 => 
                           n18379, ZN => n23845);
   U21163 : OAI221_X1 port map( B1 => n21155, B2 => n25040, C1 => n20391, C2 =>
                           n25034, A => n23827, ZN => n23824);
   U21164 : AOI22_X1 port map( A1 => n25028, A2 => n24455, B1 => n25022, B2 => 
                           n18358, ZN => n23827);
   U21165 : OAI221_X1 port map( B1 => n21154, B2 => n25040, C1 => n20390, C2 =>
                           n25034, A => n23809, ZN => n23806);
   U21166 : AOI22_X1 port map( A1 => n25028, A2 => n24457, B1 => n25022, B2 => 
                           n18337, ZN => n23809);
   U21167 : OAI221_X1 port map( B1 => n21153, B2 => n25040, C1 => n20389, C2 =>
                           n25034, A => n23791, ZN => n23788);
   U21168 : AOI22_X1 port map( A1 => n25028, A2 => n24459, B1 => n25022, B2 => 
                           n18316, ZN => n23791);
   U21169 : OAI221_X1 port map( B1 => n21152, B2 => n25040, C1 => n20388, C2 =>
                           n25034, A => n23773, ZN => n23770);
   U21170 : AOI22_X1 port map( A1 => n25028, A2 => n24461, B1 => n25022, B2 => 
                           n18295, ZN => n23773);
   U21171 : OAI221_X1 port map( B1 => n21151, B2 => n25040, C1 => n20387, C2 =>
                           n25034, A => n23755, ZN => n23752);
   U21172 : AOI22_X1 port map( A1 => n25028, A2 => n24463, B1 => n25022, B2 => 
                           n18274, ZN => n23755);
   U21173 : OAI221_X1 port map( B1 => n21150, B2 => n25040, C1 => n20386, C2 =>
                           n25034, A => n23737, ZN => n23734);
   U21174 : AOI22_X1 port map( A1 => n25028, A2 => n24465, B1 => n25022, B2 => 
                           n18253, ZN => n23737);
   U21175 : OAI221_X1 port map( B1 => n21161, B2 => n25238, C1 => n20397, C2 =>
                           n25232, A => n22750, ZN => n22746);
   U21176 : AOI22_X1 port map( A1 => n25226, A2 => n24443, B1 => n25220, B2 => 
                           n18484, ZN => n22750);
   U21177 : OAI221_X1 port map( B1 => n21160, B2 => n25238, C1 => n20396, C2 =>
                           n25232, A => n22720, ZN => n22717);
   U21178 : AOI22_X1 port map( A1 => n25226, A2 => n24445, B1 => n25220, B2 => 
                           n18463, ZN => n22720);
   U21179 : OAI221_X1 port map( B1 => n21159, B2 => n25238, C1 => n20395, C2 =>
                           n25232, A => n22702, ZN => n22699);
   U21180 : AOI22_X1 port map( A1 => n25226, A2 => n24447, B1 => n25220, B2 => 
                           n18442, ZN => n22702);
   U21181 : OAI221_X1 port map( B1 => n21158, B2 => n25238, C1 => n20394, C2 =>
                           n25232, A => n22684, ZN => n22681);
   U21182 : AOI22_X1 port map( A1 => n25226, A2 => n24449, B1 => n25220, B2 => 
                           n18421, ZN => n22684);
   U21183 : OAI221_X1 port map( B1 => n21157, B2 => n25238, C1 => n20393, C2 =>
                           n25232, A => n22666, ZN => n22663);
   U21184 : AOI22_X1 port map( A1 => n25226, A2 => n24451, B1 => n25220, B2 => 
                           n18400, ZN => n22666);
   U21185 : OAI221_X1 port map( B1 => n21156, B2 => n25238, C1 => n20392, C2 =>
                           n25232, A => n22648, ZN => n22645);
   U21186 : AOI22_X1 port map( A1 => n25226, A2 => n24453, B1 => n25220, B2 => 
                           n18379, ZN => n22648);
   U21187 : OAI221_X1 port map( B1 => n21155, B2 => n25238, C1 => n20391, C2 =>
                           n25232, A => n22630, ZN => n22627);
   U21188 : AOI22_X1 port map( A1 => n25226, A2 => n24455, B1 => n25220, B2 => 
                           n18358, ZN => n22630);
   U21189 : OAI221_X1 port map( B1 => n21154, B2 => n25238, C1 => n20390, C2 =>
                           n25232, A => n22612, ZN => n22609);
   U21190 : AOI22_X1 port map( A1 => n25226, A2 => n24457, B1 => n25220, B2 => 
                           n18337, ZN => n22612);
   U21191 : OAI221_X1 port map( B1 => n21153, B2 => n25238, C1 => n20389, C2 =>
                           n25232, A => n22594, ZN => n22591);
   U21192 : AOI22_X1 port map( A1 => n25226, A2 => n24459, B1 => n25220, B2 => 
                           n18316, ZN => n22594);
   U21193 : OAI221_X1 port map( B1 => n21152, B2 => n25238, C1 => n20388, C2 =>
                           n25232, A => n22576, ZN => n22573);
   U21194 : AOI22_X1 port map( A1 => n25226, A2 => n24461, B1 => n25220, B2 => 
                           n18295, ZN => n22576);
   U21195 : OAI221_X1 port map( B1 => n21151, B2 => n25238, C1 => n20387, C2 =>
                           n25232, A => n22558, ZN => n22555);
   U21196 : AOI22_X1 port map( A1 => n25226, A2 => n24463, B1 => n25220, B2 => 
                           n18274, ZN => n22558);
   U21197 : OAI221_X1 port map( B1 => n21150, B2 => n25238, C1 => n20386, C2 =>
                           n25232, A => n22540, ZN => n22537);
   U21198 : AOI22_X1 port map( A1 => n25226, A2 => n24465, B1 => n25220, B2 => 
                           n18253, ZN => n22540);
   U21199 : OAI221_X1 port map( B1 => n21401, B2 => n25017, C1 => n20321, C2 =>
                           n25011, A => n23720, ZN => n23715);
   U21200 : AOI22_X1 port map( A1 => n25005, A2 => n24626, B1 => n24999, B2 => 
                           n18234, ZN => n23720);
   U21201 : OAI221_X1 port map( B1 => n21400, B2 => n25017, C1 => n20320, C2 =>
                           n25011, A => n23702, ZN => n23697);
   U21202 : AOI22_X1 port map( A1 => n25005, A2 => n24627, B1 => n24999, B2 => 
                           n18213, ZN => n23702);
   U21203 : OAI221_X1 port map( B1 => n21399, B2 => n25017, C1 => n20319, C2 =>
                           n25011, A => n23684, ZN => n23679);
   U21204 : AOI22_X1 port map( A1 => n25005, A2 => n24628, B1 => n24999, B2 => 
                           n18192, ZN => n23684);
   U21205 : OAI221_X1 port map( B1 => n21398, B2 => n25017, C1 => n20318, C2 =>
                           n25011, A => n23666, ZN => n23661);
   U21206 : AOI22_X1 port map( A1 => n25005, A2 => n24629, B1 => n24999, B2 => 
                           n18171, ZN => n23666);
   U21207 : OAI221_X1 port map( B1 => n21397, B2 => n25017, C1 => n20317, C2 =>
                           n25011, A => n23648, ZN => n23643);
   U21208 : AOI22_X1 port map( A1 => n25005, A2 => n24630, B1 => n24999, B2 => 
                           n18150, ZN => n23648);
   U21209 : OAI221_X1 port map( B1 => n21396, B2 => n25017, C1 => n20316, C2 =>
                           n25011, A => n23630, ZN => n23625);
   U21210 : AOI22_X1 port map( A1 => n25005, A2 => n24631, B1 => n24999, B2 => 
                           n18129, ZN => n23630);
   U21211 : OAI221_X1 port map( B1 => n21395, B2 => n25017, C1 => n20315, C2 =>
                           n25011, A => n23612, ZN => n23607);
   U21212 : AOI22_X1 port map( A1 => n25005, A2 => n24632, B1 => n24999, B2 => 
                           n18108, ZN => n23612);
   U21213 : OAI221_X1 port map( B1 => n21394, B2 => n25017, C1 => n20314, C2 =>
                           n25011, A => n23594, ZN => n23589);
   U21214 : AOI22_X1 port map( A1 => n25005, A2 => n24633, B1 => n24999, B2 => 
                           n18087, ZN => n23594);
   U21215 : OAI221_X1 port map( B1 => n21393, B2 => n25017, C1 => n20313, C2 =>
                           n25011, A => n23576, ZN => n23571);
   U21216 : AOI22_X1 port map( A1 => n25005, A2 => n24634, B1 => n24999, B2 => 
                           n18066, ZN => n23576);
   U21217 : OAI221_X1 port map( B1 => n21392, B2 => n25017, C1 => n20312, C2 =>
                           n25011, A => n23558, ZN => n23553);
   U21218 : AOI22_X1 port map( A1 => n25005, A2 => n24635, B1 => n24999, B2 => 
                           n18045, ZN => n23558);
   U21219 : OAI221_X1 port map( B1 => n21391, B2 => n25017, C1 => n20311, C2 =>
                           n25011, A => n23540, ZN => n23535);
   U21220 : AOI22_X1 port map( A1 => n25005, A2 => n24636, B1 => n24999, B2 => 
                           n18024, ZN => n23540);
   U21221 : OAI221_X1 port map( B1 => n21390, B2 => n25017, C1 => n20310, C2 =>
                           n25011, A => n23522, ZN => n23517);
   U21222 : AOI22_X1 port map( A1 => n25005, A2 => n24637, B1 => n24999, B2 => 
                           n18003, ZN => n23522);
   U21223 : OAI221_X1 port map( B1 => n21389, B2 => n25018, C1 => n20309, C2 =>
                           n25012, A => n23504, ZN => n23499);
   U21224 : AOI22_X1 port map( A1 => n25006, A2 => n24638, B1 => n25000, B2 => 
                           n17982, ZN => n23504);
   U21225 : OAI221_X1 port map( B1 => n21388, B2 => n25018, C1 => n20308, C2 =>
                           n25012, A => n23486, ZN => n23481);
   U21226 : AOI22_X1 port map( A1 => n25006, A2 => n24639, B1 => n25000, B2 => 
                           n17961, ZN => n23486);
   U21227 : OAI221_X1 port map( B1 => n21387, B2 => n25018, C1 => n20307, C2 =>
                           n25012, A => n23468, ZN => n23463);
   U21228 : AOI22_X1 port map( A1 => n25006, A2 => n24640, B1 => n25000, B2 => 
                           n17940, ZN => n23468);
   U21229 : OAI221_X1 port map( B1 => n21386, B2 => n25018, C1 => n20306, C2 =>
                           n25012, A => n23450, ZN => n23445);
   U21230 : AOI22_X1 port map( A1 => n25006, A2 => n24641, B1 => n25000, B2 => 
                           n17919, ZN => n23450);
   U21231 : OAI221_X1 port map( B1 => n21385, B2 => n25018, C1 => n20305, C2 =>
                           n25012, A => n23432, ZN => n23427);
   U21232 : AOI22_X1 port map( A1 => n25006, A2 => n24642, B1 => n25000, B2 => 
                           n17898, ZN => n23432);
   U21233 : OAI221_X1 port map( B1 => n21384, B2 => n25018, C1 => n20304, C2 =>
                           n25012, A => n23414, ZN => n23409);
   U21234 : AOI22_X1 port map( A1 => n25006, A2 => n24643, B1 => n25000, B2 => 
                           n17877, ZN => n23414);
   U21235 : OAI221_X1 port map( B1 => n21383, B2 => n25018, C1 => n20303, C2 =>
                           n25012, A => n23396, ZN => n23391);
   U21236 : AOI22_X1 port map( A1 => n25006, A2 => n24644, B1 => n25000, B2 => 
                           n17856, ZN => n23396);
   U21237 : OAI221_X1 port map( B1 => n21382, B2 => n25018, C1 => n20302, C2 =>
                           n25012, A => n23378, ZN => n23373);
   U21238 : AOI22_X1 port map( A1 => n25006, A2 => n24645, B1 => n25000, B2 => 
                           n17835, ZN => n23378);
   U21239 : OAI221_X1 port map( B1 => n21381, B2 => n25018, C1 => n20301, C2 =>
                           n25012, A => n23360, ZN => n23355);
   U21240 : AOI22_X1 port map( A1 => n25006, A2 => n24646, B1 => n25000, B2 => 
                           n17814, ZN => n23360);
   U21241 : OAI221_X1 port map( B1 => n21380, B2 => n25018, C1 => n20300, C2 =>
                           n25012, A => n23342, ZN => n23337);
   U21242 : AOI22_X1 port map( A1 => n25006, A2 => n24647, B1 => n25000, B2 => 
                           n17793, ZN => n23342);
   U21243 : OAI221_X1 port map( B1 => n21379, B2 => n25018, C1 => n20299, C2 =>
                           n25012, A => n23324, ZN => n23319);
   U21244 : AOI22_X1 port map( A1 => n25006, A2 => n24648, B1 => n25000, B2 => 
                           n17772, ZN => n23324);
   U21245 : OAI221_X1 port map( B1 => n21378, B2 => n25018, C1 => n20298, C2 =>
                           n25012, A => n23306, ZN => n23301);
   U21246 : AOI22_X1 port map( A1 => n25006, A2 => n24649, B1 => n25000, B2 => 
                           n17751, ZN => n23306);
   U21247 : OAI221_X1 port map( B1 => n21377, B2 => n25019, C1 => n20297, C2 =>
                           n25013, A => n23288, ZN => n23283);
   U21248 : AOI22_X1 port map( A1 => n25007, A2 => n24650, B1 => n25001, B2 => 
                           n17730, ZN => n23288);
   U21249 : OAI221_X1 port map( B1 => n21376, B2 => n25019, C1 => n20296, C2 =>
                           n25013, A => n23270, ZN => n23265);
   U21250 : AOI22_X1 port map( A1 => n25007, A2 => n24651, B1 => n25001, B2 => 
                           n17709, ZN => n23270);
   U21251 : OAI221_X1 port map( B1 => n21375, B2 => n25019, C1 => n20295, C2 =>
                           n25013, A => n23252, ZN => n23247);
   U21252 : AOI22_X1 port map( A1 => n25007, A2 => n24652, B1 => n25001, B2 => 
                           n17688, ZN => n23252);
   U21253 : OAI221_X1 port map( B1 => n21374, B2 => n25019, C1 => n20294, C2 =>
                           n25013, A => n23234, ZN => n23229);
   U21254 : AOI22_X1 port map( A1 => n25007, A2 => n24653, B1 => n25001, B2 => 
                           n17667, ZN => n23234);
   U21255 : OAI221_X1 port map( B1 => n21373, B2 => n25019, C1 => n20293, C2 =>
                           n25013, A => n23216, ZN => n23211);
   U21256 : AOI22_X1 port map( A1 => n25007, A2 => n24654, B1 => n25001, B2 => 
                           n17646, ZN => n23216);
   U21257 : OAI221_X1 port map( B1 => n21372, B2 => n25019, C1 => n20292, C2 =>
                           n25013, A => n23198, ZN => n23193);
   U21258 : AOI22_X1 port map( A1 => n25007, A2 => n24655, B1 => n25001, B2 => 
                           n17625, ZN => n23198);
   U21259 : OAI221_X1 port map( B1 => n21371, B2 => n25019, C1 => n20291, C2 =>
                           n25013, A => n23180, ZN => n23175);
   U21260 : AOI22_X1 port map( A1 => n25007, A2 => n24656, B1 => n25001, B2 => 
                           n17604, ZN => n23180);
   U21261 : OAI221_X1 port map( B1 => n21370, B2 => n25019, C1 => n20290, C2 =>
                           n25013, A => n23162, ZN => n23157);
   U21262 : AOI22_X1 port map( A1 => n25007, A2 => n24657, B1 => n25001, B2 => 
                           n17583, ZN => n23162);
   U21263 : OAI221_X1 port map( B1 => n21369, B2 => n25019, C1 => n20289, C2 =>
                           n25013, A => n23144, ZN => n23139);
   U21264 : AOI22_X1 port map( A1 => n25007, A2 => n24658, B1 => n25001, B2 => 
                           n17562, ZN => n23144);
   U21265 : OAI221_X1 port map( B1 => n21368, B2 => n25019, C1 => n20288, C2 =>
                           n25013, A => n23126, ZN => n23121);
   U21266 : AOI22_X1 port map( A1 => n25007, A2 => n24659, B1 => n25001, B2 => 
                           n17541, ZN => n23126);
   U21267 : OAI221_X1 port map( B1 => n21367, B2 => n25019, C1 => n20287, C2 =>
                           n25013, A => n23108, ZN => n23103);
   U21268 : AOI22_X1 port map( A1 => n25007, A2 => n24660, B1 => n25001, B2 => 
                           n17520, ZN => n23108);
   U21269 : OAI221_X1 port map( B1 => n21366, B2 => n25019, C1 => n20286, C2 =>
                           n25013, A => n23090, ZN => n23085);
   U21270 : AOI22_X1 port map( A1 => n25007, A2 => n24661, B1 => n25001, B2 => 
                           n17499, ZN => n23090);
   U21271 : OAI221_X1 port map( B1 => n21365, B2 => n25020, C1 => n20285, C2 =>
                           n25014, A => n23072, ZN => n23067);
   U21272 : AOI22_X1 port map( A1 => n25008, A2 => n24662, B1 => n25002, B2 => 
                           n17478, ZN => n23072);
   U21273 : OAI221_X1 port map( B1 => n21364, B2 => n25020, C1 => n20284, C2 =>
                           n25014, A => n23054, ZN => n23049);
   U21274 : AOI22_X1 port map( A1 => n25008, A2 => n24663, B1 => n25002, B2 => 
                           n17457, ZN => n23054);
   U21275 : OAI221_X1 port map( B1 => n21363, B2 => n25020, C1 => n20283, C2 =>
                           n25014, A => n23036, ZN => n23031);
   U21276 : AOI22_X1 port map( A1 => n25008, A2 => n24664, B1 => n25002, B2 => 
                           n17436, ZN => n23036);
   U21277 : OAI221_X1 port map( B1 => n21362, B2 => n25020, C1 => n20282, C2 =>
                           n25014, A => n23018, ZN => n23013);
   U21278 : AOI22_X1 port map( A1 => n25008, A2 => n24665, B1 => n25002, B2 => 
                           n17415, ZN => n23018);
   U21279 : OAI221_X1 port map( B1 => n21361, B2 => n25020, C1 => n20281, C2 =>
                           n25014, A => n23000, ZN => n22995);
   U21280 : AOI22_X1 port map( A1 => n25008, A2 => n24666, B1 => n25002, B2 => 
                           n17394, ZN => n23000);
   U21281 : OAI221_X1 port map( B1 => n21360, B2 => n25020, C1 => n20280, C2 =>
                           n25014, A => n22982, ZN => n22977);
   U21282 : AOI22_X1 port map( A1 => n25008, A2 => n24667, B1 => n25002, B2 => 
                           n17373, ZN => n22982);
   U21283 : OAI221_X1 port map( B1 => n21359, B2 => n25020, C1 => n20279, C2 =>
                           n25014, A => n22964, ZN => n22959);
   U21284 : AOI22_X1 port map( A1 => n25008, A2 => n24668, B1 => n25002, B2 => 
                           n17352, ZN => n22964);
   U21285 : OAI221_X1 port map( B1 => n21358, B2 => n25020, C1 => n20278, C2 =>
                           n25014, A => n22946, ZN => n22941);
   U21286 : AOI22_X1 port map( A1 => n25008, A2 => n24669, B1 => n25002, B2 => 
                           n17331, ZN => n22946);
   U21287 : OAI221_X1 port map( B1 => n21357, B2 => n25020, C1 => n20277, C2 =>
                           n25014, A => n22928, ZN => n22923);
   U21288 : AOI22_X1 port map( A1 => n25008, A2 => n24670, B1 => n25002, B2 => 
                           n17310, ZN => n22928);
   U21289 : OAI221_X1 port map( B1 => n21356, B2 => n25020, C1 => n20276, C2 =>
                           n25014, A => n22910, ZN => n22905);
   U21290 : AOI22_X1 port map( A1 => n25008, A2 => n24671, B1 => n25002, B2 => 
                           n17289, ZN => n22910);
   U21291 : OAI221_X1 port map( B1 => n21355, B2 => n25020, C1 => n20275, C2 =>
                           n25014, A => n22892, ZN => n22887);
   U21292 : AOI22_X1 port map( A1 => n25008, A2 => n24672, B1 => n25002, B2 => 
                           n17268, ZN => n22892);
   U21293 : OAI221_X1 port map( B1 => n21354, B2 => n25020, C1 => n20274, C2 =>
                           n25014, A => n22874, ZN => n22869);
   U21294 : AOI22_X1 port map( A1 => n25008, A2 => n24673, B1 => n25002, B2 => 
                           n17247, ZN => n22874);
   U21295 : OAI221_X1 port map( B1 => n21401, B2 => n25215, C1 => n20321, C2 =>
                           n25209, A => n22523, ZN => n22518);
   U21296 : AOI22_X1 port map( A1 => n25203, A2 => n24626, B1 => n25197, B2 => 
                           n18234, ZN => n22523);
   U21297 : OAI221_X1 port map( B1 => n21400, B2 => n25215, C1 => n20320, C2 =>
                           n25209, A => n22505, ZN => n22500);
   U21298 : AOI22_X1 port map( A1 => n25203, A2 => n24627, B1 => n25197, B2 => 
                           n18213, ZN => n22505);
   U21299 : OAI221_X1 port map( B1 => n21399, B2 => n25215, C1 => n20319, C2 =>
                           n25209, A => n22487, ZN => n22482);
   U21300 : AOI22_X1 port map( A1 => n25203, A2 => n24628, B1 => n25197, B2 => 
                           n18192, ZN => n22487);
   U21301 : OAI221_X1 port map( B1 => n21398, B2 => n25215, C1 => n20318, C2 =>
                           n25209, A => n22469, ZN => n22464);
   U21302 : AOI22_X1 port map( A1 => n25203, A2 => n24629, B1 => n25197, B2 => 
                           n18171, ZN => n22469);
   U21303 : OAI221_X1 port map( B1 => n21397, B2 => n25215, C1 => n20317, C2 =>
                           n25209, A => n22451, ZN => n22446);
   U21304 : AOI22_X1 port map( A1 => n25203, A2 => n24630, B1 => n25197, B2 => 
                           n18150, ZN => n22451);
   U21305 : OAI221_X1 port map( B1 => n21396, B2 => n25215, C1 => n20316, C2 =>
                           n25209, A => n22433, ZN => n22428);
   U21306 : AOI22_X1 port map( A1 => n25203, A2 => n24631, B1 => n25197, B2 => 
                           n18129, ZN => n22433);
   U21307 : OAI221_X1 port map( B1 => n21395, B2 => n25215, C1 => n20315, C2 =>
                           n25209, A => n22415, ZN => n22410);
   U21308 : AOI22_X1 port map( A1 => n25203, A2 => n24632, B1 => n25197, B2 => 
                           n18108, ZN => n22415);
   U21309 : OAI221_X1 port map( B1 => n21394, B2 => n25215, C1 => n20314, C2 =>
                           n25209, A => n22397, ZN => n22392);
   U21310 : AOI22_X1 port map( A1 => n25203, A2 => n24633, B1 => n25197, B2 => 
                           n18087, ZN => n22397);
   U21311 : OAI221_X1 port map( B1 => n21393, B2 => n25215, C1 => n20313, C2 =>
                           n25209, A => n22379, ZN => n22374);
   U21312 : AOI22_X1 port map( A1 => n25203, A2 => n24634, B1 => n25197, B2 => 
                           n18066, ZN => n22379);
   U21313 : OAI221_X1 port map( B1 => n21392, B2 => n25215, C1 => n20312, C2 =>
                           n25209, A => n22361, ZN => n22356);
   U21314 : AOI22_X1 port map( A1 => n25203, A2 => n24635, B1 => n25197, B2 => 
                           n18045, ZN => n22361);
   U21315 : OAI221_X1 port map( B1 => n21391, B2 => n25215, C1 => n20311, C2 =>
                           n25209, A => n22343, ZN => n22338);
   U21316 : AOI22_X1 port map( A1 => n25203, A2 => n24636, B1 => n25197, B2 => 
                           n18024, ZN => n22343);
   U21317 : OAI221_X1 port map( B1 => n21390, B2 => n25215, C1 => n20310, C2 =>
                           n25209, A => n22325, ZN => n22320);
   U21318 : AOI22_X1 port map( A1 => n25203, A2 => n24637, B1 => n25197, B2 => 
                           n18003, ZN => n22325);
   U21319 : OAI221_X1 port map( B1 => n21389, B2 => n25216, C1 => n20309, C2 =>
                           n25210, A => n22307, ZN => n22302);
   U21320 : AOI22_X1 port map( A1 => n25204, A2 => n24638, B1 => n25198, B2 => 
                           n17982, ZN => n22307);
   U21321 : OAI221_X1 port map( B1 => n21388, B2 => n25216, C1 => n20308, C2 =>
                           n25210, A => n22289, ZN => n22284);
   U21322 : AOI22_X1 port map( A1 => n25204, A2 => n24639, B1 => n25198, B2 => 
                           n17961, ZN => n22289);
   U21323 : OAI221_X1 port map( B1 => n21387, B2 => n25216, C1 => n20307, C2 =>
                           n25210, A => n22271, ZN => n22266);
   U21324 : AOI22_X1 port map( A1 => n25204, A2 => n24640, B1 => n25198, B2 => 
                           n17940, ZN => n22271);
   U21325 : OAI221_X1 port map( B1 => n21386, B2 => n25216, C1 => n20306, C2 =>
                           n25210, A => n22253, ZN => n22248);
   U21326 : AOI22_X1 port map( A1 => n25204, A2 => n24641, B1 => n25198, B2 => 
                           n17919, ZN => n22253);
   U21327 : OAI221_X1 port map( B1 => n21385, B2 => n25216, C1 => n20305, C2 =>
                           n25210, A => n22235, ZN => n22230);
   U21328 : AOI22_X1 port map( A1 => n25204, A2 => n24642, B1 => n25198, B2 => 
                           n17898, ZN => n22235);
   U21329 : OAI221_X1 port map( B1 => n21384, B2 => n25216, C1 => n20304, C2 =>
                           n25210, A => n22217, ZN => n22212);
   U21330 : AOI22_X1 port map( A1 => n25204, A2 => n24643, B1 => n25198, B2 => 
                           n17877, ZN => n22217);
   U21331 : OAI221_X1 port map( B1 => n21383, B2 => n25216, C1 => n20303, C2 =>
                           n25210, A => n22199, ZN => n22194);
   U21332 : AOI22_X1 port map( A1 => n25204, A2 => n24644, B1 => n25198, B2 => 
                           n17856, ZN => n22199);
   U21333 : OAI221_X1 port map( B1 => n21382, B2 => n25216, C1 => n20302, C2 =>
                           n25210, A => n22181, ZN => n22176);
   U21334 : AOI22_X1 port map( A1 => n25204, A2 => n24645, B1 => n25198, B2 => 
                           n17835, ZN => n22181);
   U21335 : OAI221_X1 port map( B1 => n21381, B2 => n25216, C1 => n20301, C2 =>
                           n25210, A => n22163, ZN => n22158);
   U21336 : AOI22_X1 port map( A1 => n25204, A2 => n24646, B1 => n25198, B2 => 
                           n17814, ZN => n22163);
   U21337 : OAI221_X1 port map( B1 => n21380, B2 => n25216, C1 => n20300, C2 =>
                           n25210, A => n22145, ZN => n22140);
   U21338 : AOI22_X1 port map( A1 => n25204, A2 => n24647, B1 => n25198, B2 => 
                           n17793, ZN => n22145);
   U21339 : OAI221_X1 port map( B1 => n21379, B2 => n25216, C1 => n20299, C2 =>
                           n25210, A => n22127, ZN => n22122);
   U21340 : AOI22_X1 port map( A1 => n25204, A2 => n24648, B1 => n25198, B2 => 
                           n17772, ZN => n22127);
   U21341 : OAI221_X1 port map( B1 => n21378, B2 => n25216, C1 => n20298, C2 =>
                           n25210, A => n22109, ZN => n22104);
   U21342 : AOI22_X1 port map( A1 => n25204, A2 => n24649, B1 => n25198, B2 => 
                           n17751, ZN => n22109);
   U21343 : OAI221_X1 port map( B1 => n21377, B2 => n25217, C1 => n20297, C2 =>
                           n25211, A => n22091, ZN => n22086);
   U21344 : AOI22_X1 port map( A1 => n25205, A2 => n24650, B1 => n25199, B2 => 
                           n17730, ZN => n22091);
   U21345 : OAI221_X1 port map( B1 => n21376, B2 => n25217, C1 => n20296, C2 =>
                           n25211, A => n22073, ZN => n22068);
   U21346 : AOI22_X1 port map( A1 => n25205, A2 => n24651, B1 => n25199, B2 => 
                           n17709, ZN => n22073);
   U21347 : OAI221_X1 port map( B1 => n21375, B2 => n25217, C1 => n20295, C2 =>
                           n25211, A => n22055, ZN => n22050);
   U21348 : AOI22_X1 port map( A1 => n25205, A2 => n24652, B1 => n25199, B2 => 
                           n17688, ZN => n22055);
   U21349 : OAI221_X1 port map( B1 => n21374, B2 => n25217, C1 => n20294, C2 =>
                           n25211, A => n22037, ZN => n22032);
   U21350 : AOI22_X1 port map( A1 => n25205, A2 => n24653, B1 => n25199, B2 => 
                           n17667, ZN => n22037);
   U21351 : OAI221_X1 port map( B1 => n21373, B2 => n25217, C1 => n20293, C2 =>
                           n25211, A => n22019, ZN => n22014);
   U21352 : AOI22_X1 port map( A1 => n25205, A2 => n24654, B1 => n25199, B2 => 
                           n17646, ZN => n22019);
   U21353 : OAI221_X1 port map( B1 => n21372, B2 => n25217, C1 => n20292, C2 =>
                           n25211, A => n22001, ZN => n21996);
   U21354 : AOI22_X1 port map( A1 => n25205, A2 => n24655, B1 => n25199, B2 => 
                           n17625, ZN => n22001);
   U21355 : OAI221_X1 port map( B1 => n21371, B2 => n25217, C1 => n20291, C2 =>
                           n25211, A => n21983, ZN => n21978);
   U21356 : AOI22_X1 port map( A1 => n25205, A2 => n24656, B1 => n25199, B2 => 
                           n17604, ZN => n21983);
   U21357 : OAI221_X1 port map( B1 => n21370, B2 => n25217, C1 => n20290, C2 =>
                           n25211, A => n21965, ZN => n21960);
   U21358 : AOI22_X1 port map( A1 => n25205, A2 => n24657, B1 => n25199, B2 => 
                           n17583, ZN => n21965);
   U21359 : OAI221_X1 port map( B1 => n21369, B2 => n25217, C1 => n20289, C2 =>
                           n25211, A => n21947, ZN => n21942);
   U21360 : AOI22_X1 port map( A1 => n25205, A2 => n24658, B1 => n25199, B2 => 
                           n17562, ZN => n21947);
   U21361 : OAI221_X1 port map( B1 => n21368, B2 => n25217, C1 => n20288, C2 =>
                           n25211, A => n21929, ZN => n21924);
   U21362 : AOI22_X1 port map( A1 => n25205, A2 => n24659, B1 => n25199, B2 => 
                           n17541, ZN => n21929);
   U21363 : OAI221_X1 port map( B1 => n21367, B2 => n25217, C1 => n20287, C2 =>
                           n25211, A => n21911, ZN => n21906);
   U21364 : AOI22_X1 port map( A1 => n25205, A2 => n24660, B1 => n25199, B2 => 
                           n17520, ZN => n21911);
   U21365 : OAI221_X1 port map( B1 => n21366, B2 => n25217, C1 => n20286, C2 =>
                           n25211, A => n21893, ZN => n21888);
   U21366 : AOI22_X1 port map( A1 => n25205, A2 => n24661, B1 => n25199, B2 => 
                           n17499, ZN => n21893);
   U21367 : OAI221_X1 port map( B1 => n21365, B2 => n25218, C1 => n20285, C2 =>
                           n25212, A => n21875, ZN => n21870);
   U21368 : AOI22_X1 port map( A1 => n25206, A2 => n24662, B1 => n25200, B2 => 
                           n17478, ZN => n21875);
   U21369 : OAI221_X1 port map( B1 => n21364, B2 => n25218, C1 => n20284, C2 =>
                           n25212, A => n21857, ZN => n21852);
   U21370 : AOI22_X1 port map( A1 => n25206, A2 => n24663, B1 => n25200, B2 => 
                           n17457, ZN => n21857);
   U21371 : OAI221_X1 port map( B1 => n21363, B2 => n25218, C1 => n20283, C2 =>
                           n25212, A => n21839, ZN => n21834);
   U21372 : AOI22_X1 port map( A1 => n25206, A2 => n24664, B1 => n25200, B2 => 
                           n17436, ZN => n21839);
   U21373 : OAI221_X1 port map( B1 => n21362, B2 => n25218, C1 => n20282, C2 =>
                           n25212, A => n21821, ZN => n21816);
   U21374 : AOI22_X1 port map( A1 => n25206, A2 => n24665, B1 => n25200, B2 => 
                           n17415, ZN => n21821);
   U21375 : OAI221_X1 port map( B1 => n21361, B2 => n25218, C1 => n20281, C2 =>
                           n25212, A => n21803, ZN => n21798);
   U21376 : AOI22_X1 port map( A1 => n25206, A2 => n24666, B1 => n25200, B2 => 
                           n17394, ZN => n21803);
   U21377 : OAI221_X1 port map( B1 => n21360, B2 => n25218, C1 => n20280, C2 =>
                           n25212, A => n21785, ZN => n21780);
   U21378 : AOI22_X1 port map( A1 => n25206, A2 => n24667, B1 => n25200, B2 => 
                           n17373, ZN => n21785);
   U21379 : OAI221_X1 port map( B1 => n21359, B2 => n25218, C1 => n20279, C2 =>
                           n25212, A => n21767, ZN => n21762);
   U21380 : AOI22_X1 port map( A1 => n25206, A2 => n24668, B1 => n25200, B2 => 
                           n17352, ZN => n21767);
   U21381 : OAI221_X1 port map( B1 => n21358, B2 => n25218, C1 => n20278, C2 =>
                           n25212, A => n21749, ZN => n21744);
   U21382 : AOI22_X1 port map( A1 => n25206, A2 => n24669, B1 => n25200, B2 => 
                           n17331, ZN => n21749);
   U21383 : OAI221_X1 port map( B1 => n21357, B2 => n25218, C1 => n20277, C2 =>
                           n25212, A => n21731, ZN => n21726);
   U21384 : AOI22_X1 port map( A1 => n25206, A2 => n24670, B1 => n25200, B2 => 
                           n17310, ZN => n21731);
   U21385 : OAI221_X1 port map( B1 => n21356, B2 => n25218, C1 => n20276, C2 =>
                           n25212, A => n21713, ZN => n21708);
   U21386 : AOI22_X1 port map( A1 => n25206, A2 => n24671, B1 => n25200, B2 => 
                           n17289, ZN => n21713);
   U21387 : OAI221_X1 port map( B1 => n21355, B2 => n25218, C1 => n20275, C2 =>
                           n25212, A => n21695, ZN => n21690);
   U21388 : AOI22_X1 port map( A1 => n25206, A2 => n24672, B1 => n25200, B2 => 
                           n17268, ZN => n21695);
   U21389 : OAI221_X1 port map( B1 => n21354, B2 => n25218, C1 => n20274, C2 =>
                           n25212, A => n21677, ZN => n21672);
   U21390 : AOI22_X1 port map( A1 => n25206, A2 => n24673, B1 => n25200, B2 => 
                           n17247, ZN => n21677);
   U21391 : OAI221_X1 port map( B1 => n21222, B2 => n25123, C1 => n19558, C2 =>
                           n25117, A => n22771, ZN => n22756);
   U21392 : AOI22_X1 port map( A1 => n25111, A2 => n24481, B1 => n25105, B2 => 
                           n20005, ZN => n22771);
   U21393 : OAI221_X1 port map( B1 => n21350, B2 => n25021, C1 => n20270, C2 =>
                           n25015, A => n22796, ZN => n22781);
   U21394 : AOI22_X1 port map( A1 => n25009, A2 => n24613, B1 => n25003, B2 => 
                           n17163, ZN => n22796);
   U21395 : OAI221_X1 port map( B1 => n21225, B2 => n25123, C1 => n19561, C2 =>
                           n25117, A => n22848, ZN => n22843);
   U21396 : AOI22_X1 port map( A1 => n25111, A2 => n24478, B1 => n25105, B2 => 
                           n20008, ZN => n22848);
   U21397 : OAI221_X1 port map( B1 => n21353, B2 => n25021, C1 => n20273, C2 =>
                           n25015, A => n22856, ZN => n22851);
   U21398 : AOI22_X1 port map( A1 => n25009, A2 => n24607, B1 => n25003, B2 => 
                           n17226, ZN => n22856);
   U21399 : OAI221_X1 port map( B1 => n21224, B2 => n25123, C1 => n19560, C2 =>
                           n25117, A => n22830, ZN => n22825);
   U21400 : AOI22_X1 port map( A1 => n25111, A2 => n24479, B1 => n25105, B2 => 
                           n20007, ZN => n22830);
   U21401 : OAI221_X1 port map( B1 => n21352, B2 => n25021, C1 => n20272, C2 =>
                           n25015, A => n22838, ZN => n22833);
   U21402 : AOI22_X1 port map( A1 => n25009, A2 => n24609, B1 => n25003, B2 => 
                           n17205, ZN => n22838);
   U21403 : OAI221_X1 port map( B1 => n21223, B2 => n25123, C1 => n19559, C2 =>
                           n25117, A => n22812, ZN => n22807);
   U21404 : AOI22_X1 port map( A1 => n25111, A2 => n24480, B1 => n25105, B2 => 
                           n20006, ZN => n22812);
   U21405 : OAI221_X1 port map( B1 => n21351, B2 => n25021, C1 => n20271, C2 =>
                           n25015, A => n22820, ZN => n22815);
   U21406 : AOI22_X1 port map( A1 => n25009, A2 => n24611, B1 => n25003, B2 => 
                           n17184, ZN => n22820);
   U21407 : OAI221_X1 port map( B1 => n21225, B2 => n25321, C1 => n19561, C2 =>
                           n25315, A => n21651, ZN => n21646);
   U21408 : AOI22_X1 port map( A1 => n25309, A2 => n24478, B1 => n25303, B2 => 
                           n20008, ZN => n21651);
   U21409 : OAI221_X1 port map( B1 => n21353, B2 => n25219, C1 => n20273, C2 =>
                           n25213, A => n21659, ZN => n21654);
   U21410 : AOI22_X1 port map( A1 => n25207, A2 => n24607, B1 => n25201, B2 => 
                           n17226, ZN => n21659);
   U21411 : OAI221_X1 port map( B1 => n21224, B2 => n25321, C1 => n19560, C2 =>
                           n25315, A => n21633, ZN => n21628);
   U21412 : AOI22_X1 port map( A1 => n25309, A2 => n24479, B1 => n25303, B2 => 
                           n20007, ZN => n21633);
   U21413 : OAI221_X1 port map( B1 => n21352, B2 => n25219, C1 => n20272, C2 =>
                           n25213, A => n21641, ZN => n21636);
   U21414 : AOI22_X1 port map( A1 => n25207, A2 => n24609, B1 => n25201, B2 => 
                           n17205, ZN => n21641);
   U21415 : OAI221_X1 port map( B1 => n21223, B2 => n25321, C1 => n19559, C2 =>
                           n25315, A => n21615, ZN => n21610);
   U21416 : AOI22_X1 port map( A1 => n25309, A2 => n24480, B1 => n25303, B2 => 
                           n20006, ZN => n21615);
   U21417 : OAI221_X1 port map( B1 => n21351, B2 => n25219, C1 => n20271, C2 =>
                           n25213, A => n21623, ZN => n21618);
   U21418 : AOI22_X1 port map( A1 => n25207, A2 => n24611, B1 => n25201, B2 => 
                           n17184, ZN => n21623);
   U21419 : OAI221_X1 port map( B1 => n21222, B2 => n25321, C1 => n19558, C2 =>
                           n25315, A => n21574, ZN => n21559);
   U21420 : AOI22_X1 port map( A1 => n25309, A2 => n24481, B1 => n25303, B2 => 
                           n20005, ZN => n21574);
   U21421 : OAI221_X1 port map( B1 => n21350, B2 => n25219, C1 => n20270, C2 =>
                           n25213, A => n21599, ZN => n21584);
   U21422 : AOI22_X1 port map( A1 => n25207, A2 => n24613, B1 => n25201, B2 => 
                           n17163, ZN => n21599);
   U21423 : OAI221_X1 port map( B1 => n20697, B2 => n25095, C1 => n21017, C2 =>
                           n25089, A => n23713, ZN => n23706);
   U21424 : AOI222_X1 port map( A1 => n25083, A2 => n24206, B1 => n25077, B2 =>
                           n18228, C1 => n25071, C2 => n18227, ZN => n23713);
   U21425 : OAI221_X1 port map( B1 => n20696, B2 => n25095, C1 => n21016, C2 =>
                           n25089, A => n23695, ZN => n23688);
   U21426 : AOI222_X1 port map( A1 => n25083, A2 => n24208, B1 => n25077, B2 =>
                           n18207, C1 => n25071, C2 => n18206, ZN => n23695);
   U21427 : OAI221_X1 port map( B1 => n20695, B2 => n25095, C1 => n21015, C2 =>
                           n25089, A => n23677, ZN => n23670);
   U21428 : AOI222_X1 port map( A1 => n25083, A2 => n24210, B1 => n25077, B2 =>
                           n18186, C1 => n25071, C2 => n18185, ZN => n23677);
   U21429 : OAI221_X1 port map( B1 => n20694, B2 => n25095, C1 => n21014, C2 =>
                           n25089, A => n23659, ZN => n23652);
   U21430 : AOI222_X1 port map( A1 => n25083, A2 => n24212, B1 => n25077, B2 =>
                           n18165, C1 => n25071, C2 => n18164, ZN => n23659);
   U21431 : OAI221_X1 port map( B1 => n20693, B2 => n25095, C1 => n21013, C2 =>
                           n25089, A => n23641, ZN => n23634);
   U21432 : AOI222_X1 port map( A1 => n25083, A2 => n24214, B1 => n25077, B2 =>
                           n18144, C1 => n25071, C2 => n18143, ZN => n23641);
   U21433 : OAI221_X1 port map( B1 => n20692, B2 => n25095, C1 => n21012, C2 =>
                           n25089, A => n23623, ZN => n23616);
   U21434 : AOI222_X1 port map( A1 => n25083, A2 => n24216, B1 => n25077, B2 =>
                           n18123, C1 => n25071, C2 => n18122, ZN => n23623);
   U21435 : OAI221_X1 port map( B1 => n20691, B2 => n25095, C1 => n21011, C2 =>
                           n25089, A => n23605, ZN => n23598);
   U21436 : AOI222_X1 port map( A1 => n25083, A2 => n24218, B1 => n25077, B2 =>
                           n18102, C1 => n25071, C2 => n18101, ZN => n23605);
   U21437 : OAI221_X1 port map( B1 => n20690, B2 => n25095, C1 => n21010, C2 =>
                           n25089, A => n23587, ZN => n23580);
   U21438 : AOI222_X1 port map( A1 => n25083, A2 => n24220, B1 => n25077, B2 =>
                           n18081, C1 => n25071, C2 => n18080, ZN => n23587);
   U21439 : OAI221_X1 port map( B1 => n20689, B2 => n25095, C1 => n21009, C2 =>
                           n25089, A => n23569, ZN => n23562);
   U21440 : AOI222_X1 port map( A1 => n25083, A2 => n24222, B1 => n25077, B2 =>
                           n18060, C1 => n25071, C2 => n18059, ZN => n23569);
   U21441 : OAI221_X1 port map( B1 => n20688, B2 => n25095, C1 => n21008, C2 =>
                           n25089, A => n23551, ZN => n23544);
   U21442 : AOI222_X1 port map( A1 => n25083, A2 => n24224, B1 => n25077, B2 =>
                           n18039, C1 => n25071, C2 => n18038, ZN => n23551);
   U21443 : OAI221_X1 port map( B1 => n20687, B2 => n25095, C1 => n21007, C2 =>
                           n25089, A => n23533, ZN => n23526);
   U21444 : AOI222_X1 port map( A1 => n25083, A2 => n24226, B1 => n25077, B2 =>
                           n18018, C1 => n25071, C2 => n18017, ZN => n23533);
   U21445 : OAI221_X1 port map( B1 => n20686, B2 => n25095, C1 => n21006, C2 =>
                           n25089, A => n23515, ZN => n23508);
   U21446 : AOI222_X1 port map( A1 => n25083, A2 => n24228, B1 => n25077, B2 =>
                           n17997, C1 => n25071, C2 => n17996, ZN => n23515);
   U21447 : OAI221_X1 port map( B1 => n20685, B2 => n25096, C1 => n21005, C2 =>
                           n25090, A => n23497, ZN => n23490);
   U21448 : AOI222_X1 port map( A1 => n25084, A2 => n24230, B1 => n25078, B2 =>
                           n17976, C1 => n25072, C2 => n17975, ZN => n23497);
   U21449 : OAI221_X1 port map( B1 => n20684, B2 => n25096, C1 => n21004, C2 =>
                           n25090, A => n23479, ZN => n23472);
   U21450 : AOI222_X1 port map( A1 => n25084, A2 => n24232, B1 => n25078, B2 =>
                           n17955, C1 => n25072, C2 => n17954, ZN => n23479);
   U21451 : OAI221_X1 port map( B1 => n20683, B2 => n25096, C1 => n21003, C2 =>
                           n25090, A => n23461, ZN => n23454);
   U21452 : AOI222_X1 port map( A1 => n25084, A2 => n24234, B1 => n25078, B2 =>
                           n17934, C1 => n25072, C2 => n17933, ZN => n23461);
   U21453 : OAI221_X1 port map( B1 => n20682, B2 => n25096, C1 => n21002, C2 =>
                           n25090, A => n23443, ZN => n23436);
   U21454 : AOI222_X1 port map( A1 => n25084, A2 => n24236, B1 => n25078, B2 =>
                           n17913, C1 => n25072, C2 => n17912, ZN => n23443);
   U21455 : OAI221_X1 port map( B1 => n20681, B2 => n25096, C1 => n21001, C2 =>
                           n25090, A => n23425, ZN => n23418);
   U21456 : AOI222_X1 port map( A1 => n25084, A2 => n24238, B1 => n25078, B2 =>
                           n17892, C1 => n25072, C2 => n17891, ZN => n23425);
   U21457 : OAI221_X1 port map( B1 => n20680, B2 => n25096, C1 => n21000, C2 =>
                           n25090, A => n23407, ZN => n23400);
   U21458 : AOI222_X1 port map( A1 => n25084, A2 => n24240, B1 => n25078, B2 =>
                           n17871, C1 => n25072, C2 => n17870, ZN => n23407);
   U21459 : OAI221_X1 port map( B1 => n20679, B2 => n25096, C1 => n20999, C2 =>
                           n25090, A => n23389, ZN => n23382);
   U21460 : AOI222_X1 port map( A1 => n25084, A2 => n24242, B1 => n25078, B2 =>
                           n17850, C1 => n25072, C2 => n17849, ZN => n23389);
   U21461 : OAI221_X1 port map( B1 => n20678, B2 => n25096, C1 => n20998, C2 =>
                           n25090, A => n23371, ZN => n23364);
   U21462 : AOI222_X1 port map( A1 => n25084, A2 => n24244, B1 => n25078, B2 =>
                           n17829, C1 => n25072, C2 => n17828, ZN => n23371);
   U21463 : OAI221_X1 port map( B1 => n20677, B2 => n25096, C1 => n20997, C2 =>
                           n25090, A => n23353, ZN => n23346);
   U21464 : AOI222_X1 port map( A1 => n25084, A2 => n24246, B1 => n25078, B2 =>
                           n17808, C1 => n25072, C2 => n17807, ZN => n23353);
   U21465 : OAI221_X1 port map( B1 => n20676, B2 => n25096, C1 => n20996, C2 =>
                           n25090, A => n23335, ZN => n23328);
   U21466 : AOI222_X1 port map( A1 => n25084, A2 => n24248, B1 => n25078, B2 =>
                           n17787, C1 => n25072, C2 => n17786, ZN => n23335);
   U21467 : OAI221_X1 port map( B1 => n20675, B2 => n25096, C1 => n20995, C2 =>
                           n25090, A => n23317, ZN => n23310);
   U21468 : AOI222_X1 port map( A1 => n25084, A2 => n24250, B1 => n25078, B2 =>
                           n17766, C1 => n25072, C2 => n17765, ZN => n23317);
   U21469 : OAI221_X1 port map( B1 => n20674, B2 => n25096, C1 => n20994, C2 =>
                           n25090, A => n23299, ZN => n23292);
   U21470 : AOI222_X1 port map( A1 => n25084, A2 => n24252, B1 => n25078, B2 =>
                           n17745, C1 => n25072, C2 => n17744, ZN => n23299);
   U21471 : OAI221_X1 port map( B1 => n20673, B2 => n25097, C1 => n20993, C2 =>
                           n25091, A => n23281, ZN => n23274);
   U21472 : AOI222_X1 port map( A1 => n25085, A2 => n24254, B1 => n25079, B2 =>
                           n17724, C1 => n25073, C2 => n17723, ZN => n23281);
   U21473 : OAI221_X1 port map( B1 => n20672, B2 => n25097, C1 => n20992, C2 =>
                           n25091, A => n23263, ZN => n23256);
   U21474 : AOI222_X1 port map( A1 => n25085, A2 => n24256, B1 => n25079, B2 =>
                           n17703, C1 => n25073, C2 => n17702, ZN => n23263);
   U21475 : OAI221_X1 port map( B1 => n20671, B2 => n25097, C1 => n20991, C2 =>
                           n25091, A => n23245, ZN => n23238);
   U21476 : AOI222_X1 port map( A1 => n25085, A2 => n24258, B1 => n25079, B2 =>
                           n17682, C1 => n25073, C2 => n17681, ZN => n23245);
   U21477 : OAI221_X1 port map( B1 => n20670, B2 => n25097, C1 => n20990, C2 =>
                           n25091, A => n23227, ZN => n23220);
   U21478 : AOI222_X1 port map( A1 => n25085, A2 => n24260, B1 => n25079, B2 =>
                           n17661, C1 => n25073, C2 => n17660, ZN => n23227);
   U21479 : OAI221_X1 port map( B1 => n20669, B2 => n25097, C1 => n20989, C2 =>
                           n25091, A => n23209, ZN => n23202);
   U21480 : AOI222_X1 port map( A1 => n25085, A2 => n24262, B1 => n25079, B2 =>
                           n17640, C1 => n25073, C2 => n17639, ZN => n23209);
   U21481 : OAI221_X1 port map( B1 => n20668, B2 => n25097, C1 => n20988, C2 =>
                           n25091, A => n23191, ZN => n23184);
   U21482 : AOI222_X1 port map( A1 => n25085, A2 => n24264, B1 => n25079, B2 =>
                           n17619, C1 => n25073, C2 => n17618, ZN => n23191);
   U21483 : OAI221_X1 port map( B1 => n20667, B2 => n25097, C1 => n20987, C2 =>
                           n25091, A => n23173, ZN => n23166);
   U21484 : AOI222_X1 port map( A1 => n25085, A2 => n24266, B1 => n25079, B2 =>
                           n17598, C1 => n25073, C2 => n17597, ZN => n23173);
   U21485 : OAI221_X1 port map( B1 => n20666, B2 => n25097, C1 => n20986, C2 =>
                           n25091, A => n23155, ZN => n23148);
   U21486 : AOI222_X1 port map( A1 => n25085, A2 => n24268, B1 => n25079, B2 =>
                           n17577, C1 => n25073, C2 => n17576, ZN => n23155);
   U21487 : OAI221_X1 port map( B1 => n20665, B2 => n25097, C1 => n20985, C2 =>
                           n25091, A => n23137, ZN => n23130);
   U21488 : AOI222_X1 port map( A1 => n25085, A2 => n24270, B1 => n25079, B2 =>
                           n17556, C1 => n25073, C2 => n17555, ZN => n23137);
   U21489 : OAI221_X1 port map( B1 => n20664, B2 => n25097, C1 => n20984, C2 =>
                           n25091, A => n23119, ZN => n23112);
   U21490 : AOI222_X1 port map( A1 => n25085, A2 => n24272, B1 => n25079, B2 =>
                           n17535, C1 => n25073, C2 => n17534, ZN => n23119);
   U21491 : OAI221_X1 port map( B1 => n20663, B2 => n25097, C1 => n20983, C2 =>
                           n25091, A => n23101, ZN => n23094);
   U21492 : AOI222_X1 port map( A1 => n25085, A2 => n24274, B1 => n25079, B2 =>
                           n17514, C1 => n25073, C2 => n17513, ZN => n23101);
   U21493 : OAI221_X1 port map( B1 => n20662, B2 => n25097, C1 => n20982, C2 =>
                           n25091, A => n23083, ZN => n23076);
   U21494 : AOI222_X1 port map( A1 => n25085, A2 => n24276, B1 => n25079, B2 =>
                           n17493, C1 => n25073, C2 => n17492, ZN => n23083);
   U21495 : OAI221_X1 port map( B1 => n20661, B2 => n25098, C1 => n20981, C2 =>
                           n25092, A => n23065, ZN => n23058);
   U21496 : AOI222_X1 port map( A1 => n25086, A2 => n24278, B1 => n25080, B2 =>
                           n17472, C1 => n25074, C2 => n17471, ZN => n23065);
   U21497 : OAI221_X1 port map( B1 => n20660, B2 => n25098, C1 => n20980, C2 =>
                           n25092, A => n23047, ZN => n23040);
   U21498 : AOI222_X1 port map( A1 => n25086, A2 => n24280, B1 => n25080, B2 =>
                           n17451, C1 => n25074, C2 => n17450, ZN => n23047);
   U21499 : OAI221_X1 port map( B1 => n20659, B2 => n25098, C1 => n20979, C2 =>
                           n25092, A => n23029, ZN => n23022);
   U21500 : AOI222_X1 port map( A1 => n25086, A2 => n24282, B1 => n25080, B2 =>
                           n17430, C1 => n25074, C2 => n17429, ZN => n23029);
   U21501 : OAI221_X1 port map( B1 => n20658, B2 => n25098, C1 => n20978, C2 =>
                           n25092, A => n23011, ZN => n23004);
   U21502 : AOI222_X1 port map( A1 => n25086, A2 => n24284, B1 => n25080, B2 =>
                           n17409, C1 => n25074, C2 => n17408, ZN => n23011);
   U21503 : OAI221_X1 port map( B1 => n20657, B2 => n25098, C1 => n20977, C2 =>
                           n25092, A => n22993, ZN => n22986);
   U21504 : AOI222_X1 port map( A1 => n25086, A2 => n24286, B1 => n25080, B2 =>
                           n17388, C1 => n25074, C2 => n17387, ZN => n22993);
   U21505 : OAI221_X1 port map( B1 => n20656, B2 => n25098, C1 => n20976, C2 =>
                           n25092, A => n22975, ZN => n22968);
   U21506 : AOI222_X1 port map( A1 => n25086, A2 => n24288, B1 => n25080, B2 =>
                           n17367, C1 => n25074, C2 => n17366, ZN => n22975);
   U21507 : OAI221_X1 port map( B1 => n20655, B2 => n25098, C1 => n20975, C2 =>
                           n25092, A => n22957, ZN => n22950);
   U21508 : AOI222_X1 port map( A1 => n25086, A2 => n24290, B1 => n25080, B2 =>
                           n17346, C1 => n25074, C2 => n17345, ZN => n22957);
   U21509 : OAI221_X1 port map( B1 => n20654, B2 => n25098, C1 => n20974, C2 =>
                           n25092, A => n22939, ZN => n22932);
   U21510 : AOI222_X1 port map( A1 => n25086, A2 => n24292, B1 => n25080, B2 =>
                           n17325, C1 => n25074, C2 => n17324, ZN => n22939);
   U21511 : OAI221_X1 port map( B1 => n20653, B2 => n25098, C1 => n20973, C2 =>
                           n25092, A => n22921, ZN => n22914);
   U21512 : AOI222_X1 port map( A1 => n25086, A2 => n24294, B1 => n25080, B2 =>
                           n17304, C1 => n25074, C2 => n17303, ZN => n22921);
   U21513 : OAI221_X1 port map( B1 => n20652, B2 => n25098, C1 => n20972, C2 =>
                           n25092, A => n22903, ZN => n22896);
   U21514 : AOI222_X1 port map( A1 => n25086, A2 => n24296, B1 => n25080, B2 =>
                           n17283, C1 => n25074, C2 => n17282, ZN => n22903);
   U21515 : OAI221_X1 port map( B1 => n20651, B2 => n25098, C1 => n20971, C2 =>
                           n25092, A => n22885, ZN => n22878);
   U21516 : AOI222_X1 port map( A1 => n25086, A2 => n24298, B1 => n25080, B2 =>
                           n17262, C1 => n25074, C2 => n17261, ZN => n22885);
   U21517 : OAI221_X1 port map( B1 => n20650, B2 => n25098, C1 => n20970, C2 =>
                           n25092, A => n22867, ZN => n22860);
   U21518 : AOI222_X1 port map( A1 => n25086, A2 => n24300, B1 => n25080, B2 =>
                           n17241, C1 => n25074, C2 => n17240, ZN => n22867);
   U21519 : OAI221_X1 port map( B1 => n20697, B2 => n25293, C1 => n21017, C2 =>
                           n25287, A => n22516, ZN => n22509);
   U21520 : AOI222_X1 port map( A1 => n25281, A2 => n24206, B1 => n25275, B2 =>
                           n18228, C1 => n25269, C2 => n18227, ZN => n22516);
   U21521 : OAI221_X1 port map( B1 => n20696, B2 => n25293, C1 => n21016, C2 =>
                           n25287, A => n22498, ZN => n22491);
   U21522 : AOI222_X1 port map( A1 => n25281, A2 => n24208, B1 => n25275, B2 =>
                           n18207, C1 => n25269, C2 => n18206, ZN => n22498);
   U21523 : OAI221_X1 port map( B1 => n20695, B2 => n25293, C1 => n21015, C2 =>
                           n25287, A => n22480, ZN => n22473);
   U21524 : AOI222_X1 port map( A1 => n25281, A2 => n24210, B1 => n25275, B2 =>
                           n18186, C1 => n25269, C2 => n18185, ZN => n22480);
   U21525 : OAI221_X1 port map( B1 => n20694, B2 => n25293, C1 => n21014, C2 =>
                           n25287, A => n22462, ZN => n22455);
   U21526 : AOI222_X1 port map( A1 => n25281, A2 => n24212, B1 => n25275, B2 =>
                           n18165, C1 => n25269, C2 => n18164, ZN => n22462);
   U21527 : OAI221_X1 port map( B1 => n20693, B2 => n25293, C1 => n21013, C2 =>
                           n25287, A => n22444, ZN => n22437);
   U21528 : AOI222_X1 port map( A1 => n25281, A2 => n24214, B1 => n25275, B2 =>
                           n18144, C1 => n25269, C2 => n18143, ZN => n22444);
   U21529 : OAI221_X1 port map( B1 => n20692, B2 => n25293, C1 => n21012, C2 =>
                           n25287, A => n22426, ZN => n22419);
   U21530 : AOI222_X1 port map( A1 => n25281, A2 => n24216, B1 => n25275, B2 =>
                           n18123, C1 => n25269, C2 => n18122, ZN => n22426);
   U21531 : OAI221_X1 port map( B1 => n20691, B2 => n25293, C1 => n21011, C2 =>
                           n25287, A => n22408, ZN => n22401);
   U21532 : AOI222_X1 port map( A1 => n25281, A2 => n24218, B1 => n25275, B2 =>
                           n18102, C1 => n25269, C2 => n18101, ZN => n22408);
   U21533 : OAI221_X1 port map( B1 => n20690, B2 => n25293, C1 => n21010, C2 =>
                           n25287, A => n22390, ZN => n22383);
   U21534 : AOI222_X1 port map( A1 => n25281, A2 => n24220, B1 => n25275, B2 =>
                           n18081, C1 => n25269, C2 => n18080, ZN => n22390);
   U21535 : OAI221_X1 port map( B1 => n20689, B2 => n25293, C1 => n21009, C2 =>
                           n25287, A => n22372, ZN => n22365);
   U21536 : AOI222_X1 port map( A1 => n25281, A2 => n24222, B1 => n25275, B2 =>
                           n18060, C1 => n25269, C2 => n18059, ZN => n22372);
   U21537 : OAI221_X1 port map( B1 => n20688, B2 => n25293, C1 => n21008, C2 =>
                           n25287, A => n22354, ZN => n22347);
   U21538 : AOI222_X1 port map( A1 => n25281, A2 => n24224, B1 => n25275, B2 =>
                           n18039, C1 => n25269, C2 => n18038, ZN => n22354);
   U21539 : OAI221_X1 port map( B1 => n20687, B2 => n25293, C1 => n21007, C2 =>
                           n25287, A => n22336, ZN => n22329);
   U21540 : AOI222_X1 port map( A1 => n25281, A2 => n24226, B1 => n25275, B2 =>
                           n18018, C1 => n25269, C2 => n18017, ZN => n22336);
   U21541 : OAI221_X1 port map( B1 => n20686, B2 => n25293, C1 => n21006, C2 =>
                           n25287, A => n22318, ZN => n22311);
   U21542 : AOI222_X1 port map( A1 => n25281, A2 => n24228, B1 => n25275, B2 =>
                           n17997, C1 => n25269, C2 => n17996, ZN => n22318);
   U21543 : OAI221_X1 port map( B1 => n20685, B2 => n25294, C1 => n21005, C2 =>
                           n25288, A => n22300, ZN => n22293);
   U21544 : AOI222_X1 port map( A1 => n25282, A2 => n24230, B1 => n25276, B2 =>
                           n17976, C1 => n25270, C2 => n17975, ZN => n22300);
   U21545 : OAI221_X1 port map( B1 => n20684, B2 => n25294, C1 => n21004, C2 =>
                           n25288, A => n22282, ZN => n22275);
   U21546 : AOI222_X1 port map( A1 => n25282, A2 => n24232, B1 => n25276, B2 =>
                           n17955, C1 => n25270, C2 => n17954, ZN => n22282);
   U21547 : OAI221_X1 port map( B1 => n20683, B2 => n25294, C1 => n21003, C2 =>
                           n25288, A => n22264, ZN => n22257);
   U21548 : AOI222_X1 port map( A1 => n25282, A2 => n24234, B1 => n25276, B2 =>
                           n17934, C1 => n25270, C2 => n17933, ZN => n22264);
   U21549 : OAI221_X1 port map( B1 => n20682, B2 => n25294, C1 => n21002, C2 =>
                           n25288, A => n22246, ZN => n22239);
   U21550 : AOI222_X1 port map( A1 => n25282, A2 => n24236, B1 => n25276, B2 =>
                           n17913, C1 => n25270, C2 => n17912, ZN => n22246);
   U21551 : OAI221_X1 port map( B1 => n20681, B2 => n25294, C1 => n21001, C2 =>
                           n25288, A => n22228, ZN => n22221);
   U21552 : AOI222_X1 port map( A1 => n25282, A2 => n24238, B1 => n25276, B2 =>
                           n17892, C1 => n25270, C2 => n17891, ZN => n22228);
   U21553 : OAI221_X1 port map( B1 => n20680, B2 => n25294, C1 => n21000, C2 =>
                           n25288, A => n22210, ZN => n22203);
   U21554 : AOI222_X1 port map( A1 => n25282, A2 => n24240, B1 => n25276, B2 =>
                           n17871, C1 => n25270, C2 => n17870, ZN => n22210);
   U21555 : OAI221_X1 port map( B1 => n20679, B2 => n25294, C1 => n20999, C2 =>
                           n25288, A => n22192, ZN => n22185);
   U21556 : AOI222_X1 port map( A1 => n25282, A2 => n24242, B1 => n25276, B2 =>
                           n17850, C1 => n25270, C2 => n17849, ZN => n22192);
   U21557 : OAI221_X1 port map( B1 => n20678, B2 => n25294, C1 => n20998, C2 =>
                           n25288, A => n22174, ZN => n22167);
   U21558 : AOI222_X1 port map( A1 => n25282, A2 => n24244, B1 => n25276, B2 =>
                           n17829, C1 => n25270, C2 => n17828, ZN => n22174);
   U21559 : OAI221_X1 port map( B1 => n20677, B2 => n25294, C1 => n20997, C2 =>
                           n25288, A => n22156, ZN => n22149);
   U21560 : AOI222_X1 port map( A1 => n25282, A2 => n24246, B1 => n25276, B2 =>
                           n17808, C1 => n25270, C2 => n17807, ZN => n22156);
   U21561 : OAI221_X1 port map( B1 => n20676, B2 => n25294, C1 => n20996, C2 =>
                           n25288, A => n22138, ZN => n22131);
   U21562 : AOI222_X1 port map( A1 => n25282, A2 => n24248, B1 => n25276, B2 =>
                           n17787, C1 => n25270, C2 => n17786, ZN => n22138);
   U21563 : OAI221_X1 port map( B1 => n20675, B2 => n25294, C1 => n20995, C2 =>
                           n25288, A => n22120, ZN => n22113);
   U21564 : AOI222_X1 port map( A1 => n25282, A2 => n24250, B1 => n25276, B2 =>
                           n17766, C1 => n25270, C2 => n17765, ZN => n22120);
   U21565 : OAI221_X1 port map( B1 => n20674, B2 => n25294, C1 => n20994, C2 =>
                           n25288, A => n22102, ZN => n22095);
   U21566 : AOI222_X1 port map( A1 => n25282, A2 => n24252, B1 => n25276, B2 =>
                           n17745, C1 => n25270, C2 => n17744, ZN => n22102);
   U21567 : OAI221_X1 port map( B1 => n20673, B2 => n25295, C1 => n20993, C2 =>
                           n25289, A => n22084, ZN => n22077);
   U21568 : AOI222_X1 port map( A1 => n25283, A2 => n24254, B1 => n25277, B2 =>
                           n17724, C1 => n25271, C2 => n17723, ZN => n22084);
   U21569 : OAI221_X1 port map( B1 => n20672, B2 => n25295, C1 => n20992, C2 =>
                           n25289, A => n22066, ZN => n22059);
   U21570 : AOI222_X1 port map( A1 => n25283, A2 => n24256, B1 => n25277, B2 =>
                           n17703, C1 => n25271, C2 => n17702, ZN => n22066);
   U21571 : OAI221_X1 port map( B1 => n20671, B2 => n25295, C1 => n20991, C2 =>
                           n25289, A => n22048, ZN => n22041);
   U21572 : AOI222_X1 port map( A1 => n25283, A2 => n24258, B1 => n25277, B2 =>
                           n17682, C1 => n25271, C2 => n17681, ZN => n22048);
   U21573 : OAI221_X1 port map( B1 => n20670, B2 => n25295, C1 => n20990, C2 =>
                           n25289, A => n22030, ZN => n22023);
   U21574 : AOI222_X1 port map( A1 => n25283, A2 => n24260, B1 => n25277, B2 =>
                           n17661, C1 => n25271, C2 => n17660, ZN => n22030);
   U21575 : OAI221_X1 port map( B1 => n20669, B2 => n25295, C1 => n20989, C2 =>
                           n25289, A => n22012, ZN => n22005);
   U21576 : AOI222_X1 port map( A1 => n25283, A2 => n24262, B1 => n25277, B2 =>
                           n17640, C1 => n25271, C2 => n17639, ZN => n22012);
   U21577 : OAI221_X1 port map( B1 => n20668, B2 => n25295, C1 => n20988, C2 =>
                           n25289, A => n21994, ZN => n21987);
   U21578 : AOI222_X1 port map( A1 => n25283, A2 => n24264, B1 => n25277, B2 =>
                           n17619, C1 => n25271, C2 => n17618, ZN => n21994);
   U21579 : OAI221_X1 port map( B1 => n20667, B2 => n25295, C1 => n20987, C2 =>
                           n25289, A => n21976, ZN => n21969);
   U21580 : AOI222_X1 port map( A1 => n25283, A2 => n24266, B1 => n25277, B2 =>
                           n17598, C1 => n25271, C2 => n17597, ZN => n21976);
   U21581 : OAI221_X1 port map( B1 => n20666, B2 => n25295, C1 => n20986, C2 =>
                           n25289, A => n21958, ZN => n21951);
   U21582 : AOI222_X1 port map( A1 => n25283, A2 => n24268, B1 => n25277, B2 =>
                           n17577, C1 => n25271, C2 => n17576, ZN => n21958);
   U21583 : OAI221_X1 port map( B1 => n20665, B2 => n25295, C1 => n20985, C2 =>
                           n25289, A => n21940, ZN => n21933);
   U21584 : AOI222_X1 port map( A1 => n25283, A2 => n24270, B1 => n25277, B2 =>
                           n17556, C1 => n25271, C2 => n17555, ZN => n21940);
   U21585 : OAI221_X1 port map( B1 => n20664, B2 => n25295, C1 => n20984, C2 =>
                           n25289, A => n21922, ZN => n21915);
   U21586 : AOI222_X1 port map( A1 => n25283, A2 => n24272, B1 => n25277, B2 =>
                           n17535, C1 => n25271, C2 => n17534, ZN => n21922);
   U21587 : OAI221_X1 port map( B1 => n20663, B2 => n25295, C1 => n20983, C2 =>
                           n25289, A => n21904, ZN => n21897);
   U21588 : AOI222_X1 port map( A1 => n25283, A2 => n24274, B1 => n25277, B2 =>
                           n17514, C1 => n25271, C2 => n17513, ZN => n21904);
   U21589 : OAI221_X1 port map( B1 => n20662, B2 => n25295, C1 => n20982, C2 =>
                           n25289, A => n21886, ZN => n21879);
   U21590 : AOI222_X1 port map( A1 => n25283, A2 => n24276, B1 => n25277, B2 =>
                           n17493, C1 => n25271, C2 => n17492, ZN => n21886);
   U21591 : OAI221_X1 port map( B1 => n20661, B2 => n25296, C1 => n20981, C2 =>
                           n25290, A => n21868, ZN => n21861);
   U21592 : AOI222_X1 port map( A1 => n25284, A2 => n24278, B1 => n25278, B2 =>
                           n17472, C1 => n25272, C2 => n17471, ZN => n21868);
   U21593 : OAI221_X1 port map( B1 => n20660, B2 => n25296, C1 => n20980, C2 =>
                           n25290, A => n21850, ZN => n21843);
   U21594 : AOI222_X1 port map( A1 => n25284, A2 => n24280, B1 => n25278, B2 =>
                           n17451, C1 => n25272, C2 => n17450, ZN => n21850);
   U21595 : OAI221_X1 port map( B1 => n20659, B2 => n25296, C1 => n20979, C2 =>
                           n25290, A => n21832, ZN => n21825);
   U21596 : AOI222_X1 port map( A1 => n25284, A2 => n24282, B1 => n25278, B2 =>
                           n17430, C1 => n25272, C2 => n17429, ZN => n21832);
   U21597 : OAI221_X1 port map( B1 => n20658, B2 => n25296, C1 => n20978, C2 =>
                           n25290, A => n21814, ZN => n21807);
   U21598 : AOI222_X1 port map( A1 => n25284, A2 => n24284, B1 => n25278, B2 =>
                           n17409, C1 => n25272, C2 => n17408, ZN => n21814);
   U21599 : OAI221_X1 port map( B1 => n20657, B2 => n25296, C1 => n20977, C2 =>
                           n25290, A => n21796, ZN => n21789);
   U21600 : AOI222_X1 port map( A1 => n25284, A2 => n24286, B1 => n25278, B2 =>
                           n17388, C1 => n25272, C2 => n17387, ZN => n21796);
   U21601 : OAI221_X1 port map( B1 => n20656, B2 => n25296, C1 => n20976, C2 =>
                           n25290, A => n21778, ZN => n21771);
   U21602 : AOI222_X1 port map( A1 => n25284, A2 => n24288, B1 => n25278, B2 =>
                           n17367, C1 => n25272, C2 => n17366, ZN => n21778);
   U21603 : OAI221_X1 port map( B1 => n20655, B2 => n25296, C1 => n20975, C2 =>
                           n25290, A => n21760, ZN => n21753);
   U21604 : AOI222_X1 port map( A1 => n25284, A2 => n24290, B1 => n25278, B2 =>
                           n17346, C1 => n25272, C2 => n17345, ZN => n21760);
   U21605 : OAI221_X1 port map( B1 => n20654, B2 => n25296, C1 => n20974, C2 =>
                           n25290, A => n21742, ZN => n21735);
   U21606 : AOI222_X1 port map( A1 => n25284, A2 => n24292, B1 => n25278, B2 =>
                           n17325, C1 => n25272, C2 => n17324, ZN => n21742);
   U21607 : OAI221_X1 port map( B1 => n20653, B2 => n25296, C1 => n20973, C2 =>
                           n25290, A => n21724, ZN => n21717);
   U21608 : AOI222_X1 port map( A1 => n25284, A2 => n24294, B1 => n25278, B2 =>
                           n17304, C1 => n25272, C2 => n17303, ZN => n21724);
   U21609 : OAI221_X1 port map( B1 => n20652, B2 => n25296, C1 => n20972, C2 =>
                           n25290, A => n21706, ZN => n21699);
   U21610 : AOI222_X1 port map( A1 => n25284, A2 => n24296, B1 => n25278, B2 =>
                           n17283, C1 => n25272, C2 => n17282, ZN => n21706);
   U21611 : OAI221_X1 port map( B1 => n20651, B2 => n25296, C1 => n20971, C2 =>
                           n25290, A => n21688, ZN => n21681);
   U21612 : AOI222_X1 port map( A1 => n25284, A2 => n24298, B1 => n25278, B2 =>
                           n17262, C1 => n25272, C2 => n17261, ZN => n21688);
   U21613 : OAI221_X1 port map( B1 => n20650, B2 => n25296, C1 => n20970, C2 =>
                           n25290, A => n21670, ZN => n21663);
   U21614 : AOI222_X1 port map( A1 => n25284, A2 => n24300, B1 => n25278, B2 =>
                           n17241, C1 => n25272, C2 => n17240, ZN => n21670);
   U21615 : OAI221_X1 port map( B1 => n20646, B2 => n25099, C1 => n20966, C2 =>
                           n25093, A => n22776, ZN => n22755);
   U21616 : AOI222_X1 port map( A1 => n25087, A2 => n24311, B1 => n25081, B2 =>
                           n17157, C1 => n25075, C2 => n17156, ZN => n22776);
   U21617 : OAI221_X1 port map( B1 => n20649, B2 => n25099, C1 => n20969, C2 =>
                           n25093, A => n22849, ZN => n22842);
   U21618 : AOI222_X1 port map( A1 => n25087, A2 => n24302, B1 => n25081, B2 =>
                           n17220, C1 => n25075, C2 => n17219, ZN => n22849);
   U21619 : OAI221_X1 port map( B1 => n20648, B2 => n25099, C1 => n20968, C2 =>
                           n25093, A => n22831, ZN => n22824);
   U21620 : AOI222_X1 port map( A1 => n25087, A2 => n24305, B1 => n25081, B2 =>
                           n17199, C1 => n25075, C2 => n17198, ZN => n22831);
   U21621 : OAI221_X1 port map( B1 => n20647, B2 => n25099, C1 => n20967, C2 =>
                           n25093, A => n22813, ZN => n22806);
   U21622 : AOI222_X1 port map( A1 => n25087, A2 => n24308, B1 => n25081, B2 =>
                           n17178, C1 => n25075, C2 => n17177, ZN => n22813);
   U21623 : OAI221_X1 port map( B1 => n20649, B2 => n25297, C1 => n20969, C2 =>
                           n25291, A => n21652, ZN => n21645);
   U21624 : AOI222_X1 port map( A1 => n25285, A2 => n24302, B1 => n25279, B2 =>
                           n17220, C1 => n25273, C2 => n17219, ZN => n21652);
   U21625 : OAI221_X1 port map( B1 => n20648, B2 => n25297, C1 => n20968, C2 =>
                           n25291, A => n21634, ZN => n21627);
   U21626 : AOI222_X1 port map( A1 => n25285, A2 => n24305, B1 => n25279, B2 =>
                           n17199, C1 => n25273, C2 => n17198, ZN => n21634);
   U21627 : OAI221_X1 port map( B1 => n20647, B2 => n25297, C1 => n20967, C2 =>
                           n25291, A => n21616, ZN => n21609);
   U21628 : AOI222_X1 port map( A1 => n25285, A2 => n24308, B1 => n25279, B2 =>
                           n17178, C1 => n25273, C2 => n17177, ZN => n21616);
   U21629 : OAI221_X1 port map( B1 => n20646, B2 => n25297, C1 => n20966, C2 =>
                           n25291, A => n21579, ZN => n21558);
   U21630 : AOI222_X1 port map( A1 => n25285, A2 => n24311, B1 => n25279, B2 =>
                           n17157, C1 => n25273, C2 => n17156, ZN => n21579);
   U21631 : OAI221_X1 port map( B1 => n21413, B2 => n25016, C1 => n20333, C2 =>
                           n25010, A => n23948, ZN => n23942);
   U21632 : AOI22_X1 port map( A1 => n25004, A2 => n24614, B1 => n24998, B2 => 
                           n18486, ZN => n23948);
   U21633 : OAI221_X1 port map( B1 => n21412, B2 => n25016, C1 => n20332, C2 =>
                           n25010, A => n23918, ZN => n23913);
   U21634 : AOI22_X1 port map( A1 => n25004, A2 => n24615, B1 => n24998, B2 => 
                           n18465, ZN => n23918);
   U21635 : OAI221_X1 port map( B1 => n21411, B2 => n25016, C1 => n20331, C2 =>
                           n25010, A => n23900, ZN => n23895);
   U21636 : AOI22_X1 port map( A1 => n25004, A2 => n24616, B1 => n24998, B2 => 
                           n18444, ZN => n23900);
   U21637 : OAI221_X1 port map( B1 => n21410, B2 => n25016, C1 => n20330, C2 =>
                           n25010, A => n23882, ZN => n23877);
   U21638 : AOI22_X1 port map( A1 => n25004, A2 => n24617, B1 => n24998, B2 => 
                           n18423, ZN => n23882);
   U21639 : OAI221_X1 port map( B1 => n21409, B2 => n25016, C1 => n20329, C2 =>
                           n25010, A => n23864, ZN => n23859);
   U21640 : AOI22_X1 port map( A1 => n25004, A2 => n24618, B1 => n24998, B2 => 
                           n18402, ZN => n23864);
   U21641 : OAI221_X1 port map( B1 => n21408, B2 => n25016, C1 => n20328, C2 =>
                           n25010, A => n23846, ZN => n23841);
   U21642 : AOI22_X1 port map( A1 => n25004, A2 => n24619, B1 => n24998, B2 => 
                           n18381, ZN => n23846);
   U21643 : OAI221_X1 port map( B1 => n21407, B2 => n25016, C1 => n20327, C2 =>
                           n25010, A => n23828, ZN => n23823);
   U21644 : AOI22_X1 port map( A1 => n25004, A2 => n24620, B1 => n24998, B2 => 
                           n18360, ZN => n23828);
   U21645 : OAI221_X1 port map( B1 => n21406, B2 => n25016, C1 => n20326, C2 =>
                           n25010, A => n23810, ZN => n23805);
   U21646 : AOI22_X1 port map( A1 => n25004, A2 => n24621, B1 => n24998, B2 => 
                           n18339, ZN => n23810);
   U21647 : OAI221_X1 port map( B1 => n21405, B2 => n25016, C1 => n20325, C2 =>
                           n25010, A => n23792, ZN => n23787);
   U21648 : AOI22_X1 port map( A1 => n25004, A2 => n24622, B1 => n24998, B2 => 
                           n18318, ZN => n23792);
   U21649 : OAI221_X1 port map( B1 => n21404, B2 => n25016, C1 => n20324, C2 =>
                           n25010, A => n23774, ZN => n23769);
   U21650 : AOI22_X1 port map( A1 => n25004, A2 => n24623, B1 => n24998, B2 => 
                           n18297, ZN => n23774);
   U21651 : OAI221_X1 port map( B1 => n21403, B2 => n25016, C1 => n20323, C2 =>
                           n25010, A => n23756, ZN => n23751);
   U21652 : AOI22_X1 port map( A1 => n25004, A2 => n24624, B1 => n24998, B2 => 
                           n18276, ZN => n23756);
   U21653 : OAI221_X1 port map( B1 => n21402, B2 => n25016, C1 => n20322, C2 =>
                           n25010, A => n23738, ZN => n23733);
   U21654 : AOI22_X1 port map( A1 => n25004, A2 => n24625, B1 => n24998, B2 => 
                           n18255, ZN => n23738);
   U21655 : OAI221_X1 port map( B1 => n21413, B2 => n25214, C1 => n20333, C2 =>
                           n25208, A => n22751, ZN => n22745);
   U21656 : AOI22_X1 port map( A1 => n25202, A2 => n24614, B1 => n25196, B2 => 
                           n18486, ZN => n22751);
   U21657 : OAI221_X1 port map( B1 => n21412, B2 => n25214, C1 => n20332, C2 =>
                           n25208, A => n22721, ZN => n22716);
   U21658 : AOI22_X1 port map( A1 => n25202, A2 => n24615, B1 => n25196, B2 => 
                           n18465, ZN => n22721);
   U21659 : OAI221_X1 port map( B1 => n21411, B2 => n25214, C1 => n20331, C2 =>
                           n25208, A => n22703, ZN => n22698);
   U21660 : AOI22_X1 port map( A1 => n25202, A2 => n24616, B1 => n25196, B2 => 
                           n18444, ZN => n22703);
   U21661 : OAI221_X1 port map( B1 => n21410, B2 => n25214, C1 => n20330, C2 =>
                           n25208, A => n22685, ZN => n22680);
   U21662 : AOI22_X1 port map( A1 => n25202, A2 => n24617, B1 => n25196, B2 => 
                           n18423, ZN => n22685);
   U21663 : OAI221_X1 port map( B1 => n21409, B2 => n25214, C1 => n20329, C2 =>
                           n25208, A => n22667, ZN => n22662);
   U21664 : AOI22_X1 port map( A1 => n25202, A2 => n24618, B1 => n25196, B2 => 
                           n18402, ZN => n22667);
   U21665 : OAI221_X1 port map( B1 => n21408, B2 => n25214, C1 => n20328, C2 =>
                           n25208, A => n22649, ZN => n22644);
   U21666 : AOI22_X1 port map( A1 => n25202, A2 => n24619, B1 => n25196, B2 => 
                           n18381, ZN => n22649);
   U21667 : OAI221_X1 port map( B1 => n21407, B2 => n25214, C1 => n20327, C2 =>
                           n25208, A => n22631, ZN => n22626);
   U21668 : AOI22_X1 port map( A1 => n25202, A2 => n24620, B1 => n25196, B2 => 
                           n18360, ZN => n22631);
   U21669 : OAI221_X1 port map( B1 => n21406, B2 => n25214, C1 => n20326, C2 =>
                           n25208, A => n22613, ZN => n22608);
   U21670 : AOI22_X1 port map( A1 => n25202, A2 => n24621, B1 => n25196, B2 => 
                           n18339, ZN => n22613);
   U21671 : OAI221_X1 port map( B1 => n21405, B2 => n25214, C1 => n20325, C2 =>
                           n25208, A => n22595, ZN => n22590);
   U21672 : AOI22_X1 port map( A1 => n25202, A2 => n24622, B1 => n25196, B2 => 
                           n18318, ZN => n22595);
   U21673 : OAI221_X1 port map( B1 => n21404, B2 => n25214, C1 => n20324, C2 =>
                           n25208, A => n22577, ZN => n22572);
   U21674 : AOI22_X1 port map( A1 => n25202, A2 => n24623, B1 => n25196, B2 => 
                           n18297, ZN => n22577);
   U21675 : OAI221_X1 port map( B1 => n21403, B2 => n25214, C1 => n20323, C2 =>
                           n25208, A => n22559, ZN => n22554);
   U21676 : AOI22_X1 port map( A1 => n25202, A2 => n24624, B1 => n25196, B2 => 
                           n18276, ZN => n22559);
   U21677 : OAI221_X1 port map( B1 => n21402, B2 => n25214, C1 => n20322, C2 =>
                           n25208, A => n22541, ZN => n22536);
   U21678 : AOI22_X1 port map( A1 => n25202, A2 => n24625, B1 => n25196, B2 => 
                           n18255, ZN => n22541);
   U21679 : OAI221_X1 port map( B1 => n20709, B2 => n25094, C1 => n21029, C2 =>
                           n25088, A => n23938, ZN => n23922);
   U21680 : AOI222_X1 port map( A1 => n25082, A2 => n24314, B1 => n25076, B2 =>
                           n18480, C1 => n25070, C2 => n18479, ZN => n23938);
   U21681 : OAI221_X1 port map( B1 => n20708, B2 => n25094, C1 => n21028, C2 =>
                           n25088, A => n23911, ZN => n23904);
   U21682 : AOI222_X1 port map( A1 => n25082, A2 => n24316, B1 => n25076, B2 =>
                           n18459, C1 => n25070, C2 => n18458, ZN => n23911);
   U21683 : OAI221_X1 port map( B1 => n20707, B2 => n25094, C1 => n21027, C2 =>
                           n25088, A => n23893, ZN => n23886);
   U21684 : AOI222_X1 port map( A1 => n25082, A2 => n24318, B1 => n25076, B2 =>
                           n18438, C1 => n25070, C2 => n18437, ZN => n23893);
   U21685 : OAI221_X1 port map( B1 => n20706, B2 => n25094, C1 => n21026, C2 =>
                           n25088, A => n23875, ZN => n23868);
   U21686 : AOI222_X1 port map( A1 => n25082, A2 => n24320, B1 => n25076, B2 =>
                           n18417, C1 => n25070, C2 => n18416, ZN => n23875);
   U21687 : OAI221_X1 port map( B1 => n20705, B2 => n25094, C1 => n21025, C2 =>
                           n25088, A => n23857, ZN => n23850);
   U21688 : AOI222_X1 port map( A1 => n25082, A2 => n24322, B1 => n25076, B2 =>
                           n18396, C1 => n25070, C2 => n18395, ZN => n23857);
   U21689 : OAI221_X1 port map( B1 => n20704, B2 => n25094, C1 => n21024, C2 =>
                           n25088, A => n23839, ZN => n23832);
   U21690 : AOI222_X1 port map( A1 => n25082, A2 => n24324, B1 => n25076, B2 =>
                           n18375, C1 => n25070, C2 => n18374, ZN => n23839);
   U21691 : OAI221_X1 port map( B1 => n20703, B2 => n25094, C1 => n21023, C2 =>
                           n25088, A => n23821, ZN => n23814);
   U21692 : AOI222_X1 port map( A1 => n25082, A2 => n24326, B1 => n25076, B2 =>
                           n18354, C1 => n25070, C2 => n18353, ZN => n23821);
   U21693 : OAI221_X1 port map( B1 => n20702, B2 => n25094, C1 => n21022, C2 =>
                           n25088, A => n23803, ZN => n23796);
   U21694 : AOI222_X1 port map( A1 => n25082, A2 => n24328, B1 => n25076, B2 =>
                           n18333, C1 => n25070, C2 => n18332, ZN => n23803);
   U21695 : OAI221_X1 port map( B1 => n20701, B2 => n25094, C1 => n21021, C2 =>
                           n25088, A => n23785, ZN => n23778);
   U21696 : AOI222_X1 port map( A1 => n25082, A2 => n24330, B1 => n25076, B2 =>
                           n18312, C1 => n25070, C2 => n18311, ZN => n23785);
   U21697 : OAI221_X1 port map( B1 => n20700, B2 => n25094, C1 => n21020, C2 =>
                           n25088, A => n23767, ZN => n23760);
   U21698 : AOI222_X1 port map( A1 => n25082, A2 => n24332, B1 => n25076, B2 =>
                           n18291, C1 => n25070, C2 => n18290, ZN => n23767);
   U21699 : OAI221_X1 port map( B1 => n20699, B2 => n25094, C1 => n21019, C2 =>
                           n25088, A => n23749, ZN => n23742);
   U21700 : AOI222_X1 port map( A1 => n25082, A2 => n24334, B1 => n25076, B2 =>
                           n18270, C1 => n25070, C2 => n18269, ZN => n23749);
   U21701 : OAI221_X1 port map( B1 => n20698, B2 => n25094, C1 => n21018, C2 =>
                           n25088, A => n23731, ZN => n23724);
   U21702 : AOI222_X1 port map( A1 => n25082, A2 => n24336, B1 => n25076, B2 =>
                           n18249, C1 => n25070, C2 => n18248, ZN => n23731);
   U21703 : OAI221_X1 port map( B1 => n20709, B2 => n25292, C1 => n21029, C2 =>
                           n25286, A => n22741, ZN => n22725);
   U21704 : AOI222_X1 port map( A1 => n25280, A2 => n24314, B1 => n25274, B2 =>
                           n18480, C1 => n25268, C2 => n18479, ZN => n22741);
   U21705 : OAI221_X1 port map( B1 => n20708, B2 => n25292, C1 => n21028, C2 =>
                           n25286, A => n22714, ZN => n22707);
   U21706 : AOI222_X1 port map( A1 => n25280, A2 => n24316, B1 => n25274, B2 =>
                           n18459, C1 => n25268, C2 => n18458, ZN => n22714);
   U21707 : OAI221_X1 port map( B1 => n20707, B2 => n25292, C1 => n21027, C2 =>
                           n25286, A => n22696, ZN => n22689);
   U21708 : AOI222_X1 port map( A1 => n25280, A2 => n24318, B1 => n25274, B2 =>
                           n18438, C1 => n25268, C2 => n18437, ZN => n22696);
   U21709 : OAI221_X1 port map( B1 => n20706, B2 => n25292, C1 => n21026, C2 =>
                           n25286, A => n22678, ZN => n22671);
   U21710 : AOI222_X1 port map( A1 => n25280, A2 => n24320, B1 => n25274, B2 =>
                           n18417, C1 => n25268, C2 => n18416, ZN => n22678);
   U21711 : OAI221_X1 port map( B1 => n20705, B2 => n25292, C1 => n21025, C2 =>
                           n25286, A => n22660, ZN => n22653);
   U21712 : AOI222_X1 port map( A1 => n25280, A2 => n24322, B1 => n25274, B2 =>
                           n18396, C1 => n25268, C2 => n18395, ZN => n22660);
   U21713 : OAI221_X1 port map( B1 => n20704, B2 => n25292, C1 => n21024, C2 =>
                           n25286, A => n22642, ZN => n22635);
   U21714 : AOI222_X1 port map( A1 => n25280, A2 => n24324, B1 => n25274, B2 =>
                           n18375, C1 => n25268, C2 => n18374, ZN => n22642);
   U21715 : OAI221_X1 port map( B1 => n20703, B2 => n25292, C1 => n21023, C2 =>
                           n25286, A => n22624, ZN => n22617);
   U21716 : AOI222_X1 port map( A1 => n25280, A2 => n24326, B1 => n25274, B2 =>
                           n18354, C1 => n25268, C2 => n18353, ZN => n22624);
   U21717 : OAI221_X1 port map( B1 => n20702, B2 => n25292, C1 => n21022, C2 =>
                           n25286, A => n22606, ZN => n22599);
   U21718 : AOI222_X1 port map( A1 => n25280, A2 => n24328, B1 => n25274, B2 =>
                           n18333, C1 => n25268, C2 => n18332, ZN => n22606);
   U21719 : OAI221_X1 port map( B1 => n20701, B2 => n25292, C1 => n21021, C2 =>
                           n25286, A => n22588, ZN => n22581);
   U21720 : AOI222_X1 port map( A1 => n25280, A2 => n24330, B1 => n25274, B2 =>
                           n18312, C1 => n25268, C2 => n18311, ZN => n22588);
   U21721 : OAI221_X1 port map( B1 => n20700, B2 => n25292, C1 => n21020, C2 =>
                           n25286, A => n22570, ZN => n22563);
   U21722 : AOI222_X1 port map( A1 => n25280, A2 => n24332, B1 => n25274, B2 =>
                           n18291, C1 => n25268, C2 => n18290, ZN => n22570);
   U21723 : OAI221_X1 port map( B1 => n20699, B2 => n25292, C1 => n21019, C2 =>
                           n25286, A => n22552, ZN => n22545);
   U21724 : AOI222_X1 port map( A1 => n25280, A2 => n24334, B1 => n25274, B2 =>
                           n18270, C1 => n25268, C2 => n18269, ZN => n22552);
   U21725 : OAI221_X1 port map( B1 => n20698, B2 => n25292, C1 => n21018, C2 =>
                           n25286, A => n22534, ZN => n22527);
   U21726 : AOI222_X1 port map( A1 => n25280, A2 => n24336, B1 => n25274, B2 =>
                           n18249, C1 => n25268, C2 => n18248, ZN => n22534);
   U21727 : OAI22_X1 port map( A1 => n9466, A2 => n25776, B1 => n25770, B2 => 
                           n25817, ZN => n7435);
   U21728 : OAI22_X1 port map( A1 => n9465, A2 => n25776, B1 => n25770, B2 => 
                           n25820, ZN => n7436);
   U21729 : OAI22_X1 port map( A1 => n9464, A2 => n25776, B1 => n25770, B2 => 
                           n25823, ZN => n7437);
   U21730 : OAI22_X1 port map( A1 => n9463, A2 => n25776, B1 => n25770, B2 => 
                           n25826, ZN => n7438);
   U21731 : OAI22_X1 port map( A1 => n9462, A2 => n25776, B1 => n25770, B2 => 
                           n25829, ZN => n7439);
   U21732 : OAI22_X1 port map( A1 => n9461, A2 => n25776, B1 => n25770, B2 => 
                           n25832, ZN => n7440);
   U21733 : OAI22_X1 port map( A1 => n9460, A2 => n25776, B1 => n25770, B2 => 
                           n25835, ZN => n7441);
   U21734 : OAI22_X1 port map( A1 => n9459, A2 => n25776, B1 => n25770, B2 => 
                           n25838, ZN => n7442);
   U21735 : OAI22_X1 port map( A1 => n9458, A2 => n25776, B1 => n25770, B2 => 
                           n25841, ZN => n7443);
   U21736 : OAI22_X1 port map( A1 => n9457, A2 => n25776, B1 => n25770, B2 => 
                           n25844, ZN => n7444);
   U21737 : OAI22_X1 port map( A1 => n9456, A2 => n25776, B1 => n25770, B2 => 
                           n25847, ZN => n7445);
   U21738 : OAI22_X1 port map( A1 => n9455, A2 => n25777, B1 => n25770, B2 => 
                           n25850, ZN => n7446);
   U21739 : OAI22_X1 port map( A1 => n9454, A2 => n25777, B1 => n25771, B2 => 
                           n25853, ZN => n7447);
   U21740 : OAI22_X1 port map( A1 => n9453, A2 => n25777, B1 => n25771, B2 => 
                           n25856, ZN => n7448);
   U21741 : OAI22_X1 port map( A1 => n9452, A2 => n25777, B1 => n25771, B2 => 
                           n25859, ZN => n7449);
   U21742 : OAI22_X1 port map( A1 => n9451, A2 => n25777, B1 => n25771, B2 => 
                           n25862, ZN => n7450);
   U21743 : OAI22_X1 port map( A1 => n9450, A2 => n25777, B1 => n25771, B2 => 
                           n25865, ZN => n7451);
   U21744 : OAI22_X1 port map( A1 => n9449, A2 => n25777, B1 => n25771, B2 => 
                           n25868, ZN => n7452);
   U21745 : OAI22_X1 port map( A1 => n9448, A2 => n25777, B1 => n25771, B2 => 
                           n25871, ZN => n7453);
   U21746 : OAI22_X1 port map( A1 => n9447, A2 => n25777, B1 => n25771, B2 => 
                           n25874, ZN => n7454);
   U21747 : OAI22_X1 port map( A1 => n9446, A2 => n25777, B1 => n25771, B2 => 
                           n25877, ZN => n7455);
   U21748 : OAI22_X1 port map( A1 => n9445, A2 => n25777, B1 => n25771, B2 => 
                           n25880, ZN => n7456);
   U21749 : OAI22_X1 port map( A1 => n9444, A2 => n25777, B1 => n25771, B2 => 
                           n25883, ZN => n7457);
   U21750 : OAI22_X1 port map( A1 => n9443, A2 => n25778, B1 => n25771, B2 => 
                           n25886, ZN => n7458);
   U21751 : OAI22_X1 port map( A1 => n9442, A2 => n25778, B1 => n25772, B2 => 
                           n25889, ZN => n7459);
   U21752 : OAI22_X1 port map( A1 => n9441, A2 => n25778, B1 => n25772, B2 => 
                           n25892, ZN => n7460);
   U21753 : OAI22_X1 port map( A1 => n9440, A2 => n25778, B1 => n25772, B2 => 
                           n25895, ZN => n7461);
   U21754 : OAI22_X1 port map( A1 => n9439, A2 => n25778, B1 => n25772, B2 => 
                           n25898, ZN => n7462);
   U21755 : OAI22_X1 port map( A1 => n9438, A2 => n25778, B1 => n25772, B2 => 
                           n25901, ZN => n7463);
   U21756 : OAI22_X1 port map( A1 => n9437, A2 => n25778, B1 => n25772, B2 => 
                           n25904, ZN => n7464);
   U21757 : OAI22_X1 port map( A1 => n9436, A2 => n25778, B1 => n25772, B2 => 
                           n25907, ZN => n7465);
   U21758 : OAI22_X1 port map( A1 => n9435, A2 => n25778, B1 => n25772, B2 => 
                           n25910, ZN => n7466);
   U21759 : OAI22_X1 port map( A1 => n9434, A2 => n25778, B1 => n25772, B2 => 
                           n25913, ZN => n7467);
   U21760 : OAI22_X1 port map( A1 => n9433, A2 => n25778, B1 => n25772, B2 => 
                           n25916, ZN => n7468);
   U21761 : OAI22_X1 port map( A1 => n9432, A2 => n25778, B1 => n25772, B2 => 
                           n25919, ZN => n7469);
   U21762 : OAI22_X1 port map( A1 => n9431, A2 => n25779, B1 => n25772, B2 => 
                           n25922, ZN => n7470);
   U21763 : OAI22_X1 port map( A1 => n9430, A2 => n25779, B1 => n25773, B2 => 
                           n25925, ZN => n7471);
   U21764 : OAI22_X1 port map( A1 => n9429, A2 => n25779, B1 => n25773, B2 => 
                           n25928, ZN => n7472);
   U21765 : OAI22_X1 port map( A1 => n9428, A2 => n25779, B1 => n25773, B2 => 
                           n25931, ZN => n7473);
   U21766 : OAI22_X1 port map( A1 => n9427, A2 => n25779, B1 => n25773, B2 => 
                           n25934, ZN => n7474);
   U21767 : OAI22_X1 port map( A1 => n9426, A2 => n25779, B1 => n25773, B2 => 
                           n25937, ZN => n7475);
   U21768 : OAI22_X1 port map( A1 => n9425, A2 => n25779, B1 => n25773, B2 => 
                           n25940, ZN => n7476);
   U21769 : OAI22_X1 port map( A1 => n9424, A2 => n25779, B1 => n25773, B2 => 
                           n25943, ZN => n7477);
   U21770 : OAI22_X1 port map( A1 => n9423, A2 => n25779, B1 => n25773, B2 => 
                           n25946, ZN => n7478);
   U21771 : OAI22_X1 port map( A1 => n9422, A2 => n25779, B1 => n25773, B2 => 
                           n25949, ZN => n7479);
   U21772 : OAI22_X1 port map( A1 => n9421, A2 => n25779, B1 => n25773, B2 => 
                           n25952, ZN => n7480);
   U21773 : OAI22_X1 port map( A1 => n9420, A2 => n25779, B1 => n25773, B2 => 
                           n25955, ZN => n7481);
   U21774 : OAI22_X1 port map( A1 => n9419, A2 => n25780, B1 => n25773, B2 => 
                           n25958, ZN => n7482);
   U21775 : OAI22_X1 port map( A1 => n9418, A2 => n25780, B1 => n25774, B2 => 
                           n25961, ZN => n7483);
   U21776 : OAI22_X1 port map( A1 => n9417, A2 => n25780, B1 => n25774, B2 => 
                           n25964, ZN => n7484);
   U21777 : OAI22_X1 port map( A1 => n9416, A2 => n25780, B1 => n25774, B2 => 
                           n25967, ZN => n7485);
   U21778 : OAI22_X1 port map( A1 => n9415, A2 => n25780, B1 => n25774, B2 => 
                           n25970, ZN => n7486);
   U21779 : OAI22_X1 port map( A1 => n25601, A2 => n21417, B1 => n25962, B2 => 
                           n25594, ZN => n6587);
   U21780 : OAI22_X1 port map( A1 => n25601, A2 => n21416, B1 => n25965, B2 => 
                           n25594, ZN => n6588);
   U21781 : OAI22_X1 port map( A1 => n25601, A2 => n21415, B1 => n25968, B2 => 
                           n25594, ZN => n6589);
   U21782 : OAI22_X1 port map( A1 => n25601, A2 => n21414, B1 => n25971, B2 => 
                           n25594, ZN => n6590);
   U21783 : OAI22_X1 port map( A1 => n25473, A2 => n21289, B1 => n25962, B2 => 
                           n25466, ZN => n5947);
   U21784 : OAI22_X1 port map( A1 => n25473, A2 => n21288, B1 => n25965, B2 => 
                           n25466, ZN => n5948);
   U21785 : OAI22_X1 port map( A1 => n25473, A2 => n21287, B1 => n25968, B2 => 
                           n25466, ZN => n5949);
   U21786 : OAI22_X1 port map( A1 => n25473, A2 => n21286, B1 => n25971, B2 => 
                           n25466, ZN => n5950);
   U21787 : OAI22_X1 port map( A1 => n25486, A2 => n21033, B1 => n25962, B2 => 
                           n25479, ZN => n6011);
   U21788 : OAI22_X1 port map( A1 => n25486, A2 => n21032, B1 => n25965, B2 => 
                           n25479, ZN => n6012);
   U21789 : OAI22_X1 port map( A1 => n25486, A2 => n21031, B1 => n25968, B2 => 
                           n25479, ZN => n6013);
   U21790 : OAI22_X1 port map( A1 => n25486, A2 => n21030, B1 => n25971, B2 => 
                           n25479, ZN => n6014);
   U21791 : OAI22_X1 port map( A1 => n25576, A2 => n20905, B1 => n25962, B2 => 
                           n25569, ZN => n6459);
   U21792 : OAI22_X1 port map( A1 => n25576, A2 => n20904, B1 => n25965, B2 => 
                           n25569, ZN => n6460);
   U21793 : OAI22_X1 port map( A1 => n25576, A2 => n20903, B1 => n25968, B2 => 
                           n25569, ZN => n6461);
   U21794 : OAI22_X1 port map( A1 => n25576, A2 => n20902, B1 => n25971, B2 => 
                           n25569, ZN => n6462);
   U21795 : OAI22_X1 port map( A1 => n25460, A2 => n20781, B1 => n25963, B2 => 
                           n25453, ZN => n5883);
   U21796 : OAI22_X1 port map( A1 => n25460, A2 => n20780, B1 => n25966, B2 => 
                           n25453, ZN => n5884);
   U21797 : OAI22_X1 port map( A1 => n25460, A2 => n20779, B1 => n25969, B2 => 
                           n25453, ZN => n5885);
   U21798 : OAI22_X1 port map( A1 => n25460, A2 => n20778, B1 => n25972, B2 => 
                           n25453, ZN => n5886);
   U21799 : OAI22_X1 port map( A1 => n25653, A2 => n20585, B1 => n25961, B2 => 
                           n25646, ZN => n6843);
   U21800 : OAI22_X1 port map( A1 => n25653, A2 => n20584, B1 => n25964, B2 => 
                           n25646, ZN => n6844);
   U21801 : OAI22_X1 port map( A1 => n25653, A2 => n20583, B1 => n25967, B2 => 
                           n25646, ZN => n6845);
   U21802 : OAI22_X1 port map( A1 => n25653, A2 => n20582, B1 => n25970, B2 => 
                           n25646, ZN => n6846);
   U21803 : OAI22_X1 port map( A1 => n25421, A2 => n20269, B1 => n25963, B2 => 
                           n25414, ZN => n5691);
   U21804 : OAI22_X1 port map( A1 => n25421, A2 => n20268, B1 => n25966, B2 => 
                           n25414, ZN => n5692);
   U21805 : OAI22_X1 port map( A1 => n25421, A2 => n20267, B1 => n25969, B2 => 
                           n25414, ZN => n5693);
   U21806 : OAI22_X1 port map( A1 => n25421, A2 => n20266, B1 => n25972, B2 => 
                           n25414, ZN => n5694);
   U21807 : OAI22_X1 port map( A1 => n25395, A2 => n20265, B1 => n25963, B2 => 
                           n25388, ZN => n5563);
   U21808 : OAI22_X1 port map( A1 => n25395, A2 => n20264, B1 => n25966, B2 => 
                           n25388, ZN => n5564);
   U21809 : OAI22_X1 port map( A1 => n25395, A2 => n20263, B1 => n25969, B2 => 
                           n25388, ZN => n5565);
   U21810 : OAI22_X1 port map( A1 => n25395, A2 => n20262, B1 => n25972, B2 => 
                           n25388, ZN => n5566);
   U21811 : OAI22_X1 port map( A1 => n25743, A2 => n20201, B1 => n25961, B2 => 
                           n25736, ZN => n7291);
   U21812 : OAI22_X1 port map( A1 => n25743, A2 => n20200, B1 => n25964, B2 => 
                           n25736, ZN => n7292);
   U21813 : OAI22_X1 port map( A1 => n25743, A2 => n20199, B1 => n25967, B2 => 
                           n25736, ZN => n7293);
   U21814 : OAI22_X1 port map( A1 => n25743, A2 => n20198, B1 => n25970, B2 => 
                           n25736, ZN => n7294);
   U21815 : OAI22_X1 port map( A1 => n9226, A2 => n25588, B1 => n25962, B2 => 
                           n25582, ZN => n6523);
   U21816 : OAI22_X1 port map( A1 => n9225, A2 => n25588, B1 => n25965, B2 => 
                           n25582, ZN => n6524);
   U21817 : OAI22_X1 port map( A1 => n9224, A2 => n25588, B1 => n25968, B2 => 
                           n25582, ZN => n6525);
   U21818 : OAI22_X1 port map( A1 => n9223, A2 => n25588, B1 => n25971, B2 => 
                           n25582, ZN => n6526);
   U21819 : OAI22_X1 port map( A1 => n8970, A2 => n25511, B1 => n25962, B2 => 
                           n25505, ZN => n6139);
   U21820 : OAI22_X1 port map( A1 => n8969, A2 => n25511, B1 => n25965, B2 => 
                           n25505, ZN => n6140);
   U21821 : OAI22_X1 port map( A1 => n8968, A2 => n25511, B1 => n25968, B2 => 
                           n25505, ZN => n6141);
   U21822 : OAI22_X1 port map( A1 => n8967, A2 => n25511, B1 => n25971, B2 => 
                           n25505, ZN => n6142);
   U21823 : OAI22_X1 port map( A1 => n9034, A2 => n25755, B1 => n25961, B2 => 
                           n25749, ZN => n7355);
   U21824 : OAI22_X1 port map( A1 => n9033, A2 => n25755, B1 => n25964, B2 => 
                           n25749, ZN => n7356);
   U21825 : OAI22_X1 port map( A1 => n9032, A2 => n25755, B1 => n25967, B2 => 
                           n25749, ZN => n7357);
   U21826 : OAI22_X1 port map( A1 => n9031, A2 => n25755, B1 => n25970, B2 => 
                           n25749, ZN => n7358);
   U21827 : OAI22_X1 port map( A1 => n9290, A2 => n25691, B1 => n25961, B2 => 
                           n25685, ZN => n7035);
   U21828 : OAI22_X1 port map( A1 => n9289, A2 => n25691, B1 => n25964, B2 => 
                           n25685, ZN => n7036);
   U21829 : OAI22_X1 port map( A1 => n9288, A2 => n25691, B1 => n25967, B2 => 
                           n25685, ZN => n7037);
   U21830 : OAI22_X1 port map( A1 => n9287, A2 => n25691, B1 => n25970, B2 => 
                           n25685, ZN => n7038);
   U21831 : OAI22_X1 port map( A1 => n25499, A2 => n19880, B1 => n25962, B2 => 
                           n25492, ZN => n6075);
   U21832 : OAI22_X1 port map( A1 => n25499, A2 => n19879, B1 => n25965, B2 => 
                           n25492, ZN => n6076);
   U21833 : OAI22_X1 port map( A1 => n25499, A2 => n19878, B1 => n25968, B2 => 
                           n25492, ZN => n6077);
   U21834 : OAI22_X1 port map( A1 => n25499, A2 => n19877, B1 => n25971, B2 => 
                           n25492, ZN => n6078);
   U21835 : OAI22_X1 port map( A1 => n25679, A2 => n19689, B1 => n25961, B2 => 
                           n25672, ZN => n6971);
   U21836 : OAI22_X1 port map( A1 => n25679, A2 => n19688, B1 => n25964, B2 => 
                           n25672, ZN => n6972);
   U21837 : OAI22_X1 port map( A1 => n25679, A2 => n19687, B1 => n25967, B2 => 
                           n25672, ZN => n6973);
   U21838 : OAI22_X1 port map( A1 => n25679, A2 => n19686, B1 => n25970, B2 => 
                           n25672, ZN => n6974);
   U21839 : OAI22_X1 port map( A1 => n25704, A2 => n19625, B1 => n25961, B2 => 
                           n25697, ZN => n7099);
   U21840 : OAI22_X1 port map( A1 => n25704, A2 => n19624, B1 => n25964, B2 => 
                           n25697, ZN => n7100);
   U21841 : OAI22_X1 port map( A1 => n25704, A2 => n19623, B1 => n25967, B2 => 
                           n25697, ZN => n7101);
   U21842 : OAI22_X1 port map( A1 => n25704, A2 => n19622, B1 => n25970, B2 => 
                           n25697, ZN => n7102);
   U21843 : AOI22_X1 port map( A1 => n24985, A2 => n19941, B1 => n24979, B2 => 
                           n24477, ZN => n22801);
   U21844 : AOI22_X1 port map( A1 => n24980, A2 => n20004, B1 => n24974, B2 => 
                           n24794, ZN => n23949);
   U21845 : AOI22_X1 port map( A1 => n24980, A2 => n20003, B1 => n24974, B2 => 
                           n24795, ZN => n23919);
   U21846 : AOI22_X1 port map( A1 => n24980, A2 => n20002, B1 => n24974, B2 => 
                           n24796, ZN => n23901);
   U21847 : AOI22_X1 port map( A1 => n24980, A2 => n20001, B1 => n24974, B2 => 
                           n24797, ZN => n23883);
   U21848 : AOI22_X1 port map( A1 => n24980, A2 => n20000, B1 => n24974, B2 => 
                           n24798, ZN => n23865);
   U21849 : AOI22_X1 port map( A1 => n24980, A2 => n19999, B1 => n24974, B2 => 
                           n24799, ZN => n23847);
   U21850 : AOI22_X1 port map( A1 => n24980, A2 => n19998, B1 => n24974, B2 => 
                           n24800, ZN => n23829);
   U21851 : AOI22_X1 port map( A1 => n24980, A2 => n19997, B1 => n24974, B2 => 
                           n24801, ZN => n23811);
   U21852 : AOI22_X1 port map( A1 => n24980, A2 => n19996, B1 => n24974, B2 => 
                           n24802, ZN => n23793);
   U21853 : AOI22_X1 port map( A1 => n24980, A2 => n19995, B1 => n24974, B2 => 
                           n24803, ZN => n23775);
   U21854 : AOI22_X1 port map( A1 => n24980, A2 => n19994, B1 => n24974, B2 => 
                           n24804, ZN => n23757);
   U21855 : AOI22_X1 port map( A1 => n24980, A2 => n19993, B1 => n24974, B2 => 
                           n24805, ZN => n23739);
   U21856 : AOI22_X1 port map( A1 => n24981, A2 => n19992, B1 => n24975, B2 => 
                           n24806, ZN => n23721);
   U21857 : AOI22_X1 port map( A1 => n24981, A2 => n19991, B1 => n24975, B2 => 
                           n24807, ZN => n23703);
   U21858 : AOI22_X1 port map( A1 => n24981, A2 => n19990, B1 => n24975, B2 => 
                           n24808, ZN => n23685);
   U21859 : AOI22_X1 port map( A1 => n24981, A2 => n19989, B1 => n24975, B2 => 
                           n24809, ZN => n23667);
   U21860 : AOI22_X1 port map( A1 => n24981, A2 => n19988, B1 => n24975, B2 => 
                           n24810, ZN => n23649);
   U21861 : AOI22_X1 port map( A1 => n24981, A2 => n19987, B1 => n24975, B2 => 
                           n24811, ZN => n23631);
   U21862 : AOI22_X1 port map( A1 => n24981, A2 => n19986, B1 => n24975, B2 => 
                           n24812, ZN => n23613);
   U21863 : AOI22_X1 port map( A1 => n24981, A2 => n19985, B1 => n24975, B2 => 
                           n24813, ZN => n23595);
   U21864 : AOI22_X1 port map( A1 => n24981, A2 => n19984, B1 => n24975, B2 => 
                           n24814, ZN => n23577);
   U21865 : AOI22_X1 port map( A1 => n24981, A2 => n19983, B1 => n24975, B2 => 
                           n24815, ZN => n23559);
   U21866 : AOI22_X1 port map( A1 => n24981, A2 => n19982, B1 => n24975, B2 => 
                           n24816, ZN => n23541);
   U21867 : AOI22_X1 port map( A1 => n24981, A2 => n19981, B1 => n24975, B2 => 
                           n24817, ZN => n23523);
   U21868 : AOI22_X1 port map( A1 => n24982, A2 => n19980, B1 => n24976, B2 => 
                           n24818, ZN => n23505);
   U21869 : AOI22_X1 port map( A1 => n24982, A2 => n19979, B1 => n24976, B2 => 
                           n24819, ZN => n23487);
   U21870 : AOI22_X1 port map( A1 => n24982, A2 => n19978, B1 => n24976, B2 => 
                           n24820, ZN => n23469);
   U21871 : AOI22_X1 port map( A1 => n24982, A2 => n19977, B1 => n24976, B2 => 
                           n24821, ZN => n23451);
   U21872 : AOI22_X1 port map( A1 => n24982, A2 => n19976, B1 => n24976, B2 => 
                           n24822, ZN => n23433);
   U21873 : AOI22_X1 port map( A1 => n24982, A2 => n19975, B1 => n24976, B2 => 
                           n24823, ZN => n23415);
   U21874 : AOI22_X1 port map( A1 => n24982, A2 => n19974, B1 => n24976, B2 => 
                           n24824, ZN => n23397);
   U21875 : AOI22_X1 port map( A1 => n24982, A2 => n19973, B1 => n24976, B2 => 
                           n24825, ZN => n23379);
   U21876 : AOI22_X1 port map( A1 => n24982, A2 => n19972, B1 => n24976, B2 => 
                           n24826, ZN => n23361);
   U21877 : AOI22_X1 port map( A1 => n24982, A2 => n19971, B1 => n24976, B2 => 
                           n24827, ZN => n23343);
   U21878 : AOI22_X1 port map( A1 => n24982, A2 => n19970, B1 => n24976, B2 => 
                           n24828, ZN => n23325);
   U21879 : AOI22_X1 port map( A1 => n24982, A2 => n19969, B1 => n24976, B2 => 
                           n24829, ZN => n23307);
   U21880 : AOI22_X1 port map( A1 => n24983, A2 => n19968, B1 => n24977, B2 => 
                           n24830, ZN => n23289);
   U21881 : AOI22_X1 port map( A1 => n24983, A2 => n19967, B1 => n24977, B2 => 
                           n24831, ZN => n23271);
   U21882 : AOI22_X1 port map( A1 => n24983, A2 => n19966, B1 => n24977, B2 => 
                           n24832, ZN => n23253);
   U21883 : AOI22_X1 port map( A1 => n24983, A2 => n19965, B1 => n24977, B2 => 
                           n24833, ZN => n23235);
   U21884 : AOI22_X1 port map( A1 => n24983, A2 => n19964, B1 => n24977, B2 => 
                           n24834, ZN => n23217);
   U21885 : AOI22_X1 port map( A1 => n24983, A2 => n19963, B1 => n24977, B2 => 
                           n24835, ZN => n23199);
   U21886 : AOI22_X1 port map( A1 => n24983, A2 => n19962, B1 => n24977, B2 => 
                           n24836, ZN => n23181);
   U21887 : AOI22_X1 port map( A1 => n24983, A2 => n19961, B1 => n24977, B2 => 
                           n24837, ZN => n23163);
   U21888 : AOI22_X1 port map( A1 => n24983, A2 => n19960, B1 => n24977, B2 => 
                           n24838, ZN => n23145);
   U21889 : AOI22_X1 port map( A1 => n24983, A2 => n19959, B1 => n24977, B2 => 
                           n24839, ZN => n23127);
   U21890 : AOI22_X1 port map( A1 => n24983, A2 => n19958, B1 => n24977, B2 => 
                           n24840, ZN => n23109);
   U21891 : AOI22_X1 port map( A1 => n24983, A2 => n19957, B1 => n24977, B2 => 
                           n24841, ZN => n23091);
   U21892 : AOI22_X1 port map( A1 => n24984, A2 => n19956, B1 => n24978, B2 => 
                           n24842, ZN => n23073);
   U21893 : AOI22_X1 port map( A1 => n24984, A2 => n19955, B1 => n24978, B2 => 
                           n24843, ZN => n23055);
   U21894 : AOI22_X1 port map( A1 => n24984, A2 => n19954, B1 => n24978, B2 => 
                           n24844, ZN => n23037);
   U21895 : AOI22_X1 port map( A1 => n24984, A2 => n19953, B1 => n24978, B2 => 
                           n24845, ZN => n23019);
   U21896 : AOI22_X1 port map( A1 => n24984, A2 => n19952, B1 => n24978, B2 => 
                           n24846, ZN => n23001);
   U21897 : AOI22_X1 port map( A1 => n24984, A2 => n19951, B1 => n24978, B2 => 
                           n24847, ZN => n22983);
   U21898 : AOI22_X1 port map( A1 => n24984, A2 => n19950, B1 => n24978, B2 => 
                           n24848, ZN => n22965);
   U21899 : AOI22_X1 port map( A1 => n24984, A2 => n19949, B1 => n24978, B2 => 
                           n24849, ZN => n22947);
   U21900 : AOI22_X1 port map( A1 => n24984, A2 => n19948, B1 => n24978, B2 => 
                           n24850, ZN => n22929);
   U21901 : AOI22_X1 port map( A1 => n24984, A2 => n19947, B1 => n24978, B2 => 
                           n24851, ZN => n22911);
   U21902 : AOI22_X1 port map( A1 => n24984, A2 => n19946, B1 => n24978, B2 => 
                           n24852, ZN => n22893);
   U21903 : AOI22_X1 port map( A1 => n24984, A2 => n19945, B1 => n24978, B2 => 
                           n24853, ZN => n22875);
   U21904 : AOI22_X1 port map( A1 => n24985, A2 => n19944, B1 => n24979, B2 => 
                           n24474, ZN => n22857);
   U21905 : AOI22_X1 port map( A1 => n24985, A2 => n19943, B1 => n24979, B2 => 
                           n24475, ZN => n22839);
   U21906 : AOI22_X1 port map( A1 => n24985, A2 => n19942, B1 => n24979, B2 => 
                           n24476, ZN => n22821);
   U21907 : AOI22_X1 port map( A1 => n25178, A2 => n20004, B1 => n25172, B2 => 
                           n24794, ZN => n22752);
   U21908 : AOI22_X1 port map( A1 => n25178, A2 => n20003, B1 => n25172, B2 => 
                           n24795, ZN => n22722);
   U21909 : AOI22_X1 port map( A1 => n25178, A2 => n20002, B1 => n25172, B2 => 
                           n24796, ZN => n22704);
   U21910 : AOI22_X1 port map( A1 => n25178, A2 => n20001, B1 => n25172, B2 => 
                           n24797, ZN => n22686);
   U21911 : AOI22_X1 port map( A1 => n25178, A2 => n20000, B1 => n25172, B2 => 
                           n24798, ZN => n22668);
   U21912 : AOI22_X1 port map( A1 => n25178, A2 => n19999, B1 => n25172, B2 => 
                           n24799, ZN => n22650);
   U21913 : AOI22_X1 port map( A1 => n25178, A2 => n19998, B1 => n25172, B2 => 
                           n24800, ZN => n22632);
   U21914 : AOI22_X1 port map( A1 => n25178, A2 => n19997, B1 => n25172, B2 => 
                           n24801, ZN => n22614);
   U21915 : AOI22_X1 port map( A1 => n25178, A2 => n19996, B1 => n25172, B2 => 
                           n24802, ZN => n22596);
   U21916 : AOI22_X1 port map( A1 => n25178, A2 => n19995, B1 => n25172, B2 => 
                           n24803, ZN => n22578);
   U21917 : AOI22_X1 port map( A1 => n25178, A2 => n19994, B1 => n25172, B2 => 
                           n24804, ZN => n22560);
   U21918 : AOI22_X1 port map( A1 => n25178, A2 => n19993, B1 => n25172, B2 => 
                           n24805, ZN => n22542);
   U21919 : AOI22_X1 port map( A1 => n25179, A2 => n19992, B1 => n25173, B2 => 
                           n24806, ZN => n22524);
   U21920 : AOI22_X1 port map( A1 => n25179, A2 => n19991, B1 => n25173, B2 => 
                           n24807, ZN => n22506);
   U21921 : AOI22_X1 port map( A1 => n25179, A2 => n19990, B1 => n25173, B2 => 
                           n24808, ZN => n22488);
   U21922 : AOI22_X1 port map( A1 => n25179, A2 => n19989, B1 => n25173, B2 => 
                           n24809, ZN => n22470);
   U21923 : AOI22_X1 port map( A1 => n25179, A2 => n19988, B1 => n25173, B2 => 
                           n24810, ZN => n22452);
   U21924 : AOI22_X1 port map( A1 => n25179, A2 => n19987, B1 => n25173, B2 => 
                           n24811, ZN => n22434);
   U21925 : AOI22_X1 port map( A1 => n25179, A2 => n19986, B1 => n25173, B2 => 
                           n24812, ZN => n22416);
   U21926 : AOI22_X1 port map( A1 => n25179, A2 => n19985, B1 => n25173, B2 => 
                           n24813, ZN => n22398);
   U21927 : AOI22_X1 port map( A1 => n25179, A2 => n19984, B1 => n25173, B2 => 
                           n24814, ZN => n22380);
   U21928 : AOI22_X1 port map( A1 => n25179, A2 => n19983, B1 => n25173, B2 => 
                           n24815, ZN => n22362);
   U21929 : AOI22_X1 port map( A1 => n25179, A2 => n19982, B1 => n25173, B2 => 
                           n24816, ZN => n22344);
   U21930 : AOI22_X1 port map( A1 => n25179, A2 => n19981, B1 => n25173, B2 => 
                           n24817, ZN => n22326);
   U21931 : AOI22_X1 port map( A1 => n25180, A2 => n19980, B1 => n25174, B2 => 
                           n24818, ZN => n22308);
   U21932 : AOI22_X1 port map( A1 => n25180, A2 => n19979, B1 => n25174, B2 => 
                           n24819, ZN => n22290);
   U21933 : AOI22_X1 port map( A1 => n25180, A2 => n19978, B1 => n25174, B2 => 
                           n24820, ZN => n22272);
   U21934 : AOI22_X1 port map( A1 => n25180, A2 => n19977, B1 => n25174, B2 => 
                           n24821, ZN => n22254);
   U21935 : AOI22_X1 port map( A1 => n25180, A2 => n19976, B1 => n25174, B2 => 
                           n24822, ZN => n22236);
   U21936 : AOI22_X1 port map( A1 => n25180, A2 => n19975, B1 => n25174, B2 => 
                           n24823, ZN => n22218);
   U21937 : AOI22_X1 port map( A1 => n25180, A2 => n19974, B1 => n25174, B2 => 
                           n24824, ZN => n22200);
   U21938 : AOI22_X1 port map( A1 => n25180, A2 => n19973, B1 => n25174, B2 => 
                           n24825, ZN => n22182);
   U21939 : AOI22_X1 port map( A1 => n25180, A2 => n19972, B1 => n25174, B2 => 
                           n24826, ZN => n22164);
   U21940 : AOI22_X1 port map( A1 => n25180, A2 => n19971, B1 => n25174, B2 => 
                           n24827, ZN => n22146);
   U21941 : AOI22_X1 port map( A1 => n25180, A2 => n19970, B1 => n25174, B2 => 
                           n24828, ZN => n22128);
   U21942 : AOI22_X1 port map( A1 => n25180, A2 => n19969, B1 => n25174, B2 => 
                           n24829, ZN => n22110);
   U21943 : AOI22_X1 port map( A1 => n25181, A2 => n19968, B1 => n25175, B2 => 
                           n24830, ZN => n22092);
   U21944 : AOI22_X1 port map( A1 => n25181, A2 => n19967, B1 => n25175, B2 => 
                           n24831, ZN => n22074);
   U21945 : AOI22_X1 port map( A1 => n25181, A2 => n19966, B1 => n25175, B2 => 
                           n24832, ZN => n22056);
   U21946 : AOI22_X1 port map( A1 => n25181, A2 => n19965, B1 => n25175, B2 => 
                           n24833, ZN => n22038);
   U21947 : AOI22_X1 port map( A1 => n25181, A2 => n19964, B1 => n25175, B2 => 
                           n24834, ZN => n22020);
   U21948 : AOI22_X1 port map( A1 => n25181, A2 => n19963, B1 => n25175, B2 => 
                           n24835, ZN => n22002);
   U21949 : AOI22_X1 port map( A1 => n25181, A2 => n19962, B1 => n25175, B2 => 
                           n24836, ZN => n21984);
   U21950 : AOI22_X1 port map( A1 => n25181, A2 => n19961, B1 => n25175, B2 => 
                           n24837, ZN => n21966);
   U21951 : AOI22_X1 port map( A1 => n25181, A2 => n19960, B1 => n25175, B2 => 
                           n24838, ZN => n21948);
   U21952 : AOI22_X1 port map( A1 => n25181, A2 => n19959, B1 => n25175, B2 => 
                           n24839, ZN => n21930);
   U21953 : AOI22_X1 port map( A1 => n25181, A2 => n19958, B1 => n25175, B2 => 
                           n24840, ZN => n21912);
   U21954 : AOI22_X1 port map( A1 => n25181, A2 => n19957, B1 => n25175, B2 => 
                           n24841, ZN => n21894);
   U21955 : AOI22_X1 port map( A1 => n25182, A2 => n19956, B1 => n25176, B2 => 
                           n24842, ZN => n21876);
   U21956 : AOI22_X1 port map( A1 => n25182, A2 => n19955, B1 => n25176, B2 => 
                           n24843, ZN => n21858);
   U21957 : AOI22_X1 port map( A1 => n25182, A2 => n19954, B1 => n25176, B2 => 
                           n24844, ZN => n21840);
   U21958 : AOI22_X1 port map( A1 => n25182, A2 => n19953, B1 => n25176, B2 => 
                           n24845, ZN => n21822);
   U21959 : AOI22_X1 port map( A1 => n25182, A2 => n19952, B1 => n25176, B2 => 
                           n24846, ZN => n21804);
   U21960 : AOI22_X1 port map( A1 => n25182, A2 => n19951, B1 => n25176, B2 => 
                           n24847, ZN => n21786);
   U21961 : AOI22_X1 port map( A1 => n25182, A2 => n19950, B1 => n25176, B2 => 
                           n24848, ZN => n21768);
   U21962 : AOI22_X1 port map( A1 => n25182, A2 => n19949, B1 => n25176, B2 => 
                           n24849, ZN => n21750);
   U21963 : AOI22_X1 port map( A1 => n25182, A2 => n19948, B1 => n25176, B2 => 
                           n24850, ZN => n21732);
   U21964 : AOI22_X1 port map( A1 => n25182, A2 => n19947, B1 => n25176, B2 => 
                           n24851, ZN => n21714);
   U21965 : AOI22_X1 port map( A1 => n25182, A2 => n19946, B1 => n25176, B2 => 
                           n24852, ZN => n21696);
   U21966 : AOI22_X1 port map( A1 => n25182, A2 => n19945, B1 => n25176, B2 => 
                           n24853, ZN => n21678);
   U21967 : AOI22_X1 port map( A1 => n25183, A2 => n19944, B1 => n25177, B2 => 
                           n24474, ZN => n21660);
   U21968 : AOI22_X1 port map( A1 => n25183, A2 => n19943, B1 => n25177, B2 => 
                           n24475, ZN => n21642);
   U21969 : AOI22_X1 port map( A1 => n25183, A2 => n19942, B1 => n25177, B2 => 
                           n24476, ZN => n21624);
   U21970 : AOI22_X1 port map( A1 => n25183, A2 => n19941, B1 => n25177, B2 => 
                           n24477, ZN => n21604);
   U21971 : OAI221_X1 port map( B1 => n21285, B2 => n25118, C1 => n19621, C2 =>
                           n25112, A => n23936, ZN => n23923);
   U21972 : AOI22_X1 port map( A1 => n25106, A2 => n24854, B1 => n25100, B2 => 
                           n20068, ZN => n23936);
   U21973 : OAI221_X1 port map( B1 => n21221, B2 => n25064, C1 => n20197, C2 =>
                           n25058, A => n23945, ZN => n23944);
   U21974 : AOI22_X1 port map( A1 => n25052, A2 => n24087, B1 => n25046, B2 => 
                           OUT2_0_port, ZN => n23945);
   U21975 : OAI221_X1 port map( B1 => n21284, B2 => n25118, C1 => n19620, C2 =>
                           n25112, A => n23910, ZN => n23905);
   U21976 : AOI22_X1 port map( A1 => n25106, A2 => n24855, B1 => n25100, B2 => 
                           n20067, ZN => n23910);
   U21977 : OAI221_X1 port map( B1 => n21220, B2 => n25064, C1 => n20196, C2 =>
                           n25058, A => n23916, ZN => n23915);
   U21978 : AOI22_X1 port map( A1 => n25052, A2 => n24089, B1 => n25051, B2 => 
                           OUT2_1_port, ZN => n23916);
   U21979 : OAI221_X1 port map( B1 => n21283, B2 => n25118, C1 => n19619, C2 =>
                           n25112, A => n23892, ZN => n23887);
   U21980 : AOI22_X1 port map( A1 => n25106, A2 => n24856, B1 => n25100, B2 => 
                           n20066, ZN => n23892);
   U21981 : OAI221_X1 port map( B1 => n21219, B2 => n25064, C1 => n20195, C2 =>
                           n25058, A => n23898, ZN => n23897);
   U21982 : AOI22_X1 port map( A1 => n25052, A2 => n24091, B1 => n25051, B2 => 
                           OUT2_2_port, ZN => n23898);
   U21983 : OAI221_X1 port map( B1 => n21282, B2 => n25118, C1 => n19618, C2 =>
                           n25112, A => n23874, ZN => n23869);
   U21984 : AOI22_X1 port map( A1 => n25106, A2 => n24857, B1 => n25100, B2 => 
                           n20065, ZN => n23874);
   U21985 : OAI221_X1 port map( B1 => n21218, B2 => n25064, C1 => n20194, C2 =>
                           n25058, A => n23880, ZN => n23879);
   U21986 : AOI22_X1 port map( A1 => n25052, A2 => n24093, B1 => n25051, B2 => 
                           OUT2_3_port, ZN => n23880);
   U21987 : OAI221_X1 port map( B1 => n21281, B2 => n25118, C1 => n19617, C2 =>
                           n25112, A => n23856, ZN => n23851);
   U21988 : AOI22_X1 port map( A1 => n25106, A2 => n24858, B1 => n25100, B2 => 
                           n20064, ZN => n23856);
   U21989 : OAI221_X1 port map( B1 => n21217, B2 => n25064, C1 => n20193, C2 =>
                           n25058, A => n23862, ZN => n23861);
   U21990 : AOI22_X1 port map( A1 => n25052, A2 => n24095, B1 => n25050, B2 => 
                           OUT2_4_port, ZN => n23862);
   U21991 : OAI221_X1 port map( B1 => n21280, B2 => n25118, C1 => n19616, C2 =>
                           n25112, A => n23838, ZN => n23833);
   U21992 : AOI22_X1 port map( A1 => n25106, A2 => n24859, B1 => n25100, B2 => 
                           n20063, ZN => n23838);
   U21993 : OAI221_X1 port map( B1 => n21216, B2 => n25064, C1 => n20192, C2 =>
                           n25058, A => n23844, ZN => n23843);
   U21994 : AOI22_X1 port map( A1 => n25052, A2 => n24097, B1 => n25050, B2 => 
                           OUT2_5_port, ZN => n23844);
   U21995 : OAI221_X1 port map( B1 => n21279, B2 => n25118, C1 => n19615, C2 =>
                           n25112, A => n23820, ZN => n23815);
   U21996 : AOI22_X1 port map( A1 => n25106, A2 => n24860, B1 => n25100, B2 => 
                           n20062, ZN => n23820);
   U21997 : OAI221_X1 port map( B1 => n21215, B2 => n25064, C1 => n20191, C2 =>
                           n25058, A => n23826, ZN => n23825);
   U21998 : AOI22_X1 port map( A1 => n25052, A2 => n24099, B1 => n25050, B2 => 
                           OUT2_6_port, ZN => n23826);
   U21999 : OAI221_X1 port map( B1 => n21278, B2 => n25118, C1 => n19614, C2 =>
                           n25112, A => n23802, ZN => n23797);
   U22000 : AOI22_X1 port map( A1 => n25106, A2 => n24861, B1 => n25100, B2 => 
                           n20061, ZN => n23802);
   U22001 : OAI221_X1 port map( B1 => n21214, B2 => n25064, C1 => n20190, C2 =>
                           n25058, A => n23808, ZN => n23807);
   U22002 : AOI22_X1 port map( A1 => n25052, A2 => n24101, B1 => n25050, B2 => 
                           OUT2_7_port, ZN => n23808);
   U22003 : OAI221_X1 port map( B1 => n21277, B2 => n25118, C1 => n19613, C2 =>
                           n25112, A => n23784, ZN => n23779);
   U22004 : AOI22_X1 port map( A1 => n25106, A2 => n24862, B1 => n25100, B2 => 
                           n20060, ZN => n23784);
   U22005 : OAI221_X1 port map( B1 => n21213, B2 => n25064, C1 => n20189, C2 =>
                           n25058, A => n23790, ZN => n23789);
   U22006 : AOI22_X1 port map( A1 => n25052, A2 => n24103, B1 => n25050, B2 => 
                           OUT2_8_port, ZN => n23790);
   U22007 : OAI221_X1 port map( B1 => n21276, B2 => n25118, C1 => n19612, C2 =>
                           n25112, A => n23766, ZN => n23761);
   U22008 : AOI22_X1 port map( A1 => n25106, A2 => n24863, B1 => n25100, B2 => 
                           n20059, ZN => n23766);
   U22009 : OAI221_X1 port map( B1 => n21212, B2 => n25064, C1 => n20188, C2 =>
                           n25058, A => n23772, ZN => n23771);
   U22010 : AOI22_X1 port map( A1 => n25052, A2 => n24105, B1 => n25050, B2 => 
                           OUT2_9_port, ZN => n23772);
   U22011 : OAI221_X1 port map( B1 => n21275, B2 => n25118, C1 => n19611, C2 =>
                           n25112, A => n23748, ZN => n23743);
   U22012 : AOI22_X1 port map( A1 => n25106, A2 => n24864, B1 => n25100, B2 => 
                           n20058, ZN => n23748);
   U22013 : OAI221_X1 port map( B1 => n21211, B2 => n25064, C1 => n20187, C2 =>
                           n25058, A => n23754, ZN => n23753);
   U22014 : AOI22_X1 port map( A1 => n25052, A2 => n24107, B1 => n25050, B2 => 
                           OUT2_10_port, ZN => n23754);
   U22015 : OAI221_X1 port map( B1 => n21274, B2 => n25118, C1 => n19610, C2 =>
                           n25112, A => n23730, ZN => n23725);
   U22016 : AOI22_X1 port map( A1 => n25106, A2 => n24865, B1 => n25100, B2 => 
                           n20057, ZN => n23730);
   U22017 : OAI221_X1 port map( B1 => n21210, B2 => n25064, C1 => n20186, C2 =>
                           n25058, A => n23736, ZN => n23735);
   U22018 : AOI22_X1 port map( A1 => n25052, A2 => n24109, B1 => n25050, B2 => 
                           OUT2_11_port, ZN => n23736);
   U22019 : OAI221_X1 port map( B1 => n21273, B2 => n25119, C1 => n19609, C2 =>
                           n25113, A => n23712, ZN => n23707);
   U22020 : AOI22_X1 port map( A1 => n25107, A2 => n24866, B1 => n25101, B2 => 
                           n20056, ZN => n23712);
   U22021 : OAI221_X1 port map( B1 => n21209, B2 => n25065, C1 => n20185, C2 =>
                           n25059, A => n23718, ZN => n23717);
   U22022 : AOI22_X1 port map( A1 => n25053, A2 => n24111, B1 => n25050, B2 => 
                           OUT2_12_port, ZN => n23718);
   U22023 : OAI221_X1 port map( B1 => n21272, B2 => n25119, C1 => n19608, C2 =>
                           n25113, A => n23694, ZN => n23689);
   U22024 : AOI22_X1 port map( A1 => n25107, A2 => n24867, B1 => n25101, B2 => 
                           n20055, ZN => n23694);
   U22025 : OAI221_X1 port map( B1 => n21208, B2 => n25065, C1 => n20184, C2 =>
                           n25059, A => n23700, ZN => n23699);
   U22026 : AOI22_X1 port map( A1 => n25053, A2 => n24113, B1 => n25050, B2 => 
                           OUT2_13_port, ZN => n23700);
   U22027 : OAI221_X1 port map( B1 => n21271, B2 => n25119, C1 => n19607, C2 =>
                           n25113, A => n23676, ZN => n23671);
   U22028 : AOI22_X1 port map( A1 => n25107, A2 => n24868, B1 => n25101, B2 => 
                           n20054, ZN => n23676);
   U22029 : OAI221_X1 port map( B1 => n21207, B2 => n25065, C1 => n20183, C2 =>
                           n25059, A => n23682, ZN => n23681);
   U22030 : AOI22_X1 port map( A1 => n25053, A2 => n24115, B1 => n25050, B2 => 
                           OUT2_14_port, ZN => n23682);
   U22031 : OAI221_X1 port map( B1 => n21270, B2 => n25119, C1 => n19606, C2 =>
                           n25113, A => n23658, ZN => n23653);
   U22032 : AOI22_X1 port map( A1 => n25107, A2 => n24869, B1 => n25101, B2 => 
                           n20053, ZN => n23658);
   U22033 : OAI221_X1 port map( B1 => n21206, B2 => n25065, C1 => n20182, C2 =>
                           n25059, A => n23664, ZN => n23663);
   U22034 : AOI22_X1 port map( A1 => n25053, A2 => n24117, B1 => n25050, B2 => 
                           OUT2_15_port, ZN => n23664);
   U22035 : OAI221_X1 port map( B1 => n21269, B2 => n25119, C1 => n19605, C2 =>
                           n25113, A => n23640, ZN => n23635);
   U22036 : AOI22_X1 port map( A1 => n25107, A2 => n24870, B1 => n25101, B2 => 
                           n20052, ZN => n23640);
   U22037 : OAI221_X1 port map( B1 => n21205, B2 => n25065, C1 => n20181, C2 =>
                           n25059, A => n23646, ZN => n23645);
   U22038 : AOI22_X1 port map( A1 => n25053, A2 => n24119, B1 => n25050, B2 => 
                           OUT2_16_port, ZN => n23646);
   U22039 : OAI221_X1 port map( B1 => n21268, B2 => n25119, C1 => n19604, C2 =>
                           n25113, A => n23622, ZN => n23617);
   U22040 : AOI22_X1 port map( A1 => n25107, A2 => n24871, B1 => n25101, B2 => 
                           n20051, ZN => n23622);
   U22041 : OAI221_X1 port map( B1 => n21204, B2 => n25065, C1 => n20180, C2 =>
                           n25059, A => n23628, ZN => n23627);
   U22042 : AOI22_X1 port map( A1 => n25053, A2 => n24121, B1 => n25049, B2 => 
                           OUT2_17_port, ZN => n23628);
   U22043 : OAI221_X1 port map( B1 => n21267, B2 => n25119, C1 => n19603, C2 =>
                           n25113, A => n23604, ZN => n23599);
   U22044 : AOI22_X1 port map( A1 => n25107, A2 => n24872, B1 => n25101, B2 => 
                           n20050, ZN => n23604);
   U22045 : OAI221_X1 port map( B1 => n21203, B2 => n25065, C1 => n20179, C2 =>
                           n25059, A => n23610, ZN => n23609);
   U22046 : AOI22_X1 port map( A1 => n25053, A2 => n24123, B1 => n25049, B2 => 
                           OUT2_18_port, ZN => n23610);
   U22047 : OAI221_X1 port map( B1 => n21266, B2 => n25119, C1 => n19602, C2 =>
                           n25113, A => n23586, ZN => n23581);
   U22048 : AOI22_X1 port map( A1 => n25107, A2 => n24873, B1 => n25101, B2 => 
                           n20049, ZN => n23586);
   U22049 : OAI221_X1 port map( B1 => n21202, B2 => n25065, C1 => n20178, C2 =>
                           n25059, A => n23592, ZN => n23591);
   U22050 : AOI22_X1 port map( A1 => n25053, A2 => n24125, B1 => n25049, B2 => 
                           OUT2_19_port, ZN => n23592);
   U22051 : OAI221_X1 port map( B1 => n21265, B2 => n25119, C1 => n19601, C2 =>
                           n25113, A => n23568, ZN => n23563);
   U22052 : AOI22_X1 port map( A1 => n25107, A2 => n24874, B1 => n25101, B2 => 
                           n20048, ZN => n23568);
   U22053 : OAI221_X1 port map( B1 => n21201, B2 => n25065, C1 => n20177, C2 =>
                           n25059, A => n23574, ZN => n23573);
   U22054 : AOI22_X1 port map( A1 => n25053, A2 => n24127, B1 => n25049, B2 => 
                           OUT2_20_port, ZN => n23574);
   U22055 : OAI221_X1 port map( B1 => n21264, B2 => n25119, C1 => n19600, C2 =>
                           n25113, A => n23550, ZN => n23545);
   U22056 : AOI22_X1 port map( A1 => n25107, A2 => n24875, B1 => n25101, B2 => 
                           n20047, ZN => n23550);
   U22057 : OAI221_X1 port map( B1 => n21200, B2 => n25065, C1 => n20176, C2 =>
                           n25059, A => n23556, ZN => n23555);
   U22058 : AOI22_X1 port map( A1 => n25053, A2 => n24129, B1 => n25049, B2 => 
                           OUT2_21_port, ZN => n23556);
   U22059 : OAI221_X1 port map( B1 => n21263, B2 => n25119, C1 => n19599, C2 =>
                           n25113, A => n23532, ZN => n23527);
   U22060 : AOI22_X1 port map( A1 => n25107, A2 => n24876, B1 => n25101, B2 => 
                           n20046, ZN => n23532);
   U22061 : OAI221_X1 port map( B1 => n21199, B2 => n25065, C1 => n20175, C2 =>
                           n25059, A => n23538, ZN => n23537);
   U22062 : AOI22_X1 port map( A1 => n25053, A2 => n24131, B1 => n25049, B2 => 
                           OUT2_22_port, ZN => n23538);
   U22063 : OAI221_X1 port map( B1 => n21262, B2 => n25119, C1 => n19598, C2 =>
                           n25113, A => n23514, ZN => n23509);
   U22064 : AOI22_X1 port map( A1 => n25107, A2 => n24877, B1 => n25101, B2 => 
                           n20045, ZN => n23514);
   U22065 : OAI221_X1 port map( B1 => n21198, B2 => n25065, C1 => n20174, C2 =>
                           n25059, A => n23520, ZN => n23519);
   U22066 : AOI22_X1 port map( A1 => n25053, A2 => n24133, B1 => n25049, B2 => 
                           OUT2_23_port, ZN => n23520);
   U22067 : OAI221_X1 port map( B1 => n21261, B2 => n25120, C1 => n19597, C2 =>
                           n25114, A => n23496, ZN => n23491);
   U22068 : AOI22_X1 port map( A1 => n25108, A2 => n24878, B1 => n25102, B2 => 
                           n20044, ZN => n23496);
   U22069 : OAI221_X1 port map( B1 => n21197, B2 => n25066, C1 => n20173, C2 =>
                           n25060, A => n23502, ZN => n23501);
   U22070 : AOI22_X1 port map( A1 => n25054, A2 => n24135, B1 => n25049, B2 => 
                           OUT2_24_port, ZN => n23502);
   U22071 : OAI221_X1 port map( B1 => n21260, B2 => n25120, C1 => n19596, C2 =>
                           n25114, A => n23478, ZN => n23473);
   U22072 : AOI22_X1 port map( A1 => n25108, A2 => n24879, B1 => n25102, B2 => 
                           n20043, ZN => n23478);
   U22073 : OAI221_X1 port map( B1 => n21196, B2 => n25066, C1 => n20172, C2 =>
                           n25060, A => n23484, ZN => n23483);
   U22074 : AOI22_X1 port map( A1 => n25054, A2 => n24137, B1 => n25049, B2 => 
                           OUT2_25_port, ZN => n23484);
   U22075 : OAI221_X1 port map( B1 => n21259, B2 => n25120, C1 => n19595, C2 =>
                           n25114, A => n23460, ZN => n23455);
   U22076 : AOI22_X1 port map( A1 => n25108, A2 => n24880, B1 => n25102, B2 => 
                           n20042, ZN => n23460);
   U22077 : OAI221_X1 port map( B1 => n21195, B2 => n25066, C1 => n20171, C2 =>
                           n25060, A => n23466, ZN => n23465);
   U22078 : AOI22_X1 port map( A1 => n25054, A2 => n24139, B1 => n25049, B2 => 
                           OUT2_26_port, ZN => n23466);
   U22079 : OAI221_X1 port map( B1 => n21258, B2 => n25120, C1 => n19594, C2 =>
                           n25114, A => n23442, ZN => n23437);
   U22080 : AOI22_X1 port map( A1 => n25108, A2 => n24881, B1 => n25102, B2 => 
                           n20041, ZN => n23442);
   U22081 : OAI221_X1 port map( B1 => n21194, B2 => n25066, C1 => n20170, C2 =>
                           n25060, A => n23448, ZN => n23447);
   U22082 : AOI22_X1 port map( A1 => n25054, A2 => n24141, B1 => n25049, B2 => 
                           OUT2_27_port, ZN => n23448);
   U22083 : OAI221_X1 port map( B1 => n21257, B2 => n25120, C1 => n19593, C2 =>
                           n25114, A => n23424, ZN => n23419);
   U22084 : AOI22_X1 port map( A1 => n25108, A2 => n24882, B1 => n25102, B2 => 
                           n20040, ZN => n23424);
   U22085 : OAI221_X1 port map( B1 => n21193, B2 => n25066, C1 => n20169, C2 =>
                           n25060, A => n23430, ZN => n23429);
   U22086 : AOI22_X1 port map( A1 => n25054, A2 => n24143, B1 => n25049, B2 => 
                           OUT2_28_port, ZN => n23430);
   U22087 : OAI221_X1 port map( B1 => n21256, B2 => n25120, C1 => n19592, C2 =>
                           n25114, A => n23406, ZN => n23401);
   U22088 : AOI22_X1 port map( A1 => n25108, A2 => n24883, B1 => n25102, B2 => 
                           n20039, ZN => n23406);
   U22089 : OAI221_X1 port map( B1 => n21192, B2 => n25066, C1 => n20168, C2 =>
                           n25060, A => n23412, ZN => n23411);
   U22090 : AOI22_X1 port map( A1 => n25054, A2 => n24145, B1 => n25049, B2 => 
                           OUT2_29_port, ZN => n23412);
   U22091 : OAI221_X1 port map( B1 => n21255, B2 => n25120, C1 => n19591, C2 =>
                           n25114, A => n23388, ZN => n23383);
   U22092 : AOI22_X1 port map( A1 => n25108, A2 => n24884, B1 => n25102, B2 => 
                           n20038, ZN => n23388);
   U22093 : OAI221_X1 port map( B1 => n21191, B2 => n25066, C1 => n20167, C2 =>
                           n25060, A => n23394, ZN => n23393);
   U22094 : AOI22_X1 port map( A1 => n25054, A2 => n24147, B1 => n25048, B2 => 
                           OUT2_30_port, ZN => n23394);
   U22095 : OAI221_X1 port map( B1 => n21254, B2 => n25120, C1 => n19590, C2 =>
                           n25114, A => n23370, ZN => n23365);
   U22096 : AOI22_X1 port map( A1 => n25108, A2 => n24885, B1 => n25102, B2 => 
                           n20037, ZN => n23370);
   U22097 : OAI221_X1 port map( B1 => n21190, B2 => n25066, C1 => n20166, C2 =>
                           n25060, A => n23376, ZN => n23375);
   U22098 : AOI22_X1 port map( A1 => n25054, A2 => n24149, B1 => n25048, B2 => 
                           OUT2_31_port, ZN => n23376);
   U22099 : OAI221_X1 port map( B1 => n21253, B2 => n25120, C1 => n19589, C2 =>
                           n25114, A => n23352, ZN => n23347);
   U22100 : AOI22_X1 port map( A1 => n25108, A2 => n24886, B1 => n25102, B2 => 
                           n20036, ZN => n23352);
   U22101 : OAI221_X1 port map( B1 => n21189, B2 => n25066, C1 => n20165, C2 =>
                           n25060, A => n23358, ZN => n23357);
   U22102 : AOI22_X1 port map( A1 => n25054, A2 => n24151, B1 => n25048, B2 => 
                           OUT2_32_port, ZN => n23358);
   U22103 : OAI221_X1 port map( B1 => n21252, B2 => n25120, C1 => n19588, C2 =>
                           n25114, A => n23334, ZN => n23329);
   U22104 : AOI22_X1 port map( A1 => n25108, A2 => n24887, B1 => n25102, B2 => 
                           n20035, ZN => n23334);
   U22105 : OAI221_X1 port map( B1 => n21188, B2 => n25066, C1 => n20164, C2 =>
                           n25060, A => n23340, ZN => n23339);
   U22106 : AOI22_X1 port map( A1 => n25054, A2 => n24153, B1 => n25048, B2 => 
                           OUT2_33_port, ZN => n23340);
   U22107 : OAI221_X1 port map( B1 => n21251, B2 => n25120, C1 => n19587, C2 =>
                           n25114, A => n23316, ZN => n23311);
   U22108 : AOI22_X1 port map( A1 => n25108, A2 => n24888, B1 => n25102, B2 => 
                           n20034, ZN => n23316);
   U22109 : OAI221_X1 port map( B1 => n21187, B2 => n25066, C1 => n20163, C2 =>
                           n25060, A => n23322, ZN => n23321);
   U22110 : AOI22_X1 port map( A1 => n25054, A2 => n24155, B1 => n25048, B2 => 
                           OUT2_34_port, ZN => n23322);
   U22111 : OAI221_X1 port map( B1 => n21250, B2 => n25120, C1 => n19586, C2 =>
                           n25114, A => n23298, ZN => n23293);
   U22112 : AOI22_X1 port map( A1 => n25108, A2 => n24889, B1 => n25102, B2 => 
                           n20033, ZN => n23298);
   U22113 : OAI221_X1 port map( B1 => n21186, B2 => n25066, C1 => n20162, C2 =>
                           n25060, A => n23304, ZN => n23303);
   U22114 : AOI22_X1 port map( A1 => n25054, A2 => n24157, B1 => n25048, B2 => 
                           OUT2_35_port, ZN => n23304);
   U22115 : OAI221_X1 port map( B1 => n21249, B2 => n25121, C1 => n19585, C2 =>
                           n25115, A => n23280, ZN => n23275);
   U22116 : AOI22_X1 port map( A1 => n25109, A2 => n24890, B1 => n25103, B2 => 
                           n20032, ZN => n23280);
   U22117 : OAI221_X1 port map( B1 => n21185, B2 => n25067, C1 => n20161, C2 =>
                           n25061, A => n23286, ZN => n23285);
   U22118 : AOI22_X1 port map( A1 => n25055, A2 => n24159, B1 => n25048, B2 => 
                           OUT2_36_port, ZN => n23286);
   U22119 : OAI221_X1 port map( B1 => n21248, B2 => n25121, C1 => n19584, C2 =>
                           n25115, A => n23262, ZN => n23257);
   U22120 : AOI22_X1 port map( A1 => n25109, A2 => n24891, B1 => n25103, B2 => 
                           n20031, ZN => n23262);
   U22121 : OAI221_X1 port map( B1 => n21184, B2 => n25067, C1 => n20160, C2 =>
                           n25061, A => n23268, ZN => n23267);
   U22122 : AOI22_X1 port map( A1 => n25055, A2 => n24161, B1 => n25048, B2 => 
                           OUT2_37_port, ZN => n23268);
   U22123 : OAI221_X1 port map( B1 => n21247, B2 => n25121, C1 => n19583, C2 =>
                           n25115, A => n23244, ZN => n23239);
   U22124 : AOI22_X1 port map( A1 => n25109, A2 => n24892, B1 => n25103, B2 => 
                           n20030, ZN => n23244);
   U22125 : OAI221_X1 port map( B1 => n21183, B2 => n25067, C1 => n20159, C2 =>
                           n25061, A => n23250, ZN => n23249);
   U22126 : AOI22_X1 port map( A1 => n25055, A2 => n24163, B1 => n25048, B2 => 
                           OUT2_38_port, ZN => n23250);
   U22127 : OAI221_X1 port map( B1 => n21246, B2 => n25121, C1 => n19582, C2 =>
                           n25115, A => n23226, ZN => n23221);
   U22128 : AOI22_X1 port map( A1 => n25109, A2 => n24893, B1 => n25103, B2 => 
                           n20029, ZN => n23226);
   U22129 : OAI221_X1 port map( B1 => n21182, B2 => n25067, C1 => n20158, C2 =>
                           n25061, A => n23232, ZN => n23231);
   U22130 : AOI22_X1 port map( A1 => n25055, A2 => n24165, B1 => n25048, B2 => 
                           OUT2_39_port, ZN => n23232);
   U22131 : OAI221_X1 port map( B1 => n21245, B2 => n25121, C1 => n19581, C2 =>
                           n25115, A => n23208, ZN => n23203);
   U22132 : AOI22_X1 port map( A1 => n25109, A2 => n24894, B1 => n25103, B2 => 
                           n20028, ZN => n23208);
   U22133 : OAI221_X1 port map( B1 => n21181, B2 => n25067, C1 => n20157, C2 =>
                           n25061, A => n23214, ZN => n23213);
   U22134 : AOI22_X1 port map( A1 => n25055, A2 => n24167, B1 => n25048, B2 => 
                           OUT2_40_port, ZN => n23214);
   U22135 : OAI221_X1 port map( B1 => n21244, B2 => n25121, C1 => n19580, C2 =>
                           n25115, A => n23190, ZN => n23185);
   U22136 : AOI22_X1 port map( A1 => n25109, A2 => n24895, B1 => n25103, B2 => 
                           n20027, ZN => n23190);
   U22137 : OAI221_X1 port map( B1 => n21180, B2 => n25067, C1 => n20156, C2 =>
                           n25061, A => n23196, ZN => n23195);
   U22138 : AOI22_X1 port map( A1 => n25055, A2 => n24169, B1 => n25048, B2 => 
                           OUT2_41_port, ZN => n23196);
   U22139 : OAI221_X1 port map( B1 => n21243, B2 => n25121, C1 => n19579, C2 =>
                           n25115, A => n23172, ZN => n23167);
   U22140 : AOI22_X1 port map( A1 => n25109, A2 => n24896, B1 => n25103, B2 => 
                           n20026, ZN => n23172);
   U22141 : OAI221_X1 port map( B1 => n21179, B2 => n25067, C1 => n20155, C2 =>
                           n25061, A => n23178, ZN => n23177);
   U22142 : AOI22_X1 port map( A1 => n25055, A2 => n24171, B1 => n25047, B2 => 
                           OUT2_42_port, ZN => n23178);
   U22143 : OAI221_X1 port map( B1 => n21242, B2 => n25121, C1 => n19578, C2 =>
                           n25115, A => n23154, ZN => n23149);
   U22144 : AOI22_X1 port map( A1 => n25109, A2 => n24897, B1 => n25103, B2 => 
                           n20025, ZN => n23154);
   U22145 : OAI221_X1 port map( B1 => n21178, B2 => n25067, C1 => n20154, C2 =>
                           n25061, A => n23160, ZN => n23159);
   U22146 : AOI22_X1 port map( A1 => n25055, A2 => n24173, B1 => n25047, B2 => 
                           OUT2_43_port, ZN => n23160);
   U22147 : OAI221_X1 port map( B1 => n21241, B2 => n25121, C1 => n19577, C2 =>
                           n25115, A => n23136, ZN => n23131);
   U22148 : AOI22_X1 port map( A1 => n25109, A2 => n24898, B1 => n25103, B2 => 
                           n20024, ZN => n23136);
   U22149 : OAI221_X1 port map( B1 => n21177, B2 => n25067, C1 => n20153, C2 =>
                           n25061, A => n23142, ZN => n23141);
   U22150 : AOI22_X1 port map( A1 => n25055, A2 => n24175, B1 => n25047, B2 => 
                           OUT2_44_port, ZN => n23142);
   U22151 : OAI221_X1 port map( B1 => n21240, B2 => n25121, C1 => n19576, C2 =>
                           n25115, A => n23118, ZN => n23113);
   U22152 : AOI22_X1 port map( A1 => n25109, A2 => n24899, B1 => n25103, B2 => 
                           n20023, ZN => n23118);
   U22153 : OAI221_X1 port map( B1 => n21176, B2 => n25067, C1 => n20152, C2 =>
                           n25061, A => n23124, ZN => n23123);
   U22154 : AOI22_X1 port map( A1 => n25055, A2 => n24177, B1 => n25047, B2 => 
                           OUT2_45_port, ZN => n23124);
   U22155 : OAI221_X1 port map( B1 => n21239, B2 => n25121, C1 => n19575, C2 =>
                           n25115, A => n23100, ZN => n23095);
   U22156 : AOI22_X1 port map( A1 => n25109, A2 => n24900, B1 => n25103, B2 => 
                           n20022, ZN => n23100);
   U22157 : OAI221_X1 port map( B1 => n21175, B2 => n25067, C1 => n20151, C2 =>
                           n25061, A => n23106, ZN => n23105);
   U22158 : AOI22_X1 port map( A1 => n25055, A2 => n24179, B1 => n25047, B2 => 
                           OUT2_46_port, ZN => n23106);
   U22159 : OAI221_X1 port map( B1 => n21238, B2 => n25121, C1 => n19574, C2 =>
                           n25115, A => n23082, ZN => n23077);
   U22160 : AOI22_X1 port map( A1 => n25109, A2 => n24901, B1 => n25103, B2 => 
                           n20021, ZN => n23082);
   U22161 : OAI221_X1 port map( B1 => n21174, B2 => n25067, C1 => n20150, C2 =>
                           n25061, A => n23088, ZN => n23087);
   U22162 : AOI22_X1 port map( A1 => n25055, A2 => n24181, B1 => n25047, B2 => 
                           OUT2_47_port, ZN => n23088);
   U22163 : OAI221_X1 port map( B1 => n21237, B2 => n25122, C1 => n19573, C2 =>
                           n25116, A => n23064, ZN => n23059);
   U22164 : AOI22_X1 port map( A1 => n25110, A2 => n24902, B1 => n25104, B2 => 
                           n20020, ZN => n23064);
   U22165 : OAI221_X1 port map( B1 => n21173, B2 => n25068, C1 => n20149, C2 =>
                           n25062, A => n23070, ZN => n23069);
   U22166 : AOI22_X1 port map( A1 => n25056, A2 => n24183, B1 => n25047, B2 => 
                           OUT2_48_port, ZN => n23070);
   U22167 : OAI221_X1 port map( B1 => n21236, B2 => n25122, C1 => n19572, C2 =>
                           n25116, A => n23046, ZN => n23041);
   U22168 : AOI22_X1 port map( A1 => n25110, A2 => n24903, B1 => n25104, B2 => 
                           n20019, ZN => n23046);
   U22169 : OAI221_X1 port map( B1 => n21172, B2 => n25068, C1 => n20148, C2 =>
                           n25062, A => n23052, ZN => n23051);
   U22170 : AOI22_X1 port map( A1 => n25056, A2 => n24185, B1 => n25047, B2 => 
                           OUT2_49_port, ZN => n23052);
   U22171 : OAI221_X1 port map( B1 => n21235, B2 => n25122, C1 => n19571, C2 =>
                           n25116, A => n23028, ZN => n23023);
   U22172 : AOI22_X1 port map( A1 => n25110, A2 => n24904, B1 => n25104, B2 => 
                           n20018, ZN => n23028);
   U22173 : OAI221_X1 port map( B1 => n21171, B2 => n25068, C1 => n20147, C2 =>
                           n25062, A => n23034, ZN => n23033);
   U22174 : AOI22_X1 port map( A1 => n25056, A2 => n24187, B1 => n25047, B2 => 
                           OUT2_50_port, ZN => n23034);
   U22175 : OAI221_X1 port map( B1 => n21234, B2 => n25122, C1 => n19570, C2 =>
                           n25116, A => n23010, ZN => n23005);
   U22176 : AOI22_X1 port map( A1 => n25110, A2 => n24905, B1 => n25104, B2 => 
                           n20017, ZN => n23010);
   U22177 : OAI221_X1 port map( B1 => n21170, B2 => n25068, C1 => n20146, C2 =>
                           n25062, A => n23016, ZN => n23015);
   U22178 : AOI22_X1 port map( A1 => n25056, A2 => n24189, B1 => n25047, B2 => 
                           OUT2_51_port, ZN => n23016);
   U22179 : OAI221_X1 port map( B1 => n21233, B2 => n25122, C1 => n19569, C2 =>
                           n25116, A => n22992, ZN => n22987);
   U22180 : AOI22_X1 port map( A1 => n25110, A2 => n24906, B1 => n25104, B2 => 
                           n20016, ZN => n22992);
   U22181 : OAI221_X1 port map( B1 => n21169, B2 => n25068, C1 => n20145, C2 =>
                           n25062, A => n22998, ZN => n22997);
   U22182 : AOI22_X1 port map( A1 => n25056, A2 => n24191, B1 => n25047, B2 => 
                           OUT2_52_port, ZN => n22998);
   U22183 : OAI221_X1 port map( B1 => n21232, B2 => n25122, C1 => n19568, C2 =>
                           n25116, A => n22974, ZN => n22969);
   U22184 : AOI22_X1 port map( A1 => n25110, A2 => n24907, B1 => n25104, B2 => 
                           n20015, ZN => n22974);
   U22185 : OAI221_X1 port map( B1 => n21168, B2 => n25068, C1 => n20144, C2 =>
                           n25062, A => n22980, ZN => n22979);
   U22186 : AOI22_X1 port map( A1 => n25056, A2 => n24193, B1 => n25047, B2 => 
                           OUT2_53_port, ZN => n22980);
   U22187 : OAI221_X1 port map( B1 => n21231, B2 => n25122, C1 => n19567, C2 =>
                           n25116, A => n22956, ZN => n22951);
   U22188 : AOI22_X1 port map( A1 => n25110, A2 => n24908, B1 => n25104, B2 => 
                           n20014, ZN => n22956);
   U22189 : OAI221_X1 port map( B1 => n21167, B2 => n25068, C1 => n20143, C2 =>
                           n25062, A => n22962, ZN => n22961);
   U22190 : AOI22_X1 port map( A1 => n25056, A2 => n24195, B1 => n25047, B2 => 
                           OUT2_54_port, ZN => n22962);
   U22191 : OAI221_X1 port map( B1 => n21230, B2 => n25122, C1 => n19566, C2 =>
                           n25116, A => n22938, ZN => n22933);
   U22192 : AOI22_X1 port map( A1 => n25110, A2 => n24909, B1 => n25104, B2 => 
                           n20013, ZN => n22938);
   U22193 : OAI221_X1 port map( B1 => n21166, B2 => n25068, C1 => n20142, C2 =>
                           n25062, A => n22944, ZN => n22943);
   U22194 : AOI22_X1 port map( A1 => n25056, A2 => n24197, B1 => n25046, B2 => 
                           OUT2_55_port, ZN => n22944);
   U22195 : OAI221_X1 port map( B1 => n21229, B2 => n25122, C1 => n19565, C2 =>
                           n25116, A => n22920, ZN => n22915);
   U22196 : AOI22_X1 port map( A1 => n25110, A2 => n24910, B1 => n25104, B2 => 
                           n20012, ZN => n22920);
   U22197 : OAI221_X1 port map( B1 => n21165, B2 => n25068, C1 => n20141, C2 =>
                           n25062, A => n22926, ZN => n22925);
   U22198 : AOI22_X1 port map( A1 => n25056, A2 => n24199, B1 => n25046, B2 => 
                           OUT2_56_port, ZN => n22926);
   U22199 : OAI221_X1 port map( B1 => n21228, B2 => n25122, C1 => n19564, C2 =>
                           n25116, A => n22902, ZN => n22897);
   U22200 : AOI22_X1 port map( A1 => n25110, A2 => n24911, B1 => n25104, B2 => 
                           n20011, ZN => n22902);
   U22201 : OAI221_X1 port map( B1 => n21164, B2 => n25068, C1 => n20140, C2 =>
                           n25062, A => n22908, ZN => n22907);
   U22202 : AOI22_X1 port map( A1 => n25056, A2 => n24201, B1 => n25046, B2 => 
                           OUT2_57_port, ZN => n22908);
   U22203 : OAI221_X1 port map( B1 => n21227, B2 => n25122, C1 => n19563, C2 =>
                           n25116, A => n22884, ZN => n22879);
   U22204 : AOI22_X1 port map( A1 => n25110, A2 => n24912, B1 => n25104, B2 => 
                           n20010, ZN => n22884);
   U22205 : OAI221_X1 port map( B1 => n21163, B2 => n25068, C1 => n20139, C2 =>
                           n25062, A => n22890, ZN => n22889);
   U22206 : AOI22_X1 port map( A1 => n25056, A2 => n24203, B1 => n25046, B2 => 
                           OUT2_58_port, ZN => n22890);
   U22207 : OAI221_X1 port map( B1 => n21226, B2 => n25122, C1 => n19562, C2 =>
                           n25116, A => n22866, ZN => n22861);
   U22208 : AOI22_X1 port map( A1 => n25110, A2 => n24913, B1 => n25104, B2 => 
                           n20009, ZN => n22866);
   U22209 : OAI221_X1 port map( B1 => n21162, B2 => n25068, C1 => n20138, C2 =>
                           n25062, A => n22872, ZN => n22871);
   U22210 : AOI22_X1 port map( A1 => n25056, A2 => n24205, B1 => n25046, B2 => 
                           OUT2_59_port, ZN => n22872);
   U22211 : OAI221_X1 port map( B1 => n21285, B2 => n25316, C1 => n19621, C2 =>
                           n25310, A => n22739, ZN => n22726);
   U22212 : AOI22_X1 port map( A1 => n25304, A2 => n24854, B1 => n25298, B2 => 
                           n20068, ZN => n22739);
   U22213 : OAI221_X1 port map( B1 => n21221, B2 => n25262, C1 => n20197, C2 =>
                           n25256, A => n22748, ZN => n22747);
   U22214 : AOI22_X1 port map( A1 => n25250, A2 => n24087, B1 => n25244, B2 => 
                           OUT1_0_port, ZN => n22748);
   U22215 : OAI221_X1 port map( B1 => n21284, B2 => n25316, C1 => n19620, C2 =>
                           n25310, A => n22713, ZN => n22708);
   U22216 : AOI22_X1 port map( A1 => n25304, A2 => n24855, B1 => n25298, B2 => 
                           n20067, ZN => n22713);
   U22217 : OAI221_X1 port map( B1 => n21220, B2 => n25262, C1 => n20196, C2 =>
                           n25256, A => n22719, ZN => n22718);
   U22218 : AOI22_X1 port map( A1 => n25250, A2 => n24089, B1 => n25249, B2 => 
                           OUT1_1_port, ZN => n22719);
   U22219 : OAI221_X1 port map( B1 => n21283, B2 => n25316, C1 => n19619, C2 =>
                           n25310, A => n22695, ZN => n22690);
   U22220 : AOI22_X1 port map( A1 => n25304, A2 => n24856, B1 => n25298, B2 => 
                           n20066, ZN => n22695);
   U22221 : OAI221_X1 port map( B1 => n21219, B2 => n25262, C1 => n20195, C2 =>
                           n25256, A => n22701, ZN => n22700);
   U22222 : AOI22_X1 port map( A1 => n25250, A2 => n24091, B1 => n25249, B2 => 
                           OUT1_2_port, ZN => n22701);
   U22223 : OAI221_X1 port map( B1 => n21282, B2 => n25316, C1 => n19618, C2 =>
                           n25310, A => n22677, ZN => n22672);
   U22224 : AOI22_X1 port map( A1 => n25304, A2 => n24857, B1 => n25298, B2 => 
                           n20065, ZN => n22677);
   U22225 : OAI221_X1 port map( B1 => n21218, B2 => n25262, C1 => n20194, C2 =>
                           n25256, A => n22683, ZN => n22682);
   U22226 : AOI22_X1 port map( A1 => n25250, A2 => n24093, B1 => n25249, B2 => 
                           OUT1_3_port, ZN => n22683);
   U22227 : OAI221_X1 port map( B1 => n21281, B2 => n25316, C1 => n19617, C2 =>
                           n25310, A => n22659, ZN => n22654);
   U22228 : AOI22_X1 port map( A1 => n25304, A2 => n24858, B1 => n25298, B2 => 
                           n20064, ZN => n22659);
   U22229 : OAI221_X1 port map( B1 => n21217, B2 => n25262, C1 => n20193, C2 =>
                           n25256, A => n22665, ZN => n22664);
   U22230 : AOI22_X1 port map( A1 => n25250, A2 => n24095, B1 => n25248, B2 => 
                           OUT1_4_port, ZN => n22665);
   U22231 : OAI221_X1 port map( B1 => n21280, B2 => n25316, C1 => n19616, C2 =>
                           n25310, A => n22641, ZN => n22636);
   U22232 : AOI22_X1 port map( A1 => n25304, A2 => n24859, B1 => n25298, B2 => 
                           n20063, ZN => n22641);
   U22233 : OAI221_X1 port map( B1 => n21216, B2 => n25262, C1 => n20192, C2 =>
                           n25256, A => n22647, ZN => n22646);
   U22234 : AOI22_X1 port map( A1 => n25250, A2 => n24097, B1 => n25248, B2 => 
                           OUT1_5_port, ZN => n22647);
   U22235 : OAI221_X1 port map( B1 => n21279, B2 => n25316, C1 => n19615, C2 =>
                           n25310, A => n22623, ZN => n22618);
   U22236 : AOI22_X1 port map( A1 => n25304, A2 => n24860, B1 => n25298, B2 => 
                           n20062, ZN => n22623);
   U22237 : OAI221_X1 port map( B1 => n21215, B2 => n25262, C1 => n20191, C2 =>
                           n25256, A => n22629, ZN => n22628);
   U22238 : AOI22_X1 port map( A1 => n25250, A2 => n24099, B1 => n25248, B2 => 
                           OUT1_6_port, ZN => n22629);
   U22239 : OAI221_X1 port map( B1 => n21278, B2 => n25316, C1 => n19614, C2 =>
                           n25310, A => n22605, ZN => n22600);
   U22240 : AOI22_X1 port map( A1 => n25304, A2 => n24861, B1 => n25298, B2 => 
                           n20061, ZN => n22605);
   U22241 : OAI221_X1 port map( B1 => n21214, B2 => n25262, C1 => n20190, C2 =>
                           n25256, A => n22611, ZN => n22610);
   U22242 : AOI22_X1 port map( A1 => n25250, A2 => n24101, B1 => n25248, B2 => 
                           OUT1_7_port, ZN => n22611);
   U22243 : OAI221_X1 port map( B1 => n21277, B2 => n25316, C1 => n19613, C2 =>
                           n25310, A => n22587, ZN => n22582);
   U22244 : AOI22_X1 port map( A1 => n25304, A2 => n24862, B1 => n25298, B2 => 
                           n20060, ZN => n22587);
   U22245 : OAI221_X1 port map( B1 => n21213, B2 => n25262, C1 => n20189, C2 =>
                           n25256, A => n22593, ZN => n22592);
   U22246 : AOI22_X1 port map( A1 => n25250, A2 => n24103, B1 => n25248, B2 => 
                           OUT1_8_port, ZN => n22593);
   U22247 : OAI221_X1 port map( B1 => n21276, B2 => n25316, C1 => n19612, C2 =>
                           n25310, A => n22569, ZN => n22564);
   U22248 : AOI22_X1 port map( A1 => n25304, A2 => n24863, B1 => n25298, B2 => 
                           n20059, ZN => n22569);
   U22249 : OAI221_X1 port map( B1 => n21212, B2 => n25262, C1 => n20188, C2 =>
                           n25256, A => n22575, ZN => n22574);
   U22250 : AOI22_X1 port map( A1 => n25250, A2 => n24105, B1 => n25248, B2 => 
                           OUT1_9_port, ZN => n22575);
   U22251 : OAI221_X1 port map( B1 => n21275, B2 => n25316, C1 => n19611, C2 =>
                           n25310, A => n22551, ZN => n22546);
   U22252 : AOI22_X1 port map( A1 => n25304, A2 => n24864, B1 => n25298, B2 => 
                           n20058, ZN => n22551);
   U22253 : OAI221_X1 port map( B1 => n21211, B2 => n25262, C1 => n20187, C2 =>
                           n25256, A => n22557, ZN => n22556);
   U22254 : AOI22_X1 port map( A1 => n25250, A2 => n24107, B1 => n25248, B2 => 
                           OUT1_10_port, ZN => n22557);
   U22255 : OAI221_X1 port map( B1 => n21274, B2 => n25316, C1 => n19610, C2 =>
                           n25310, A => n22533, ZN => n22528);
   U22256 : AOI22_X1 port map( A1 => n25304, A2 => n24865, B1 => n25298, B2 => 
                           n20057, ZN => n22533);
   U22257 : OAI221_X1 port map( B1 => n21210, B2 => n25262, C1 => n20186, C2 =>
                           n25256, A => n22539, ZN => n22538);
   U22258 : AOI22_X1 port map( A1 => n25250, A2 => n24109, B1 => n25248, B2 => 
                           OUT1_11_port, ZN => n22539);
   U22259 : OAI221_X1 port map( B1 => n21273, B2 => n25317, C1 => n19609, C2 =>
                           n25311, A => n22515, ZN => n22510);
   U22260 : AOI22_X1 port map( A1 => n25305, A2 => n24866, B1 => n25299, B2 => 
                           n20056, ZN => n22515);
   U22261 : OAI221_X1 port map( B1 => n21209, B2 => n25263, C1 => n20185, C2 =>
                           n25257, A => n22521, ZN => n22520);
   U22262 : AOI22_X1 port map( A1 => n25251, A2 => n24111, B1 => n25248, B2 => 
                           OUT1_12_port, ZN => n22521);
   U22263 : OAI221_X1 port map( B1 => n21272, B2 => n25317, C1 => n19608, C2 =>
                           n25311, A => n22497, ZN => n22492);
   U22264 : AOI22_X1 port map( A1 => n25305, A2 => n24867, B1 => n25299, B2 => 
                           n20055, ZN => n22497);
   U22265 : OAI221_X1 port map( B1 => n21208, B2 => n25263, C1 => n20184, C2 =>
                           n25257, A => n22503, ZN => n22502);
   U22266 : AOI22_X1 port map( A1 => n25251, A2 => n24113, B1 => n25248, B2 => 
                           OUT1_13_port, ZN => n22503);
   U22267 : OAI221_X1 port map( B1 => n21271, B2 => n25317, C1 => n19607, C2 =>
                           n25311, A => n22479, ZN => n22474);
   U22268 : AOI22_X1 port map( A1 => n25305, A2 => n24868, B1 => n25299, B2 => 
                           n20054, ZN => n22479);
   U22269 : OAI221_X1 port map( B1 => n21207, B2 => n25263, C1 => n20183, C2 =>
                           n25257, A => n22485, ZN => n22484);
   U22270 : AOI22_X1 port map( A1 => n25251, A2 => n24115, B1 => n25248, B2 => 
                           OUT1_14_port, ZN => n22485);
   U22271 : OAI221_X1 port map( B1 => n21270, B2 => n25317, C1 => n19606, C2 =>
                           n25311, A => n22461, ZN => n22456);
   U22272 : AOI22_X1 port map( A1 => n25305, A2 => n24869, B1 => n25299, B2 => 
                           n20053, ZN => n22461);
   U22273 : OAI221_X1 port map( B1 => n21206, B2 => n25263, C1 => n20182, C2 =>
                           n25257, A => n22467, ZN => n22466);
   U22274 : AOI22_X1 port map( A1 => n25251, A2 => n24117, B1 => n25248, B2 => 
                           OUT1_15_port, ZN => n22467);
   U22275 : OAI221_X1 port map( B1 => n21269, B2 => n25317, C1 => n19605, C2 =>
                           n25311, A => n22443, ZN => n22438);
   U22276 : AOI22_X1 port map( A1 => n25305, A2 => n24870, B1 => n25299, B2 => 
                           n20052, ZN => n22443);
   U22277 : OAI221_X1 port map( B1 => n21205, B2 => n25263, C1 => n20181, C2 =>
                           n25257, A => n22449, ZN => n22448);
   U22278 : AOI22_X1 port map( A1 => n25251, A2 => n24119, B1 => n25248, B2 => 
                           OUT1_16_port, ZN => n22449);
   U22279 : OAI221_X1 port map( B1 => n21268, B2 => n25317, C1 => n19604, C2 =>
                           n25311, A => n22425, ZN => n22420);
   U22280 : AOI22_X1 port map( A1 => n25305, A2 => n24871, B1 => n25299, B2 => 
                           n20051, ZN => n22425);
   U22281 : OAI221_X1 port map( B1 => n21204, B2 => n25263, C1 => n20180, C2 =>
                           n25257, A => n22431, ZN => n22430);
   U22282 : AOI22_X1 port map( A1 => n25251, A2 => n24121, B1 => n25247, B2 => 
                           OUT1_17_port, ZN => n22431);
   U22283 : OAI221_X1 port map( B1 => n21267, B2 => n25317, C1 => n19603, C2 =>
                           n25311, A => n22407, ZN => n22402);
   U22284 : AOI22_X1 port map( A1 => n25305, A2 => n24872, B1 => n25299, B2 => 
                           n20050, ZN => n22407);
   U22285 : OAI221_X1 port map( B1 => n21203, B2 => n25263, C1 => n20179, C2 =>
                           n25257, A => n22413, ZN => n22412);
   U22286 : AOI22_X1 port map( A1 => n25251, A2 => n24123, B1 => n25247, B2 => 
                           OUT1_18_port, ZN => n22413);
   U22287 : OAI221_X1 port map( B1 => n21266, B2 => n25317, C1 => n19602, C2 =>
                           n25311, A => n22389, ZN => n22384);
   U22288 : AOI22_X1 port map( A1 => n25305, A2 => n24873, B1 => n25299, B2 => 
                           n20049, ZN => n22389);
   U22289 : OAI221_X1 port map( B1 => n21202, B2 => n25263, C1 => n20178, C2 =>
                           n25257, A => n22395, ZN => n22394);
   U22290 : AOI22_X1 port map( A1 => n25251, A2 => n24125, B1 => n25247, B2 => 
                           OUT1_19_port, ZN => n22395);
   U22291 : OAI221_X1 port map( B1 => n21265, B2 => n25317, C1 => n19601, C2 =>
                           n25311, A => n22371, ZN => n22366);
   U22292 : AOI22_X1 port map( A1 => n25305, A2 => n24874, B1 => n25299, B2 => 
                           n20048, ZN => n22371);
   U22293 : OAI221_X1 port map( B1 => n21201, B2 => n25263, C1 => n20177, C2 =>
                           n25257, A => n22377, ZN => n22376);
   U22294 : AOI22_X1 port map( A1 => n25251, A2 => n24127, B1 => n25247, B2 => 
                           OUT1_20_port, ZN => n22377);
   U22295 : OAI221_X1 port map( B1 => n21264, B2 => n25317, C1 => n19600, C2 =>
                           n25311, A => n22353, ZN => n22348);
   U22296 : AOI22_X1 port map( A1 => n25305, A2 => n24875, B1 => n25299, B2 => 
                           n20047, ZN => n22353);
   U22297 : OAI221_X1 port map( B1 => n21200, B2 => n25263, C1 => n20176, C2 =>
                           n25257, A => n22359, ZN => n22358);
   U22298 : AOI22_X1 port map( A1 => n25251, A2 => n24129, B1 => n25247, B2 => 
                           OUT1_21_port, ZN => n22359);
   U22299 : OAI221_X1 port map( B1 => n21263, B2 => n25317, C1 => n19599, C2 =>
                           n25311, A => n22335, ZN => n22330);
   U22300 : AOI22_X1 port map( A1 => n25305, A2 => n24876, B1 => n25299, B2 => 
                           n20046, ZN => n22335);
   U22301 : OAI221_X1 port map( B1 => n21199, B2 => n25263, C1 => n20175, C2 =>
                           n25257, A => n22341, ZN => n22340);
   U22302 : AOI22_X1 port map( A1 => n25251, A2 => n24131, B1 => n25247, B2 => 
                           OUT1_22_port, ZN => n22341);
   U22303 : OAI221_X1 port map( B1 => n21262, B2 => n25317, C1 => n19598, C2 =>
                           n25311, A => n22317, ZN => n22312);
   U22304 : AOI22_X1 port map( A1 => n25305, A2 => n24877, B1 => n25299, B2 => 
                           n20045, ZN => n22317);
   U22305 : OAI221_X1 port map( B1 => n21198, B2 => n25263, C1 => n20174, C2 =>
                           n25257, A => n22323, ZN => n22322);
   U22306 : AOI22_X1 port map( A1 => n25251, A2 => n24133, B1 => n25247, B2 => 
                           OUT1_23_port, ZN => n22323);
   U22307 : OAI221_X1 port map( B1 => n21261, B2 => n25318, C1 => n19597, C2 =>
                           n25312, A => n22299, ZN => n22294);
   U22308 : AOI22_X1 port map( A1 => n25306, A2 => n24878, B1 => n25300, B2 => 
                           n20044, ZN => n22299);
   U22309 : OAI221_X1 port map( B1 => n21197, B2 => n25264, C1 => n20173, C2 =>
                           n25258, A => n22305, ZN => n22304);
   U22310 : AOI22_X1 port map( A1 => n25252, A2 => n24135, B1 => n25247, B2 => 
                           OUT1_24_port, ZN => n22305);
   U22311 : OAI221_X1 port map( B1 => n21260, B2 => n25318, C1 => n19596, C2 =>
                           n25312, A => n22281, ZN => n22276);
   U22312 : AOI22_X1 port map( A1 => n25306, A2 => n24879, B1 => n25300, B2 => 
                           n20043, ZN => n22281);
   U22313 : OAI221_X1 port map( B1 => n21196, B2 => n25264, C1 => n20172, C2 =>
                           n25258, A => n22287, ZN => n22286);
   U22314 : AOI22_X1 port map( A1 => n25252, A2 => n24137, B1 => n25247, B2 => 
                           OUT1_25_port, ZN => n22287);
   U22315 : OAI221_X1 port map( B1 => n21259, B2 => n25318, C1 => n19595, C2 =>
                           n25312, A => n22263, ZN => n22258);
   U22316 : AOI22_X1 port map( A1 => n25306, A2 => n24880, B1 => n25300, B2 => 
                           n20042, ZN => n22263);
   U22317 : OAI221_X1 port map( B1 => n21195, B2 => n25264, C1 => n20171, C2 =>
                           n25258, A => n22269, ZN => n22268);
   U22318 : AOI22_X1 port map( A1 => n25252, A2 => n24139, B1 => n25247, B2 => 
                           OUT1_26_port, ZN => n22269);
   U22319 : OAI221_X1 port map( B1 => n21258, B2 => n25318, C1 => n19594, C2 =>
                           n25312, A => n22245, ZN => n22240);
   U22320 : AOI22_X1 port map( A1 => n25306, A2 => n24881, B1 => n25300, B2 => 
                           n20041, ZN => n22245);
   U22321 : OAI221_X1 port map( B1 => n21194, B2 => n25264, C1 => n20170, C2 =>
                           n25258, A => n22251, ZN => n22250);
   U22322 : AOI22_X1 port map( A1 => n25252, A2 => n24141, B1 => n25247, B2 => 
                           OUT1_27_port, ZN => n22251);
   U22323 : OAI221_X1 port map( B1 => n21257, B2 => n25318, C1 => n19593, C2 =>
                           n25312, A => n22227, ZN => n22222);
   U22324 : AOI22_X1 port map( A1 => n25306, A2 => n24882, B1 => n25300, B2 => 
                           n20040, ZN => n22227);
   U22325 : OAI221_X1 port map( B1 => n21193, B2 => n25264, C1 => n20169, C2 =>
                           n25258, A => n22233, ZN => n22232);
   U22326 : AOI22_X1 port map( A1 => n25252, A2 => n24143, B1 => n25247, B2 => 
                           OUT1_28_port, ZN => n22233);
   U22327 : OAI221_X1 port map( B1 => n21256, B2 => n25318, C1 => n19592, C2 =>
                           n25312, A => n22209, ZN => n22204);
   U22328 : AOI22_X1 port map( A1 => n25306, A2 => n24883, B1 => n25300, B2 => 
                           n20039, ZN => n22209);
   U22329 : OAI221_X1 port map( B1 => n21192, B2 => n25264, C1 => n20168, C2 =>
                           n25258, A => n22215, ZN => n22214);
   U22330 : AOI22_X1 port map( A1 => n25252, A2 => n24145, B1 => n25247, B2 => 
                           OUT1_29_port, ZN => n22215);
   U22331 : OAI221_X1 port map( B1 => n21255, B2 => n25318, C1 => n19591, C2 =>
                           n25312, A => n22191, ZN => n22186);
   U22332 : AOI22_X1 port map( A1 => n25306, A2 => n24884, B1 => n25300, B2 => 
                           n20038, ZN => n22191);
   U22333 : OAI221_X1 port map( B1 => n21191, B2 => n25264, C1 => n20167, C2 =>
                           n25258, A => n22197, ZN => n22196);
   U22334 : AOI22_X1 port map( A1 => n25252, A2 => n24147, B1 => n25246, B2 => 
                           OUT1_30_port, ZN => n22197);
   U22335 : OAI221_X1 port map( B1 => n21254, B2 => n25318, C1 => n19590, C2 =>
                           n25312, A => n22173, ZN => n22168);
   U22336 : AOI22_X1 port map( A1 => n25306, A2 => n24885, B1 => n25300, B2 => 
                           n20037, ZN => n22173);
   U22337 : OAI221_X1 port map( B1 => n21190, B2 => n25264, C1 => n20166, C2 =>
                           n25258, A => n22179, ZN => n22178);
   U22338 : AOI22_X1 port map( A1 => n25252, A2 => n24149, B1 => n25246, B2 => 
                           OUT1_31_port, ZN => n22179);
   U22339 : OAI221_X1 port map( B1 => n21253, B2 => n25318, C1 => n19589, C2 =>
                           n25312, A => n22155, ZN => n22150);
   U22340 : AOI22_X1 port map( A1 => n25306, A2 => n24886, B1 => n25300, B2 => 
                           n20036, ZN => n22155);
   U22341 : OAI221_X1 port map( B1 => n21189, B2 => n25264, C1 => n20165, C2 =>
                           n25258, A => n22161, ZN => n22160);
   U22342 : AOI22_X1 port map( A1 => n25252, A2 => n24151, B1 => n25246, B2 => 
                           OUT1_32_port, ZN => n22161);
   U22343 : OAI221_X1 port map( B1 => n21252, B2 => n25318, C1 => n19588, C2 =>
                           n25312, A => n22137, ZN => n22132);
   U22344 : AOI22_X1 port map( A1 => n25306, A2 => n24887, B1 => n25300, B2 => 
                           n20035, ZN => n22137);
   U22345 : OAI221_X1 port map( B1 => n21188, B2 => n25264, C1 => n20164, C2 =>
                           n25258, A => n22143, ZN => n22142);
   U22346 : AOI22_X1 port map( A1 => n25252, A2 => n24153, B1 => n25246, B2 => 
                           OUT1_33_port, ZN => n22143);
   U22347 : OAI221_X1 port map( B1 => n21251, B2 => n25318, C1 => n19587, C2 =>
                           n25312, A => n22119, ZN => n22114);
   U22348 : AOI22_X1 port map( A1 => n25306, A2 => n24888, B1 => n25300, B2 => 
                           n20034, ZN => n22119);
   U22349 : OAI221_X1 port map( B1 => n21187, B2 => n25264, C1 => n20163, C2 =>
                           n25258, A => n22125, ZN => n22124);
   U22350 : AOI22_X1 port map( A1 => n25252, A2 => n24155, B1 => n25246, B2 => 
                           OUT1_34_port, ZN => n22125);
   U22351 : OAI221_X1 port map( B1 => n21250, B2 => n25318, C1 => n19586, C2 =>
                           n25312, A => n22101, ZN => n22096);
   U22352 : AOI22_X1 port map( A1 => n25306, A2 => n24889, B1 => n25300, B2 => 
                           n20033, ZN => n22101);
   U22353 : OAI221_X1 port map( B1 => n21186, B2 => n25264, C1 => n20162, C2 =>
                           n25258, A => n22107, ZN => n22106);
   U22354 : AOI22_X1 port map( A1 => n25252, A2 => n24157, B1 => n25246, B2 => 
                           OUT1_35_port, ZN => n22107);
   U22355 : OAI221_X1 port map( B1 => n21249, B2 => n25319, C1 => n19585, C2 =>
                           n25313, A => n22083, ZN => n22078);
   U22356 : AOI22_X1 port map( A1 => n25307, A2 => n24890, B1 => n25301, B2 => 
                           n20032, ZN => n22083);
   U22357 : OAI221_X1 port map( B1 => n21185, B2 => n25265, C1 => n20161, C2 =>
                           n25259, A => n22089, ZN => n22088);
   U22358 : AOI22_X1 port map( A1 => n25253, A2 => n24159, B1 => n25246, B2 => 
                           OUT1_36_port, ZN => n22089);
   U22359 : OAI221_X1 port map( B1 => n21248, B2 => n25319, C1 => n19584, C2 =>
                           n25313, A => n22065, ZN => n22060);
   U22360 : AOI22_X1 port map( A1 => n25307, A2 => n24891, B1 => n25301, B2 => 
                           n20031, ZN => n22065);
   U22361 : OAI221_X1 port map( B1 => n21184, B2 => n25265, C1 => n20160, C2 =>
                           n25259, A => n22071, ZN => n22070);
   U22362 : AOI22_X1 port map( A1 => n25253, A2 => n24161, B1 => n25246, B2 => 
                           OUT1_37_port, ZN => n22071);
   U22363 : OAI221_X1 port map( B1 => n21247, B2 => n25319, C1 => n19583, C2 =>
                           n25313, A => n22047, ZN => n22042);
   U22364 : AOI22_X1 port map( A1 => n25307, A2 => n24892, B1 => n25301, B2 => 
                           n20030, ZN => n22047);
   U22365 : OAI221_X1 port map( B1 => n21183, B2 => n25265, C1 => n20159, C2 =>
                           n25259, A => n22053, ZN => n22052);
   U22366 : AOI22_X1 port map( A1 => n25253, A2 => n24163, B1 => n25246, B2 => 
                           OUT1_38_port, ZN => n22053);
   U22367 : OAI221_X1 port map( B1 => n21246, B2 => n25319, C1 => n19582, C2 =>
                           n25313, A => n22029, ZN => n22024);
   U22368 : AOI22_X1 port map( A1 => n25307, A2 => n24893, B1 => n25301, B2 => 
                           n20029, ZN => n22029);
   U22369 : OAI221_X1 port map( B1 => n21182, B2 => n25265, C1 => n20158, C2 =>
                           n25259, A => n22035, ZN => n22034);
   U22370 : AOI22_X1 port map( A1 => n25253, A2 => n24165, B1 => n25246, B2 => 
                           OUT1_39_port, ZN => n22035);
   U22371 : OAI221_X1 port map( B1 => n21245, B2 => n25319, C1 => n19581, C2 =>
                           n25313, A => n22011, ZN => n22006);
   U22372 : AOI22_X1 port map( A1 => n25307, A2 => n24894, B1 => n25301, B2 => 
                           n20028, ZN => n22011);
   U22373 : OAI221_X1 port map( B1 => n21181, B2 => n25265, C1 => n20157, C2 =>
                           n25259, A => n22017, ZN => n22016);
   U22374 : AOI22_X1 port map( A1 => n25253, A2 => n24167, B1 => n25246, B2 => 
                           OUT1_40_port, ZN => n22017);
   U22375 : OAI221_X1 port map( B1 => n21244, B2 => n25319, C1 => n19580, C2 =>
                           n25313, A => n21993, ZN => n21988);
   U22376 : AOI22_X1 port map( A1 => n25307, A2 => n24895, B1 => n25301, B2 => 
                           n20027, ZN => n21993);
   U22377 : OAI221_X1 port map( B1 => n21180, B2 => n25265, C1 => n20156, C2 =>
                           n25259, A => n21999, ZN => n21998);
   U22378 : AOI22_X1 port map( A1 => n25253, A2 => n24169, B1 => n25246, B2 => 
                           OUT1_41_port, ZN => n21999);
   U22379 : OAI221_X1 port map( B1 => n21243, B2 => n25319, C1 => n19579, C2 =>
                           n25313, A => n21975, ZN => n21970);
   U22380 : AOI22_X1 port map( A1 => n25307, A2 => n24896, B1 => n25301, B2 => 
                           n20026, ZN => n21975);
   U22381 : OAI221_X1 port map( B1 => n21179, B2 => n25265, C1 => n20155, C2 =>
                           n25259, A => n21981, ZN => n21980);
   U22382 : AOI22_X1 port map( A1 => n25253, A2 => n24171, B1 => n25245, B2 => 
                           OUT1_42_port, ZN => n21981);
   U22383 : OAI221_X1 port map( B1 => n21242, B2 => n25319, C1 => n19578, C2 =>
                           n25313, A => n21957, ZN => n21952);
   U22384 : AOI22_X1 port map( A1 => n25307, A2 => n24897, B1 => n25301, B2 => 
                           n20025, ZN => n21957);
   U22385 : OAI221_X1 port map( B1 => n21178, B2 => n25265, C1 => n20154, C2 =>
                           n25259, A => n21963, ZN => n21962);
   U22386 : AOI22_X1 port map( A1 => n25253, A2 => n24173, B1 => n25245, B2 => 
                           OUT1_43_port, ZN => n21963);
   U22387 : OAI221_X1 port map( B1 => n21241, B2 => n25319, C1 => n19577, C2 =>
                           n25313, A => n21939, ZN => n21934);
   U22388 : AOI22_X1 port map( A1 => n25307, A2 => n24898, B1 => n25301, B2 => 
                           n20024, ZN => n21939);
   U22389 : OAI221_X1 port map( B1 => n21177, B2 => n25265, C1 => n20153, C2 =>
                           n25259, A => n21945, ZN => n21944);
   U22390 : AOI22_X1 port map( A1 => n25253, A2 => n24175, B1 => n25245, B2 => 
                           OUT1_44_port, ZN => n21945);
   U22391 : OAI221_X1 port map( B1 => n21240, B2 => n25319, C1 => n19576, C2 =>
                           n25313, A => n21921, ZN => n21916);
   U22392 : AOI22_X1 port map( A1 => n25307, A2 => n24899, B1 => n25301, B2 => 
                           n20023, ZN => n21921);
   U22393 : OAI221_X1 port map( B1 => n21176, B2 => n25265, C1 => n20152, C2 =>
                           n25259, A => n21927, ZN => n21926);
   U22394 : AOI22_X1 port map( A1 => n25253, A2 => n24177, B1 => n25245, B2 => 
                           OUT1_45_port, ZN => n21927);
   U22395 : OAI221_X1 port map( B1 => n21239, B2 => n25319, C1 => n19575, C2 =>
                           n25313, A => n21903, ZN => n21898);
   U22396 : AOI22_X1 port map( A1 => n25307, A2 => n24900, B1 => n25301, B2 => 
                           n20022, ZN => n21903);
   U22397 : OAI221_X1 port map( B1 => n21175, B2 => n25265, C1 => n20151, C2 =>
                           n25259, A => n21909, ZN => n21908);
   U22398 : AOI22_X1 port map( A1 => n25253, A2 => n24179, B1 => n25245, B2 => 
                           OUT1_46_port, ZN => n21909);
   U22399 : OAI221_X1 port map( B1 => n21238, B2 => n25319, C1 => n19574, C2 =>
                           n25313, A => n21885, ZN => n21880);
   U22400 : AOI22_X1 port map( A1 => n25307, A2 => n24901, B1 => n25301, B2 => 
                           n20021, ZN => n21885);
   U22401 : OAI221_X1 port map( B1 => n21174, B2 => n25265, C1 => n20150, C2 =>
                           n25259, A => n21891, ZN => n21890);
   U22402 : AOI22_X1 port map( A1 => n25253, A2 => n24181, B1 => n25245, B2 => 
                           OUT1_47_port, ZN => n21891);
   U22403 : OAI221_X1 port map( B1 => n21237, B2 => n25320, C1 => n19573, C2 =>
                           n25314, A => n21867, ZN => n21862);
   U22404 : AOI22_X1 port map( A1 => n25308, A2 => n24902, B1 => n25302, B2 => 
                           n20020, ZN => n21867);
   U22405 : OAI221_X1 port map( B1 => n21173, B2 => n25266, C1 => n20149, C2 =>
                           n25260, A => n21873, ZN => n21872);
   U22406 : AOI22_X1 port map( A1 => n25254, A2 => n24183, B1 => n25245, B2 => 
                           OUT1_48_port, ZN => n21873);
   U22407 : OAI221_X1 port map( B1 => n21236, B2 => n25320, C1 => n19572, C2 =>
                           n25314, A => n21849, ZN => n21844);
   U22408 : AOI22_X1 port map( A1 => n25308, A2 => n24903, B1 => n25302, B2 => 
                           n20019, ZN => n21849);
   U22409 : OAI221_X1 port map( B1 => n21172, B2 => n25266, C1 => n20148, C2 =>
                           n25260, A => n21855, ZN => n21854);
   U22410 : AOI22_X1 port map( A1 => n25254, A2 => n24185, B1 => n25245, B2 => 
                           OUT1_49_port, ZN => n21855);
   U22411 : OAI221_X1 port map( B1 => n21235, B2 => n25320, C1 => n19571, C2 =>
                           n25314, A => n21831, ZN => n21826);
   U22412 : AOI22_X1 port map( A1 => n25308, A2 => n24904, B1 => n25302, B2 => 
                           n20018, ZN => n21831);
   U22413 : OAI221_X1 port map( B1 => n21171, B2 => n25266, C1 => n20147, C2 =>
                           n25260, A => n21837, ZN => n21836);
   U22414 : AOI22_X1 port map( A1 => n25254, A2 => n24187, B1 => n25245, B2 => 
                           OUT1_50_port, ZN => n21837);
   U22415 : OAI221_X1 port map( B1 => n21234, B2 => n25320, C1 => n19570, C2 =>
                           n25314, A => n21813, ZN => n21808);
   U22416 : AOI22_X1 port map( A1 => n25308, A2 => n24905, B1 => n25302, B2 => 
                           n20017, ZN => n21813);
   U22417 : OAI221_X1 port map( B1 => n21170, B2 => n25266, C1 => n20146, C2 =>
                           n25260, A => n21819, ZN => n21818);
   U22418 : AOI22_X1 port map( A1 => n25254, A2 => n24189, B1 => n25245, B2 => 
                           OUT1_51_port, ZN => n21819);
   U22419 : OAI221_X1 port map( B1 => n21233, B2 => n25320, C1 => n19569, C2 =>
                           n25314, A => n21795, ZN => n21790);
   U22420 : AOI22_X1 port map( A1 => n25308, A2 => n24906, B1 => n25302, B2 => 
                           n20016, ZN => n21795);
   U22421 : OAI221_X1 port map( B1 => n21169, B2 => n25266, C1 => n20145, C2 =>
                           n25260, A => n21801, ZN => n21800);
   U22422 : AOI22_X1 port map( A1 => n25254, A2 => n24191, B1 => n25245, B2 => 
                           OUT1_52_port, ZN => n21801);
   U22423 : OAI221_X1 port map( B1 => n21232, B2 => n25320, C1 => n19568, C2 =>
                           n25314, A => n21777, ZN => n21772);
   U22424 : AOI22_X1 port map( A1 => n25308, A2 => n24907, B1 => n25302, B2 => 
                           n20015, ZN => n21777);
   U22425 : OAI221_X1 port map( B1 => n21168, B2 => n25266, C1 => n20144, C2 =>
                           n25260, A => n21783, ZN => n21782);
   U22426 : AOI22_X1 port map( A1 => n25254, A2 => n24193, B1 => n25245, B2 => 
                           OUT1_53_port, ZN => n21783);
   U22427 : OAI221_X1 port map( B1 => n21231, B2 => n25320, C1 => n19567, C2 =>
                           n25314, A => n21759, ZN => n21754);
   U22428 : AOI22_X1 port map( A1 => n25308, A2 => n24908, B1 => n25302, B2 => 
                           n20014, ZN => n21759);
   U22429 : OAI221_X1 port map( B1 => n21167, B2 => n25266, C1 => n20143, C2 =>
                           n25260, A => n21765, ZN => n21764);
   U22430 : AOI22_X1 port map( A1 => n25254, A2 => n24195, B1 => n25245, B2 => 
                           OUT1_54_port, ZN => n21765);
   U22431 : OAI221_X1 port map( B1 => n21230, B2 => n25320, C1 => n19566, C2 =>
                           n25314, A => n21741, ZN => n21736);
   U22432 : AOI22_X1 port map( A1 => n25308, A2 => n24909, B1 => n25302, B2 => 
                           n20013, ZN => n21741);
   U22433 : OAI221_X1 port map( B1 => n21166, B2 => n25266, C1 => n20142, C2 =>
                           n25260, A => n21747, ZN => n21746);
   U22434 : AOI22_X1 port map( A1 => n25254, A2 => n24197, B1 => n25244, B2 => 
                           OUT1_55_port, ZN => n21747);
   U22435 : OAI221_X1 port map( B1 => n21229, B2 => n25320, C1 => n19565, C2 =>
                           n25314, A => n21723, ZN => n21718);
   U22436 : AOI22_X1 port map( A1 => n25308, A2 => n24910, B1 => n25302, B2 => 
                           n20012, ZN => n21723);
   U22437 : OAI221_X1 port map( B1 => n21165, B2 => n25266, C1 => n20141, C2 =>
                           n25260, A => n21729, ZN => n21728);
   U22438 : AOI22_X1 port map( A1 => n25254, A2 => n24199, B1 => n25244, B2 => 
                           OUT1_56_port, ZN => n21729);
   U22439 : OAI221_X1 port map( B1 => n21228, B2 => n25320, C1 => n19564, C2 =>
                           n25314, A => n21705, ZN => n21700);
   U22440 : AOI22_X1 port map( A1 => n25308, A2 => n24911, B1 => n25302, B2 => 
                           n20011, ZN => n21705);
   U22441 : OAI221_X1 port map( B1 => n21164, B2 => n25266, C1 => n20140, C2 =>
                           n25260, A => n21711, ZN => n21710);
   U22442 : AOI22_X1 port map( A1 => n25254, A2 => n24201, B1 => n25244, B2 => 
                           OUT1_57_port, ZN => n21711);
   U22443 : OAI221_X1 port map( B1 => n21227, B2 => n25320, C1 => n19563, C2 =>
                           n25314, A => n21687, ZN => n21682);
   U22444 : AOI22_X1 port map( A1 => n25308, A2 => n24912, B1 => n25302, B2 => 
                           n20010, ZN => n21687);
   U22445 : OAI221_X1 port map( B1 => n21163, B2 => n25266, C1 => n20139, C2 =>
                           n25260, A => n21693, ZN => n21692);
   U22446 : AOI22_X1 port map( A1 => n25254, A2 => n24203, B1 => n25244, B2 => 
                           OUT1_58_port, ZN => n21693);
   U22447 : OAI221_X1 port map( B1 => n21226, B2 => n25320, C1 => n19562, C2 =>
                           n25314, A => n21669, ZN => n21664);
   U22448 : AOI22_X1 port map( A1 => n25308, A2 => n24913, B1 => n25302, B2 => 
                           n20009, ZN => n21669);
   U22449 : OAI221_X1 port map( B1 => n21162, B2 => n25266, C1 => n20138, C2 =>
                           n25260, A => n21675, ZN => n21674);
   U22450 : AOI22_X1 port map( A1 => n25254, A2 => n24205, B1 => n25244, B2 => 
                           OUT1_59_port, ZN => n21675);
   U22451 : OAI22_X1 port map( A1 => n25456, A2 => n20901, B1 => n25783, B2 => 
                           n25448, ZN => n5823);
   U22452 : OAI22_X1 port map( A1 => n25456, A2 => n20900, B1 => n25786, B2 => 
                           n25448, ZN => n5824);
   U22453 : OAI22_X1 port map( A1 => n25456, A2 => n20899, B1 => n25789, B2 => 
                           n25448, ZN => n5825);
   U22454 : OAI22_X1 port map( A1 => n25456, A2 => n20898, B1 => n25792, B2 => 
                           n25448, ZN => n5826);
   U22455 : OAI22_X1 port map( A1 => n25456, A2 => n20897, B1 => n25795, B2 => 
                           n25448, ZN => n5827);
   U22456 : OAI22_X1 port map( A1 => n25456, A2 => n20896, B1 => n25798, B2 => 
                           n25448, ZN => n5828);
   U22457 : OAI22_X1 port map( A1 => n25456, A2 => n20895, B1 => n25801, B2 => 
                           n25448, ZN => n5829);
   U22458 : OAI22_X1 port map( A1 => n25456, A2 => n20894, B1 => n25804, B2 => 
                           n25448, ZN => n5830);
   U22459 : OAI22_X1 port map( A1 => n25456, A2 => n20893, B1 => n25807, B2 => 
                           n25448, ZN => n5831);
   U22460 : OAI22_X1 port map( A1 => n25456, A2 => n20892, B1 => n25810, B2 => 
                           n25448, ZN => n5832);
   U22461 : OAI22_X1 port map( A1 => n25456, A2 => n20891, B1 => n25813, B2 => 
                           n25448, ZN => n5833);
   U22462 : OAI22_X1 port map( A1 => n25456, A2 => n20890, B1 => n25816, B2 => 
                           n25448, ZN => n5834);
   U22463 : OAI22_X1 port map( A1 => n25457, A2 => n20889, B1 => n25819, B2 => 
                           n25449, ZN => n5835);
   U22464 : OAI22_X1 port map( A1 => n25457, A2 => n20888, B1 => n25822, B2 => 
                           n25449, ZN => n5836);
   U22465 : OAI22_X1 port map( A1 => n25457, A2 => n20887, B1 => n25825, B2 => 
                           n25449, ZN => n5837);
   U22466 : OAI22_X1 port map( A1 => n25457, A2 => n20886, B1 => n25828, B2 => 
                           n25449, ZN => n5838);
   U22467 : OAI22_X1 port map( A1 => n25457, A2 => n20885, B1 => n25831, B2 => 
                           n25449, ZN => n5839);
   U22468 : OAI22_X1 port map( A1 => n25457, A2 => n20884, B1 => n25834, B2 => 
                           n25449, ZN => n5840);
   U22469 : OAI22_X1 port map( A1 => n25457, A2 => n20883, B1 => n25837, B2 => 
                           n25449, ZN => n5841);
   U22470 : OAI22_X1 port map( A1 => n25457, A2 => n20882, B1 => n25840, B2 => 
                           n25449, ZN => n5842);
   U22471 : OAI22_X1 port map( A1 => n25457, A2 => n20881, B1 => n25843, B2 => 
                           n25449, ZN => n5843);
   U22472 : OAI22_X1 port map( A1 => n25457, A2 => n20880, B1 => n25846, B2 => 
                           n25449, ZN => n5844);
   U22473 : OAI22_X1 port map( A1 => n25457, A2 => n20879, B1 => n25849, B2 => 
                           n25449, ZN => n5845);
   U22474 : OAI22_X1 port map( A1 => n25457, A2 => n20878, B1 => n25852, B2 => 
                           n25449, ZN => n5846);
   U22475 : OAI22_X1 port map( A1 => n25457, A2 => n20877, B1 => n25855, B2 => 
                           n25450, ZN => n5847);
   U22476 : OAI22_X1 port map( A1 => n25458, A2 => n20876, B1 => n25858, B2 => 
                           n25450, ZN => n5848);
   U22477 : OAI22_X1 port map( A1 => n25458, A2 => n20875, B1 => n25861, B2 => 
                           n25450, ZN => n5849);
   U22478 : OAI22_X1 port map( A1 => n25458, A2 => n20874, B1 => n25864, B2 => 
                           n25450, ZN => n5850);
   U22479 : OAI22_X1 port map( A1 => n25458, A2 => n20873, B1 => n25867, B2 => 
                           n25450, ZN => n5851);
   U22480 : OAI22_X1 port map( A1 => n25458, A2 => n20872, B1 => n25870, B2 => 
                           n25450, ZN => n5852);
   U22481 : OAI22_X1 port map( A1 => n25458, A2 => n20871, B1 => n25873, B2 => 
                           n25450, ZN => n5853);
   U22482 : OAI22_X1 port map( A1 => n25458, A2 => n20870, B1 => n25876, B2 => 
                           n25450, ZN => n5854);
   U22483 : OAI22_X1 port map( A1 => n25458, A2 => n20869, B1 => n25879, B2 => 
                           n25450, ZN => n5855);
   U22484 : OAI22_X1 port map( A1 => n25458, A2 => n20868, B1 => n25882, B2 => 
                           n25450, ZN => n5856);
   U22485 : OAI22_X1 port map( A1 => n25458, A2 => n20867, B1 => n25885, B2 => 
                           n25450, ZN => n5857);
   U22486 : OAI22_X1 port map( A1 => n25458, A2 => n20866, B1 => n25888, B2 => 
                           n25450, ZN => n5858);
   U22487 : OAI22_X1 port map( A1 => n25458, A2 => n20865, B1 => n25891, B2 => 
                           n25451, ZN => n5859);
   U22488 : OAI22_X1 port map( A1 => n25458, A2 => n20864, B1 => n25894, B2 => 
                           n25451, ZN => n5860);
   U22489 : OAI22_X1 port map( A1 => n25459, A2 => n20863, B1 => n25897, B2 => 
                           n25451, ZN => n5861);
   U22490 : OAI22_X1 port map( A1 => n25459, A2 => n20862, B1 => n25900, B2 => 
                           n25451, ZN => n5862);
   U22491 : OAI22_X1 port map( A1 => n25459, A2 => n20861, B1 => n25903, B2 => 
                           n25451, ZN => n5863);
   U22492 : OAI22_X1 port map( A1 => n25459, A2 => n20860, B1 => n25906, B2 => 
                           n25451, ZN => n5864);
   U22493 : OAI22_X1 port map( A1 => n25459, A2 => n20859, B1 => n25909, B2 => 
                           n25451, ZN => n5865);
   U22494 : OAI22_X1 port map( A1 => n25459, A2 => n20858, B1 => n25912, B2 => 
                           n25451, ZN => n5866);
   U22495 : OAI22_X1 port map( A1 => n25459, A2 => n20857, B1 => n25915, B2 => 
                           n25451, ZN => n5867);
   U22496 : OAI22_X1 port map( A1 => n25459, A2 => n20856, B1 => n25918, B2 => 
                           n25451, ZN => n5868);
   U22497 : OAI22_X1 port map( A1 => n25459, A2 => n20855, B1 => n25921, B2 => 
                           n25451, ZN => n5869);
   U22498 : OAI22_X1 port map( A1 => n25459, A2 => n20854, B1 => n25924, B2 => 
                           n25451, ZN => n5870);
   U22499 : OAI22_X1 port map( A1 => n25459, A2 => n20853, B1 => n25927, B2 => 
                           n25452, ZN => n5871);
   U22500 : OAI22_X1 port map( A1 => n25459, A2 => n20852, B1 => n25930, B2 => 
                           n25452, ZN => n5872);
   U22501 : OAI22_X1 port map( A1 => n25459, A2 => n20851, B1 => n25933, B2 => 
                           n25452, ZN => n5873);
   U22502 : OAI22_X1 port map( A1 => n25460, A2 => n20850, B1 => n25936, B2 => 
                           n25452, ZN => n5874);
   U22503 : OAI22_X1 port map( A1 => n25460, A2 => n20849, B1 => n25939, B2 => 
                           n25452, ZN => n5875);
   U22504 : OAI22_X1 port map( A1 => n25460, A2 => n20848, B1 => n25942, B2 => 
                           n25452, ZN => n5876);
   U22505 : OAI22_X1 port map( A1 => n25460, A2 => n20847, B1 => n25945, B2 => 
                           n25452, ZN => n5877);
   U22506 : OAI22_X1 port map( A1 => n25460, A2 => n20846, B1 => n25948, B2 => 
                           n25452, ZN => n5878);
   U22507 : OAI22_X1 port map( A1 => n25460, A2 => n20845, B1 => n25951, B2 => 
                           n25452, ZN => n5879);
   U22508 : OAI22_X1 port map( A1 => n25460, A2 => n20844, B1 => n25954, B2 => 
                           n25452, ZN => n5880);
   U22509 : OAI22_X1 port map( A1 => n25460, A2 => n20843, B1 => n25957, B2 => 
                           n25452, ZN => n5881);
   U22510 : OAI22_X1 port map( A1 => n25460, A2 => n20842, B1 => n25960, B2 => 
                           n25452, ZN => n5882);
   U22511 : OAI22_X1 port map( A1 => n25378, A2 => n20841, B1 => n25783, B2 => 
                           n25370, ZN => n5439);
   U22512 : OAI22_X1 port map( A1 => n25378, A2 => n20840, B1 => n25786, B2 => 
                           n25370, ZN => n5440);
   U22513 : OAI22_X1 port map( A1 => n25378, A2 => n20839, B1 => n25789, B2 => 
                           n25370, ZN => n5441);
   U22514 : OAI22_X1 port map( A1 => n25378, A2 => n20838, B1 => n25792, B2 => 
                           n25370, ZN => n5442);
   U22515 : OAI22_X1 port map( A1 => n25378, A2 => n20837, B1 => n25795, B2 => 
                           n25370, ZN => n5443);
   U22516 : OAI22_X1 port map( A1 => n25378, A2 => n20836, B1 => n25798, B2 => 
                           n25370, ZN => n5444);
   U22517 : OAI22_X1 port map( A1 => n25378, A2 => n20835, B1 => n25801, B2 => 
                           n25370, ZN => n5445);
   U22518 : OAI22_X1 port map( A1 => n25378, A2 => n20834, B1 => n25804, B2 => 
                           n25370, ZN => n5446);
   U22519 : OAI22_X1 port map( A1 => n25378, A2 => n20833, B1 => n25807, B2 => 
                           n25370, ZN => n5447);
   U22520 : OAI22_X1 port map( A1 => n25378, A2 => n20832, B1 => n25810, B2 => 
                           n25370, ZN => n5448);
   U22521 : OAI22_X1 port map( A1 => n25378, A2 => n20831, B1 => n25813, B2 => 
                           n25370, ZN => n5449);
   U22522 : OAI22_X1 port map( A1 => n25378, A2 => n20830, B1 => n25816, B2 => 
                           n25370, ZN => n5450);
   U22523 : OAI22_X1 port map( A1 => n25379, A2 => n20829, B1 => n25819, B2 => 
                           n25371, ZN => n5451);
   U22524 : OAI22_X1 port map( A1 => n25379, A2 => n20828, B1 => n25822, B2 => 
                           n25371, ZN => n5452);
   U22525 : OAI22_X1 port map( A1 => n25379, A2 => n20827, B1 => n25825, B2 => 
                           n25371, ZN => n5453);
   U22526 : OAI22_X1 port map( A1 => n25379, A2 => n20826, B1 => n25828, B2 => 
                           n25371, ZN => n5454);
   U22527 : OAI22_X1 port map( A1 => n25379, A2 => n20825, B1 => n25831, B2 => 
                           n25371, ZN => n5455);
   U22528 : OAI22_X1 port map( A1 => n25379, A2 => n20824, B1 => n25834, B2 => 
                           n25371, ZN => n5456);
   U22529 : OAI22_X1 port map( A1 => n25379, A2 => n20823, B1 => n25837, B2 => 
                           n25371, ZN => n5457);
   U22530 : OAI22_X1 port map( A1 => n25379, A2 => n20822, B1 => n25840, B2 => 
                           n25371, ZN => n5458);
   U22531 : OAI22_X1 port map( A1 => n25379, A2 => n20821, B1 => n25843, B2 => 
                           n25371, ZN => n5459);
   U22532 : OAI22_X1 port map( A1 => n25379, A2 => n20820, B1 => n25846, B2 => 
                           n25371, ZN => n5460);
   U22533 : OAI22_X1 port map( A1 => n25379, A2 => n20819, B1 => n25849, B2 => 
                           n25371, ZN => n5461);
   U22534 : OAI22_X1 port map( A1 => n25379, A2 => n20818, B1 => n25852, B2 => 
                           n25371, ZN => n5462);
   U22535 : OAI22_X1 port map( A1 => n25379, A2 => n20817, B1 => n25855, B2 => 
                           n25372, ZN => n5463);
   U22536 : OAI22_X1 port map( A1 => n25380, A2 => n20816, B1 => n25858, B2 => 
                           n25372, ZN => n5464);
   U22537 : OAI22_X1 port map( A1 => n25380, A2 => n20815, B1 => n25861, B2 => 
                           n25372, ZN => n5465);
   U22538 : OAI22_X1 port map( A1 => n25380, A2 => n20814, B1 => n25864, B2 => 
                           n25372, ZN => n5466);
   U22539 : OAI22_X1 port map( A1 => n25380, A2 => n20813, B1 => n25867, B2 => 
                           n25372, ZN => n5467);
   U22540 : OAI22_X1 port map( A1 => n25380, A2 => n20812, B1 => n25870, B2 => 
                           n25372, ZN => n5468);
   U22541 : OAI22_X1 port map( A1 => n25380, A2 => n20811, B1 => n25873, B2 => 
                           n25372, ZN => n5469);
   U22542 : OAI22_X1 port map( A1 => n25380, A2 => n20810, B1 => n25876, B2 => 
                           n25372, ZN => n5470);
   U22543 : OAI22_X1 port map( A1 => n25380, A2 => n20809, B1 => n25879, B2 => 
                           n25372, ZN => n5471);
   U22544 : OAI22_X1 port map( A1 => n25380, A2 => n20808, B1 => n25882, B2 => 
                           n25372, ZN => n5472);
   U22545 : OAI22_X1 port map( A1 => n25380, A2 => n20807, B1 => n25885, B2 => 
                           n25372, ZN => n5473);
   U22546 : OAI22_X1 port map( A1 => n25380, A2 => n20806, B1 => n25888, B2 => 
                           n25372, ZN => n5474);
   U22547 : OAI22_X1 port map( A1 => n25380, A2 => n20805, B1 => n25891, B2 => 
                           n25373, ZN => n5475);
   U22548 : OAI22_X1 port map( A1 => n25380, A2 => n20804, B1 => n25894, B2 => 
                           n25373, ZN => n5476);
   U22549 : OAI22_X1 port map( A1 => n25381, A2 => n20803, B1 => n25897, B2 => 
                           n25373, ZN => n5477);
   U22550 : OAI22_X1 port map( A1 => n25381, A2 => n20802, B1 => n25900, B2 => 
                           n25373, ZN => n5478);
   U22551 : OAI22_X1 port map( A1 => n25381, A2 => n20801, B1 => n25903, B2 => 
                           n25373, ZN => n5479);
   U22552 : OAI22_X1 port map( A1 => n25381, A2 => n20800, B1 => n25906, B2 => 
                           n25373, ZN => n5480);
   U22553 : OAI22_X1 port map( A1 => n25381, A2 => n20799, B1 => n25909, B2 => 
                           n25373, ZN => n5481);
   U22554 : OAI22_X1 port map( A1 => n25381, A2 => n20798, B1 => n25912, B2 => 
                           n25373, ZN => n5482);
   U22555 : OAI22_X1 port map( A1 => n25381, A2 => n20797, B1 => n25915, B2 => 
                           n25373, ZN => n5483);
   U22556 : OAI22_X1 port map( A1 => n25381, A2 => n20796, B1 => n25918, B2 => 
                           n25373, ZN => n5484);
   U22557 : OAI22_X1 port map( A1 => n25381, A2 => n20795, B1 => n25921, B2 => 
                           n25373, ZN => n5485);
   U22558 : OAI22_X1 port map( A1 => n25381, A2 => n20794, B1 => n25924, B2 => 
                           n25373, ZN => n5486);
   U22559 : OAI22_X1 port map( A1 => n25381, A2 => n20793, B1 => n25927, B2 => 
                           n25374, ZN => n5487);
   U22560 : OAI22_X1 port map( A1 => n25381, A2 => n20792, B1 => n25930, B2 => 
                           n25374, ZN => n5488);
   U22561 : OAI22_X1 port map( A1 => n25381, A2 => n20791, B1 => n25933, B2 => 
                           n25374, ZN => n5489);
   U22562 : OAI22_X1 port map( A1 => n25382, A2 => n20790, B1 => n25936, B2 => 
                           n25374, ZN => n5490);
   U22563 : OAI22_X1 port map( A1 => n25382, A2 => n20789, B1 => n25939, B2 => 
                           n25374, ZN => n5491);
   U22564 : OAI22_X1 port map( A1 => n25382, A2 => n20788, B1 => n25942, B2 => 
                           n25374, ZN => n5492);
   U22565 : OAI22_X1 port map( A1 => n25382, A2 => n20787, B1 => n25945, B2 => 
                           n25374, ZN => n5493);
   U22566 : OAI22_X1 port map( A1 => n25382, A2 => n20786, B1 => n25948, B2 => 
                           n25374, ZN => n5494);
   U22567 : OAI22_X1 port map( A1 => n25382, A2 => n20785, B1 => n25951, B2 => 
                           n25374, ZN => n5495);
   U22568 : OAI22_X1 port map( A1 => n25382, A2 => n20784, B1 => n25954, B2 => 
                           n25374, ZN => n5496);
   U22569 : OAI22_X1 port map( A1 => n25382, A2 => n20783, B1 => n25957, B2 => 
                           n25374, ZN => n5497);
   U22570 : OAI22_X1 port map( A1 => n25382, A2 => n20782, B1 => n25960, B2 => 
                           n25374, ZN => n5498);
   U22571 : OAI22_X1 port map( A1 => n25417, A2 => n20581, B1 => n25783, B2 => 
                           n25409, ZN => n5631);
   U22572 : OAI22_X1 port map( A1 => n25417, A2 => n20580, B1 => n25786, B2 => 
                           n25409, ZN => n5632);
   U22573 : OAI22_X1 port map( A1 => n25417, A2 => n20579, B1 => n25789, B2 => 
                           n25409, ZN => n5633);
   U22574 : OAI22_X1 port map( A1 => n25417, A2 => n20578, B1 => n25792, B2 => 
                           n25409, ZN => n5634);
   U22575 : OAI22_X1 port map( A1 => n25417, A2 => n20577, B1 => n25795, B2 => 
                           n25409, ZN => n5635);
   U22576 : OAI22_X1 port map( A1 => n25417, A2 => n20576, B1 => n25798, B2 => 
                           n25409, ZN => n5636);
   U22577 : OAI22_X1 port map( A1 => n25417, A2 => n20575, B1 => n25801, B2 => 
                           n25409, ZN => n5637);
   U22578 : OAI22_X1 port map( A1 => n25417, A2 => n20574, B1 => n25804, B2 => 
                           n25409, ZN => n5638);
   U22579 : OAI22_X1 port map( A1 => n25417, A2 => n20573, B1 => n25807, B2 => 
                           n25409, ZN => n5639);
   U22580 : OAI22_X1 port map( A1 => n25417, A2 => n20572, B1 => n25810, B2 => 
                           n25409, ZN => n5640);
   U22581 : OAI22_X1 port map( A1 => n25417, A2 => n20571, B1 => n25813, B2 => 
                           n25409, ZN => n5641);
   U22582 : OAI22_X1 port map( A1 => n25417, A2 => n20570, B1 => n25816, B2 => 
                           n25409, ZN => n5642);
   U22583 : OAI22_X1 port map( A1 => n25418, A2 => n20569, B1 => n25819, B2 => 
                           n25410, ZN => n5643);
   U22584 : OAI22_X1 port map( A1 => n25418, A2 => n20568, B1 => n25822, B2 => 
                           n25410, ZN => n5644);
   U22585 : OAI22_X1 port map( A1 => n25418, A2 => n20567, B1 => n25825, B2 => 
                           n25410, ZN => n5645);
   U22586 : OAI22_X1 port map( A1 => n25418, A2 => n20566, B1 => n25828, B2 => 
                           n25410, ZN => n5646);
   U22587 : OAI22_X1 port map( A1 => n25418, A2 => n20565, B1 => n25831, B2 => 
                           n25410, ZN => n5647);
   U22588 : OAI22_X1 port map( A1 => n25418, A2 => n20564, B1 => n25834, B2 => 
                           n25410, ZN => n5648);
   U22589 : OAI22_X1 port map( A1 => n25418, A2 => n20563, B1 => n25837, B2 => 
                           n25410, ZN => n5649);
   U22590 : OAI22_X1 port map( A1 => n25418, A2 => n20562, B1 => n25840, B2 => 
                           n25410, ZN => n5650);
   U22591 : OAI22_X1 port map( A1 => n25418, A2 => n20561, B1 => n25843, B2 => 
                           n25410, ZN => n5651);
   U22592 : OAI22_X1 port map( A1 => n25418, A2 => n20560, B1 => n25846, B2 => 
                           n25410, ZN => n5652);
   U22593 : OAI22_X1 port map( A1 => n25418, A2 => n20559, B1 => n25849, B2 => 
                           n25410, ZN => n5653);
   U22594 : OAI22_X1 port map( A1 => n25418, A2 => n20558, B1 => n25852, B2 => 
                           n25410, ZN => n5654);
   U22595 : OAI22_X1 port map( A1 => n25418, A2 => n20557, B1 => n25855, B2 => 
                           n25411, ZN => n5655);
   U22596 : OAI22_X1 port map( A1 => n25419, A2 => n20556, B1 => n25858, B2 => 
                           n25411, ZN => n5656);
   U22597 : OAI22_X1 port map( A1 => n25419, A2 => n20555, B1 => n25861, B2 => 
                           n25411, ZN => n5657);
   U22598 : OAI22_X1 port map( A1 => n25419, A2 => n20554, B1 => n25864, B2 => 
                           n25411, ZN => n5658);
   U22599 : OAI22_X1 port map( A1 => n25419, A2 => n20553, B1 => n25867, B2 => 
                           n25411, ZN => n5659);
   U22600 : OAI22_X1 port map( A1 => n25419, A2 => n20552, B1 => n25870, B2 => 
                           n25411, ZN => n5660);
   U22601 : OAI22_X1 port map( A1 => n25419, A2 => n20551, B1 => n25873, B2 => 
                           n25411, ZN => n5661);
   U22602 : OAI22_X1 port map( A1 => n25419, A2 => n20550, B1 => n25876, B2 => 
                           n25411, ZN => n5662);
   U22603 : OAI22_X1 port map( A1 => n25419, A2 => n20549, B1 => n25879, B2 => 
                           n25411, ZN => n5663);
   U22604 : OAI22_X1 port map( A1 => n25419, A2 => n20548, B1 => n25882, B2 => 
                           n25411, ZN => n5664);
   U22605 : OAI22_X1 port map( A1 => n25419, A2 => n20547, B1 => n25885, B2 => 
                           n25411, ZN => n5665);
   U22606 : OAI22_X1 port map( A1 => n25419, A2 => n20546, B1 => n25888, B2 => 
                           n25411, ZN => n5666);
   U22607 : OAI22_X1 port map( A1 => n25419, A2 => n20545, B1 => n25891, B2 => 
                           n25412, ZN => n5667);
   U22608 : OAI22_X1 port map( A1 => n25419, A2 => n20544, B1 => n25894, B2 => 
                           n25412, ZN => n5668);
   U22609 : OAI22_X1 port map( A1 => n25420, A2 => n20543, B1 => n25897, B2 => 
                           n25412, ZN => n5669);
   U22610 : OAI22_X1 port map( A1 => n25420, A2 => n20542, B1 => n25900, B2 => 
                           n25412, ZN => n5670);
   U22611 : OAI22_X1 port map( A1 => n25420, A2 => n20541, B1 => n25903, B2 => 
                           n25412, ZN => n5671);
   U22612 : OAI22_X1 port map( A1 => n25420, A2 => n20540, B1 => n25906, B2 => 
                           n25412, ZN => n5672);
   U22613 : OAI22_X1 port map( A1 => n25420, A2 => n20539, B1 => n25909, B2 => 
                           n25412, ZN => n5673);
   U22614 : OAI22_X1 port map( A1 => n25420, A2 => n20538, B1 => n25912, B2 => 
                           n25412, ZN => n5674);
   U22615 : OAI22_X1 port map( A1 => n25420, A2 => n20537, B1 => n25915, B2 => 
                           n25412, ZN => n5675);
   U22616 : OAI22_X1 port map( A1 => n25420, A2 => n20536, B1 => n25918, B2 => 
                           n25412, ZN => n5676);
   U22617 : OAI22_X1 port map( A1 => n25420, A2 => n20535, B1 => n25921, B2 => 
                           n25412, ZN => n5677);
   U22618 : OAI22_X1 port map( A1 => n25420, A2 => n20534, B1 => n25924, B2 => 
                           n25412, ZN => n5678);
   U22619 : OAI22_X1 port map( A1 => n25420, A2 => n20533, B1 => n25927, B2 => 
                           n25413, ZN => n5679);
   U22620 : OAI22_X1 port map( A1 => n25420, A2 => n20532, B1 => n25930, B2 => 
                           n25413, ZN => n5680);
   U22621 : OAI22_X1 port map( A1 => n25420, A2 => n20531, B1 => n25933, B2 => 
                           n25413, ZN => n5681);
   U22622 : OAI22_X1 port map( A1 => n25421, A2 => n20530, B1 => n25936, B2 => 
                           n25413, ZN => n5682);
   U22623 : OAI22_X1 port map( A1 => n25421, A2 => n20529, B1 => n25939, B2 => 
                           n25413, ZN => n5683);
   U22624 : OAI22_X1 port map( A1 => n25421, A2 => n20528, B1 => n25942, B2 => 
                           n25413, ZN => n5684);
   U22625 : OAI22_X1 port map( A1 => n25421, A2 => n20527, B1 => n25945, B2 => 
                           n25413, ZN => n5685);
   U22626 : OAI22_X1 port map( A1 => n25421, A2 => n20526, B1 => n25948, B2 => 
                           n25413, ZN => n5686);
   U22627 : OAI22_X1 port map( A1 => n25421, A2 => n20525, B1 => n25951, B2 => 
                           n25413, ZN => n5687);
   U22628 : OAI22_X1 port map( A1 => n25421, A2 => n20524, B1 => n25954, B2 => 
                           n25413, ZN => n5688);
   U22629 : OAI22_X1 port map( A1 => n25421, A2 => n20523, B1 => n25957, B2 => 
                           n25413, ZN => n5689);
   U22630 : OAI22_X1 port map( A1 => n25421, A2 => n20522, B1 => n25960, B2 => 
                           n25413, ZN => n5690);
   U22631 : OAI22_X1 port map( A1 => n25391, A2 => n20521, B1 => n25783, B2 => 
                           n25383, ZN => n5503);
   U22632 : OAI22_X1 port map( A1 => n25391, A2 => n20520, B1 => n25786, B2 => 
                           n25383, ZN => n5504);
   U22633 : OAI22_X1 port map( A1 => n25391, A2 => n20519, B1 => n25789, B2 => 
                           n25383, ZN => n5505);
   U22634 : OAI22_X1 port map( A1 => n25391, A2 => n20518, B1 => n25792, B2 => 
                           n25383, ZN => n5506);
   U22635 : OAI22_X1 port map( A1 => n25391, A2 => n20517, B1 => n25795, B2 => 
                           n25383, ZN => n5507);
   U22636 : OAI22_X1 port map( A1 => n25391, A2 => n20516, B1 => n25798, B2 => 
                           n25383, ZN => n5508);
   U22637 : OAI22_X1 port map( A1 => n25391, A2 => n20515, B1 => n25801, B2 => 
                           n25383, ZN => n5509);
   U22638 : OAI22_X1 port map( A1 => n25391, A2 => n20514, B1 => n25804, B2 => 
                           n25383, ZN => n5510);
   U22639 : OAI22_X1 port map( A1 => n25391, A2 => n20513, B1 => n25807, B2 => 
                           n25383, ZN => n5511);
   U22640 : OAI22_X1 port map( A1 => n25391, A2 => n20512, B1 => n25810, B2 => 
                           n25383, ZN => n5512);
   U22641 : OAI22_X1 port map( A1 => n25391, A2 => n20511, B1 => n25813, B2 => 
                           n25383, ZN => n5513);
   U22642 : OAI22_X1 port map( A1 => n25391, A2 => n20510, B1 => n25816, B2 => 
                           n25383, ZN => n5514);
   U22643 : OAI22_X1 port map( A1 => n25392, A2 => n20509, B1 => n25819, B2 => 
                           n25384, ZN => n5515);
   U22644 : OAI22_X1 port map( A1 => n25392, A2 => n20508, B1 => n25822, B2 => 
                           n25384, ZN => n5516);
   U22645 : OAI22_X1 port map( A1 => n25392, A2 => n20507, B1 => n25825, B2 => 
                           n25384, ZN => n5517);
   U22646 : OAI22_X1 port map( A1 => n25392, A2 => n20506, B1 => n25828, B2 => 
                           n25384, ZN => n5518);
   U22647 : OAI22_X1 port map( A1 => n25392, A2 => n20505, B1 => n25831, B2 => 
                           n25384, ZN => n5519);
   U22648 : OAI22_X1 port map( A1 => n25392, A2 => n20504, B1 => n25834, B2 => 
                           n25384, ZN => n5520);
   U22649 : OAI22_X1 port map( A1 => n25392, A2 => n20503, B1 => n25837, B2 => 
                           n25384, ZN => n5521);
   U22650 : OAI22_X1 port map( A1 => n25392, A2 => n20502, B1 => n25840, B2 => 
                           n25384, ZN => n5522);
   U22651 : OAI22_X1 port map( A1 => n25392, A2 => n20501, B1 => n25843, B2 => 
                           n25384, ZN => n5523);
   U22652 : OAI22_X1 port map( A1 => n25392, A2 => n20500, B1 => n25846, B2 => 
                           n25384, ZN => n5524);
   U22653 : OAI22_X1 port map( A1 => n25392, A2 => n20499, B1 => n25849, B2 => 
                           n25384, ZN => n5525);
   U22654 : OAI22_X1 port map( A1 => n25392, A2 => n20498, B1 => n25852, B2 => 
                           n25384, ZN => n5526);
   U22655 : OAI22_X1 port map( A1 => n25392, A2 => n20497, B1 => n25855, B2 => 
                           n25385, ZN => n5527);
   U22656 : OAI22_X1 port map( A1 => n25393, A2 => n20496, B1 => n25858, B2 => 
                           n25385, ZN => n5528);
   U22657 : OAI22_X1 port map( A1 => n25393, A2 => n20495, B1 => n25861, B2 => 
                           n25385, ZN => n5529);
   U22658 : OAI22_X1 port map( A1 => n25393, A2 => n20494, B1 => n25864, B2 => 
                           n25385, ZN => n5530);
   U22659 : OAI22_X1 port map( A1 => n25393, A2 => n20493, B1 => n25867, B2 => 
                           n25385, ZN => n5531);
   U22660 : OAI22_X1 port map( A1 => n25393, A2 => n20492, B1 => n25870, B2 => 
                           n25385, ZN => n5532);
   U22661 : OAI22_X1 port map( A1 => n25393, A2 => n20491, B1 => n25873, B2 => 
                           n25385, ZN => n5533);
   U22662 : OAI22_X1 port map( A1 => n25393, A2 => n20490, B1 => n25876, B2 => 
                           n25385, ZN => n5534);
   U22663 : OAI22_X1 port map( A1 => n25393, A2 => n20489, B1 => n25879, B2 => 
                           n25385, ZN => n5535);
   U22664 : OAI22_X1 port map( A1 => n25393, A2 => n20488, B1 => n25882, B2 => 
                           n25385, ZN => n5536);
   U22665 : OAI22_X1 port map( A1 => n25393, A2 => n20487, B1 => n25885, B2 => 
                           n25385, ZN => n5537);
   U22666 : OAI22_X1 port map( A1 => n25393, A2 => n20486, B1 => n25888, B2 => 
                           n25385, ZN => n5538);
   U22667 : OAI22_X1 port map( A1 => n25393, A2 => n20485, B1 => n25891, B2 => 
                           n25386, ZN => n5539);
   U22668 : OAI22_X1 port map( A1 => n25393, A2 => n20484, B1 => n25894, B2 => 
                           n25386, ZN => n5540);
   U22669 : OAI22_X1 port map( A1 => n25394, A2 => n20483, B1 => n25897, B2 => 
                           n25386, ZN => n5541);
   U22670 : OAI22_X1 port map( A1 => n25394, A2 => n20482, B1 => n25900, B2 => 
                           n25386, ZN => n5542);
   U22671 : OAI22_X1 port map( A1 => n25394, A2 => n20481, B1 => n25903, B2 => 
                           n25386, ZN => n5543);
   U22672 : OAI22_X1 port map( A1 => n25394, A2 => n20480, B1 => n25906, B2 => 
                           n25386, ZN => n5544);
   U22673 : OAI22_X1 port map( A1 => n25394, A2 => n20479, B1 => n25909, B2 => 
                           n25386, ZN => n5545);
   U22674 : OAI22_X1 port map( A1 => n25394, A2 => n20478, B1 => n25912, B2 => 
                           n25386, ZN => n5546);
   U22675 : OAI22_X1 port map( A1 => n25394, A2 => n20477, B1 => n25915, B2 => 
                           n25386, ZN => n5547);
   U22676 : OAI22_X1 port map( A1 => n25394, A2 => n20476, B1 => n25918, B2 => 
                           n25386, ZN => n5548);
   U22677 : OAI22_X1 port map( A1 => n25394, A2 => n20475, B1 => n25921, B2 => 
                           n25386, ZN => n5549);
   U22678 : OAI22_X1 port map( A1 => n25394, A2 => n20474, B1 => n25924, B2 => 
                           n25386, ZN => n5550);
   U22679 : OAI22_X1 port map( A1 => n25394, A2 => n20473, B1 => n25927, B2 => 
                           n25387, ZN => n5551);
   U22680 : OAI22_X1 port map( A1 => n25394, A2 => n20472, B1 => n25930, B2 => 
                           n25387, ZN => n5552);
   U22681 : OAI22_X1 port map( A1 => n25394, A2 => n20471, B1 => n25933, B2 => 
                           n25387, ZN => n5553);
   U22682 : OAI22_X1 port map( A1 => n25395, A2 => n20470, B1 => n25936, B2 => 
                           n25387, ZN => n5554);
   U22683 : OAI22_X1 port map( A1 => n25395, A2 => n20469, B1 => n25939, B2 => 
                           n25387, ZN => n5555);
   U22684 : OAI22_X1 port map( A1 => n25395, A2 => n20468, B1 => n25942, B2 => 
                           n25387, ZN => n5556);
   U22685 : OAI22_X1 port map( A1 => n25395, A2 => n20467, B1 => n25945, B2 => 
                           n25387, ZN => n5557);
   U22686 : OAI22_X1 port map( A1 => n25395, A2 => n20466, B1 => n25948, B2 => 
                           n25387, ZN => n5558);
   U22687 : OAI22_X1 port map( A1 => n25395, A2 => n20465, B1 => n25951, B2 => 
                           n25387, ZN => n5559);
   U22688 : OAI22_X1 port map( A1 => n25395, A2 => n20464, B1 => n25954, B2 => 
                           n25387, ZN => n5560);
   U22689 : OAI22_X1 port map( A1 => n25395, A2 => n20463, B1 => n25957, B2 => 
                           n25387, ZN => n5561);
   U22690 : OAI22_X1 port map( A1 => n25395, A2 => n20462, B1 => n25960, B2 => 
                           n25387, ZN => n5562);
   U22691 : OAI22_X1 port map( A1 => n25469, A2 => n21349, B1 => n25782, B2 => 
                           n25461, ZN => n5887);
   U22692 : OAI22_X1 port map( A1 => n25469, A2 => n21348, B1 => n25785, B2 => 
                           n25461, ZN => n5888);
   U22693 : OAI22_X1 port map( A1 => n25469, A2 => n21347, B1 => n25788, B2 => 
                           n25461, ZN => n5889);
   U22694 : OAI22_X1 port map( A1 => n25469, A2 => n21346, B1 => n25791, B2 => 
                           n25461, ZN => n5890);
   U22695 : OAI22_X1 port map( A1 => n25469, A2 => n21345, B1 => n25794, B2 => 
                           n25461, ZN => n5891);
   U22696 : OAI22_X1 port map( A1 => n25469, A2 => n21344, B1 => n25797, B2 => 
                           n25461, ZN => n5892);
   U22697 : OAI22_X1 port map( A1 => n25469, A2 => n21343, B1 => n25800, B2 => 
                           n25461, ZN => n5893);
   U22698 : OAI22_X1 port map( A1 => n25469, A2 => n21342, B1 => n25803, B2 => 
                           n25461, ZN => n5894);
   U22699 : OAI22_X1 port map( A1 => n25469, A2 => n21341, B1 => n25806, B2 => 
                           n25461, ZN => n5895);
   U22700 : OAI22_X1 port map( A1 => n25469, A2 => n21340, B1 => n25809, B2 => 
                           n25461, ZN => n5896);
   U22701 : OAI22_X1 port map( A1 => n25469, A2 => n21339, B1 => n25812, B2 => 
                           n25461, ZN => n5897);
   U22702 : OAI22_X1 port map( A1 => n25469, A2 => n21338, B1 => n25815, B2 => 
                           n25461, ZN => n5898);
   U22703 : OAI22_X1 port map( A1 => n25470, A2 => n21337, B1 => n25818, B2 => 
                           n25462, ZN => n5899);
   U22704 : OAI22_X1 port map( A1 => n25470, A2 => n21336, B1 => n25821, B2 => 
                           n25462, ZN => n5900);
   U22705 : OAI22_X1 port map( A1 => n25470, A2 => n21335, B1 => n25824, B2 => 
                           n25462, ZN => n5901);
   U22706 : OAI22_X1 port map( A1 => n25470, A2 => n21334, B1 => n25827, B2 => 
                           n25462, ZN => n5902);
   U22707 : OAI22_X1 port map( A1 => n25470, A2 => n21333, B1 => n25830, B2 => 
                           n25462, ZN => n5903);
   U22708 : OAI22_X1 port map( A1 => n25470, A2 => n21332, B1 => n25833, B2 => 
                           n25462, ZN => n5904);
   U22709 : OAI22_X1 port map( A1 => n25470, A2 => n21331, B1 => n25836, B2 => 
                           n25462, ZN => n5905);
   U22710 : OAI22_X1 port map( A1 => n25470, A2 => n21330, B1 => n25839, B2 => 
                           n25462, ZN => n5906);
   U22711 : OAI22_X1 port map( A1 => n25470, A2 => n21329, B1 => n25842, B2 => 
                           n25462, ZN => n5907);
   U22712 : OAI22_X1 port map( A1 => n25470, A2 => n21328, B1 => n25845, B2 => 
                           n25462, ZN => n5908);
   U22713 : OAI22_X1 port map( A1 => n25470, A2 => n21327, B1 => n25848, B2 => 
                           n25462, ZN => n5909);
   U22714 : OAI22_X1 port map( A1 => n25470, A2 => n21326, B1 => n25851, B2 => 
                           n25462, ZN => n5910);
   U22715 : OAI22_X1 port map( A1 => n25470, A2 => n21325, B1 => n25854, B2 => 
                           n25463, ZN => n5911);
   U22716 : OAI22_X1 port map( A1 => n25471, A2 => n21324, B1 => n25857, B2 => 
                           n25463, ZN => n5912);
   U22717 : OAI22_X1 port map( A1 => n25471, A2 => n21323, B1 => n25860, B2 => 
                           n25463, ZN => n5913);
   U22718 : OAI22_X1 port map( A1 => n25471, A2 => n21322, B1 => n25863, B2 => 
                           n25463, ZN => n5914);
   U22719 : OAI22_X1 port map( A1 => n25471, A2 => n21321, B1 => n25866, B2 => 
                           n25463, ZN => n5915);
   U22720 : OAI22_X1 port map( A1 => n25471, A2 => n21320, B1 => n25869, B2 => 
                           n25463, ZN => n5916);
   U22721 : OAI22_X1 port map( A1 => n25471, A2 => n21319, B1 => n25872, B2 => 
                           n25463, ZN => n5917);
   U22722 : OAI22_X1 port map( A1 => n25471, A2 => n21318, B1 => n25875, B2 => 
                           n25463, ZN => n5918);
   U22723 : OAI22_X1 port map( A1 => n25471, A2 => n21317, B1 => n25878, B2 => 
                           n25463, ZN => n5919);
   U22724 : OAI22_X1 port map( A1 => n25471, A2 => n21316, B1 => n25881, B2 => 
                           n25463, ZN => n5920);
   U22725 : OAI22_X1 port map( A1 => n25471, A2 => n21315, B1 => n25884, B2 => 
                           n25463, ZN => n5921);
   U22726 : OAI22_X1 port map( A1 => n25471, A2 => n21314, B1 => n25887, B2 => 
                           n25463, ZN => n5922);
   U22727 : OAI22_X1 port map( A1 => n25471, A2 => n21313, B1 => n25890, B2 => 
                           n25464, ZN => n5923);
   U22728 : OAI22_X1 port map( A1 => n25471, A2 => n21312, B1 => n25893, B2 => 
                           n25464, ZN => n5924);
   U22729 : OAI22_X1 port map( A1 => n25472, A2 => n21311, B1 => n25896, B2 => 
                           n25464, ZN => n5925);
   U22730 : OAI22_X1 port map( A1 => n25472, A2 => n21310, B1 => n25899, B2 => 
                           n25464, ZN => n5926);
   U22731 : OAI22_X1 port map( A1 => n25472, A2 => n21309, B1 => n25902, B2 => 
                           n25464, ZN => n5927);
   U22732 : OAI22_X1 port map( A1 => n25472, A2 => n21308, B1 => n25905, B2 => 
                           n25464, ZN => n5928);
   U22733 : OAI22_X1 port map( A1 => n25472, A2 => n21307, B1 => n25908, B2 => 
                           n25464, ZN => n5929);
   U22734 : OAI22_X1 port map( A1 => n25472, A2 => n21306, B1 => n25911, B2 => 
                           n25464, ZN => n5930);
   U22735 : OAI22_X1 port map( A1 => n25472, A2 => n21305, B1 => n25914, B2 => 
                           n25464, ZN => n5931);
   U22736 : OAI22_X1 port map( A1 => n25472, A2 => n21304, B1 => n25917, B2 => 
                           n25464, ZN => n5932);
   U22737 : OAI22_X1 port map( A1 => n25472, A2 => n21303, B1 => n25920, B2 => 
                           n25464, ZN => n5933);
   U22738 : OAI22_X1 port map( A1 => n25472, A2 => n21302, B1 => n25923, B2 => 
                           n25464, ZN => n5934);
   U22739 : OAI22_X1 port map( A1 => n25472, A2 => n21301, B1 => n25926, B2 => 
                           n25465, ZN => n5935);
   U22740 : OAI22_X1 port map( A1 => n25472, A2 => n21300, B1 => n25929, B2 => 
                           n25465, ZN => n5936);
   U22741 : OAI22_X1 port map( A1 => n25472, A2 => n21299, B1 => n25932, B2 => 
                           n25465, ZN => n5937);
   U22742 : OAI22_X1 port map( A1 => n25473, A2 => n21298, B1 => n25935, B2 => 
                           n25465, ZN => n5938);
   U22743 : OAI22_X1 port map( A1 => n25473, A2 => n21297, B1 => n25938, B2 => 
                           n25465, ZN => n5939);
   U22744 : OAI22_X1 port map( A1 => n25473, A2 => n21296, B1 => n25941, B2 => 
                           n25465, ZN => n5940);
   U22745 : OAI22_X1 port map( A1 => n25473, A2 => n21295, B1 => n25944, B2 => 
                           n25465, ZN => n5941);
   U22746 : OAI22_X1 port map( A1 => n25473, A2 => n21294, B1 => n25947, B2 => 
                           n25465, ZN => n5942);
   U22747 : OAI22_X1 port map( A1 => n25473, A2 => n21293, B1 => n25950, B2 => 
                           n25465, ZN => n5943);
   U22748 : OAI22_X1 port map( A1 => n25473, A2 => n21292, B1 => n25953, B2 => 
                           n25465, ZN => n5944);
   U22749 : OAI22_X1 port map( A1 => n25473, A2 => n21291, B1 => n25956, B2 => 
                           n25465, ZN => n5945);
   U22750 : OAI22_X1 port map( A1 => n25473, A2 => n21290, B1 => n25959, B2 => 
                           n25465, ZN => n5946);
   U22751 : OAI22_X1 port map( A1 => n25649, A2 => n20645, B1 => n25781, B2 => 
                           n25641, ZN => n6783);
   U22752 : OAI22_X1 port map( A1 => n25649, A2 => n20644, B1 => n25784, B2 => 
                           n25641, ZN => n6784);
   U22753 : OAI22_X1 port map( A1 => n25649, A2 => n20643, B1 => n25787, B2 => 
                           n25641, ZN => n6785);
   U22754 : OAI22_X1 port map( A1 => n25649, A2 => n20642, B1 => n25790, B2 => 
                           n25641, ZN => n6786);
   U22755 : OAI22_X1 port map( A1 => n25649, A2 => n20641, B1 => n25793, B2 => 
                           n25641, ZN => n6787);
   U22756 : OAI22_X1 port map( A1 => n25649, A2 => n20640, B1 => n25796, B2 => 
                           n25641, ZN => n6788);
   U22757 : OAI22_X1 port map( A1 => n25649, A2 => n20639, B1 => n25799, B2 => 
                           n25641, ZN => n6789);
   U22758 : OAI22_X1 port map( A1 => n25649, A2 => n20638, B1 => n25802, B2 => 
                           n25641, ZN => n6790);
   U22759 : OAI22_X1 port map( A1 => n25649, A2 => n20637, B1 => n25805, B2 => 
                           n25641, ZN => n6791);
   U22760 : OAI22_X1 port map( A1 => n25649, A2 => n20636, B1 => n25808, B2 => 
                           n25641, ZN => n6792);
   U22761 : OAI22_X1 port map( A1 => n25649, A2 => n20635, B1 => n25811, B2 => 
                           n25641, ZN => n6793);
   U22762 : OAI22_X1 port map( A1 => n25649, A2 => n20634, B1 => n25814, B2 => 
                           n25641, ZN => n6794);
   U22763 : OAI22_X1 port map( A1 => n25650, A2 => n20633, B1 => n25817, B2 => 
                           n25642, ZN => n6795);
   U22764 : OAI22_X1 port map( A1 => n25650, A2 => n20632, B1 => n25820, B2 => 
                           n25642, ZN => n6796);
   U22765 : OAI22_X1 port map( A1 => n25650, A2 => n20631, B1 => n25823, B2 => 
                           n25642, ZN => n6797);
   U22766 : OAI22_X1 port map( A1 => n25650, A2 => n20630, B1 => n25826, B2 => 
                           n25642, ZN => n6798);
   U22767 : OAI22_X1 port map( A1 => n25650, A2 => n20629, B1 => n25829, B2 => 
                           n25642, ZN => n6799);
   U22768 : OAI22_X1 port map( A1 => n25650, A2 => n20628, B1 => n25832, B2 => 
                           n25642, ZN => n6800);
   U22769 : OAI22_X1 port map( A1 => n25650, A2 => n20627, B1 => n25835, B2 => 
                           n25642, ZN => n6801);
   U22770 : OAI22_X1 port map( A1 => n25650, A2 => n20626, B1 => n25838, B2 => 
                           n25642, ZN => n6802);
   U22771 : OAI22_X1 port map( A1 => n25650, A2 => n20625, B1 => n25841, B2 => 
                           n25642, ZN => n6803);
   U22772 : OAI22_X1 port map( A1 => n25650, A2 => n20624, B1 => n25844, B2 => 
                           n25642, ZN => n6804);
   U22773 : OAI22_X1 port map( A1 => n25650, A2 => n20623, B1 => n25847, B2 => 
                           n25642, ZN => n6805);
   U22774 : OAI22_X1 port map( A1 => n25650, A2 => n20622, B1 => n25850, B2 => 
                           n25642, ZN => n6806);
   U22775 : OAI22_X1 port map( A1 => n25650, A2 => n20621, B1 => n25853, B2 => 
                           n25643, ZN => n6807);
   U22776 : OAI22_X1 port map( A1 => n25651, A2 => n20620, B1 => n25856, B2 => 
                           n25643, ZN => n6808);
   U22777 : OAI22_X1 port map( A1 => n25651, A2 => n20619, B1 => n25859, B2 => 
                           n25643, ZN => n6809);
   U22778 : OAI22_X1 port map( A1 => n25651, A2 => n20618, B1 => n25862, B2 => 
                           n25643, ZN => n6810);
   U22779 : OAI22_X1 port map( A1 => n25651, A2 => n20617, B1 => n25865, B2 => 
                           n25643, ZN => n6811);
   U22780 : OAI22_X1 port map( A1 => n25651, A2 => n20616, B1 => n25868, B2 => 
                           n25643, ZN => n6812);
   U22781 : OAI22_X1 port map( A1 => n25651, A2 => n20615, B1 => n25871, B2 => 
                           n25643, ZN => n6813);
   U22782 : OAI22_X1 port map( A1 => n25651, A2 => n20614, B1 => n25874, B2 => 
                           n25643, ZN => n6814);
   U22783 : OAI22_X1 port map( A1 => n25651, A2 => n20613, B1 => n25877, B2 => 
                           n25643, ZN => n6815);
   U22784 : OAI22_X1 port map( A1 => n25651, A2 => n20612, B1 => n25880, B2 => 
                           n25643, ZN => n6816);
   U22785 : OAI22_X1 port map( A1 => n25651, A2 => n20611, B1 => n25883, B2 => 
                           n25643, ZN => n6817);
   U22786 : OAI22_X1 port map( A1 => n25651, A2 => n20610, B1 => n25886, B2 => 
                           n25643, ZN => n6818);
   U22787 : OAI22_X1 port map( A1 => n25651, A2 => n20609, B1 => n25889, B2 => 
                           n25644, ZN => n6819);
   U22788 : OAI22_X1 port map( A1 => n25651, A2 => n20608, B1 => n25892, B2 => 
                           n25644, ZN => n6820);
   U22789 : OAI22_X1 port map( A1 => n25652, A2 => n20607, B1 => n25895, B2 => 
                           n25644, ZN => n6821);
   U22790 : OAI22_X1 port map( A1 => n25652, A2 => n20606, B1 => n25898, B2 => 
                           n25644, ZN => n6822);
   U22791 : OAI22_X1 port map( A1 => n25652, A2 => n20605, B1 => n25901, B2 => 
                           n25644, ZN => n6823);
   U22792 : OAI22_X1 port map( A1 => n25652, A2 => n20604, B1 => n25904, B2 => 
                           n25644, ZN => n6824);
   U22793 : OAI22_X1 port map( A1 => n25652, A2 => n20603, B1 => n25907, B2 => 
                           n25644, ZN => n6825);
   U22794 : OAI22_X1 port map( A1 => n25652, A2 => n20602, B1 => n25910, B2 => 
                           n25644, ZN => n6826);
   U22795 : OAI22_X1 port map( A1 => n25652, A2 => n20601, B1 => n25913, B2 => 
                           n25644, ZN => n6827);
   U22796 : OAI22_X1 port map( A1 => n25652, A2 => n20600, B1 => n25916, B2 => 
                           n25644, ZN => n6828);
   U22797 : OAI22_X1 port map( A1 => n25652, A2 => n20599, B1 => n25919, B2 => 
                           n25644, ZN => n6829);
   U22798 : OAI22_X1 port map( A1 => n25652, A2 => n20598, B1 => n25922, B2 => 
                           n25644, ZN => n6830);
   U22799 : OAI22_X1 port map( A1 => n25652, A2 => n20597, B1 => n25925, B2 => 
                           n25645, ZN => n6831);
   U22800 : OAI22_X1 port map( A1 => n25652, A2 => n20596, B1 => n25928, B2 => 
                           n25645, ZN => n6832);
   U22801 : OAI22_X1 port map( A1 => n25652, A2 => n20595, B1 => n25931, B2 => 
                           n25645, ZN => n6833);
   U22802 : OAI22_X1 port map( A1 => n25653, A2 => n20594, B1 => n25934, B2 => 
                           n25645, ZN => n6834);
   U22803 : OAI22_X1 port map( A1 => n25653, A2 => n20593, B1 => n25937, B2 => 
                           n25645, ZN => n6835);
   U22804 : OAI22_X1 port map( A1 => n25653, A2 => n20592, B1 => n25940, B2 => 
                           n25645, ZN => n6836);
   U22805 : OAI22_X1 port map( A1 => n25653, A2 => n20591, B1 => n25943, B2 => 
                           n25645, ZN => n6837);
   U22806 : OAI22_X1 port map( A1 => n25653, A2 => n20590, B1 => n25946, B2 => 
                           n25645, ZN => n6838);
   U22807 : OAI22_X1 port map( A1 => n25653, A2 => n20589, B1 => n25949, B2 => 
                           n25645, ZN => n6839);
   U22808 : OAI22_X1 port map( A1 => n25653, A2 => n20588, B1 => n25952, B2 => 
                           n25645, ZN => n6840);
   U22809 : OAI22_X1 port map( A1 => n25653, A2 => n20587, B1 => n25955, B2 => 
                           n25645, ZN => n6841);
   U22810 : OAI22_X1 port map( A1 => n25653, A2 => n20586, B1 => n25958, B2 => 
                           n25645, ZN => n6842);
   U22811 : OAI22_X1 port map( A1 => n25739, A2 => n20261, B1 => n25781, B2 => 
                           n25731, ZN => n7231);
   U22812 : OAI22_X1 port map( A1 => n25739, A2 => n20260, B1 => n25784, B2 => 
                           n25731, ZN => n7232);
   U22813 : OAI22_X1 port map( A1 => n25739, A2 => n20259, B1 => n25787, B2 => 
                           n25731, ZN => n7233);
   U22814 : OAI22_X1 port map( A1 => n25739, A2 => n20258, B1 => n25790, B2 => 
                           n25731, ZN => n7234);
   U22815 : OAI22_X1 port map( A1 => n25739, A2 => n20257, B1 => n25793, B2 => 
                           n25731, ZN => n7235);
   U22816 : OAI22_X1 port map( A1 => n25739, A2 => n20256, B1 => n25796, B2 => 
                           n25731, ZN => n7236);
   U22817 : OAI22_X1 port map( A1 => n25739, A2 => n20255, B1 => n25799, B2 => 
                           n25731, ZN => n7237);
   U22818 : OAI22_X1 port map( A1 => n25739, A2 => n20254, B1 => n25802, B2 => 
                           n25731, ZN => n7238);
   U22819 : OAI22_X1 port map( A1 => n25739, A2 => n20253, B1 => n25805, B2 => 
                           n25731, ZN => n7239);
   U22820 : OAI22_X1 port map( A1 => n25739, A2 => n20252, B1 => n25808, B2 => 
                           n25731, ZN => n7240);
   U22821 : OAI22_X1 port map( A1 => n25739, A2 => n20251, B1 => n25811, B2 => 
                           n25731, ZN => n7241);
   U22822 : OAI22_X1 port map( A1 => n25739, A2 => n20250, B1 => n25814, B2 => 
                           n25731, ZN => n7242);
   U22823 : OAI22_X1 port map( A1 => n25740, A2 => n20249, B1 => n25817, B2 => 
                           n25732, ZN => n7243);
   U22824 : OAI22_X1 port map( A1 => n25740, A2 => n20248, B1 => n25820, B2 => 
                           n25732, ZN => n7244);
   U22825 : OAI22_X1 port map( A1 => n25740, A2 => n20247, B1 => n25823, B2 => 
                           n25732, ZN => n7245);
   U22826 : OAI22_X1 port map( A1 => n25740, A2 => n20246, B1 => n25826, B2 => 
                           n25732, ZN => n7246);
   U22827 : OAI22_X1 port map( A1 => n25740, A2 => n20245, B1 => n25829, B2 => 
                           n25732, ZN => n7247);
   U22828 : OAI22_X1 port map( A1 => n25740, A2 => n20244, B1 => n25832, B2 => 
                           n25732, ZN => n7248);
   U22829 : OAI22_X1 port map( A1 => n25740, A2 => n20243, B1 => n25835, B2 => 
                           n25732, ZN => n7249);
   U22830 : OAI22_X1 port map( A1 => n25740, A2 => n20242, B1 => n25838, B2 => 
                           n25732, ZN => n7250);
   U22831 : OAI22_X1 port map( A1 => n25740, A2 => n20241, B1 => n25841, B2 => 
                           n25732, ZN => n7251);
   U22832 : OAI22_X1 port map( A1 => n25740, A2 => n20240, B1 => n25844, B2 => 
                           n25732, ZN => n7252);
   U22833 : OAI22_X1 port map( A1 => n25740, A2 => n20239, B1 => n25847, B2 => 
                           n25732, ZN => n7253);
   U22834 : OAI22_X1 port map( A1 => n25740, A2 => n20238, B1 => n25850, B2 => 
                           n25732, ZN => n7254);
   U22835 : OAI22_X1 port map( A1 => n25740, A2 => n20237, B1 => n25853, B2 => 
                           n25733, ZN => n7255);
   U22836 : OAI22_X1 port map( A1 => n25741, A2 => n20236, B1 => n25856, B2 => 
                           n25733, ZN => n7256);
   U22837 : OAI22_X1 port map( A1 => n25741, A2 => n20235, B1 => n25859, B2 => 
                           n25733, ZN => n7257);
   U22838 : OAI22_X1 port map( A1 => n25741, A2 => n20234, B1 => n25862, B2 => 
                           n25733, ZN => n7258);
   U22839 : OAI22_X1 port map( A1 => n25741, A2 => n20233, B1 => n25865, B2 => 
                           n25733, ZN => n7259);
   U22840 : OAI22_X1 port map( A1 => n25741, A2 => n20232, B1 => n25868, B2 => 
                           n25733, ZN => n7260);
   U22841 : OAI22_X1 port map( A1 => n25741, A2 => n20231, B1 => n25871, B2 => 
                           n25733, ZN => n7261);
   U22842 : OAI22_X1 port map( A1 => n25741, A2 => n20230, B1 => n25874, B2 => 
                           n25733, ZN => n7262);
   U22843 : OAI22_X1 port map( A1 => n25741, A2 => n20229, B1 => n25877, B2 => 
                           n25733, ZN => n7263);
   U22844 : OAI22_X1 port map( A1 => n25741, A2 => n20228, B1 => n25880, B2 => 
                           n25733, ZN => n7264);
   U22845 : OAI22_X1 port map( A1 => n25741, A2 => n20227, B1 => n25883, B2 => 
                           n25733, ZN => n7265);
   U22846 : OAI22_X1 port map( A1 => n25741, A2 => n20226, B1 => n25886, B2 => 
                           n25733, ZN => n7266);
   U22847 : OAI22_X1 port map( A1 => n25741, A2 => n20225, B1 => n25889, B2 => 
                           n25734, ZN => n7267);
   U22848 : OAI22_X1 port map( A1 => n25741, A2 => n20224, B1 => n25892, B2 => 
                           n25734, ZN => n7268);
   U22849 : OAI22_X1 port map( A1 => n25742, A2 => n20223, B1 => n25895, B2 => 
                           n25734, ZN => n7269);
   U22850 : OAI22_X1 port map( A1 => n25742, A2 => n20222, B1 => n25898, B2 => 
                           n25734, ZN => n7270);
   U22851 : OAI22_X1 port map( A1 => n25742, A2 => n20221, B1 => n25901, B2 => 
                           n25734, ZN => n7271);
   U22852 : OAI22_X1 port map( A1 => n25742, A2 => n20220, B1 => n25904, B2 => 
                           n25734, ZN => n7272);
   U22853 : OAI22_X1 port map( A1 => n25742, A2 => n20219, B1 => n25907, B2 => 
                           n25734, ZN => n7273);
   U22854 : OAI22_X1 port map( A1 => n25742, A2 => n20218, B1 => n25910, B2 => 
                           n25734, ZN => n7274);
   U22855 : OAI22_X1 port map( A1 => n25742, A2 => n20217, B1 => n25913, B2 => 
                           n25734, ZN => n7275);
   U22856 : OAI22_X1 port map( A1 => n25742, A2 => n20216, B1 => n25916, B2 => 
                           n25734, ZN => n7276);
   U22857 : OAI22_X1 port map( A1 => n25742, A2 => n20215, B1 => n25919, B2 => 
                           n25734, ZN => n7277);
   U22858 : OAI22_X1 port map( A1 => n25742, A2 => n20214, B1 => n25922, B2 => 
                           n25734, ZN => n7278);
   U22859 : OAI22_X1 port map( A1 => n25742, A2 => n20213, B1 => n25925, B2 => 
                           n25735, ZN => n7279);
   U22860 : OAI22_X1 port map( A1 => n25742, A2 => n20212, B1 => n25928, B2 => 
                           n25735, ZN => n7280);
   U22861 : OAI22_X1 port map( A1 => n25742, A2 => n20211, B1 => n25931, B2 => 
                           n25735, ZN => n7281);
   U22862 : OAI22_X1 port map( A1 => n25743, A2 => n20210, B1 => n25934, B2 => 
                           n25735, ZN => n7282);
   U22863 : OAI22_X1 port map( A1 => n25743, A2 => n20209, B1 => n25937, B2 => 
                           n25735, ZN => n7283);
   U22864 : OAI22_X1 port map( A1 => n25743, A2 => n20208, B1 => n25940, B2 => 
                           n25735, ZN => n7284);
   U22865 : OAI22_X1 port map( A1 => n25743, A2 => n20207, B1 => n25943, B2 => 
                           n25735, ZN => n7285);
   U22866 : OAI22_X1 port map( A1 => n25743, A2 => n20206, B1 => n25946, B2 => 
                           n25735, ZN => n7286);
   U22867 : OAI22_X1 port map( A1 => n25743, A2 => n20205, B1 => n25949, B2 => 
                           n25735, ZN => n7287);
   U22868 : OAI22_X1 port map( A1 => n25743, A2 => n20204, B1 => n25952, B2 => 
                           n25735, ZN => n7288);
   U22869 : OAI22_X1 port map( A1 => n25743, A2 => n20203, B1 => n25955, B2 => 
                           n25735, ZN => n7289);
   U22870 : OAI22_X1 port map( A1 => n25743, A2 => n20202, B1 => n25958, B2 => 
                           n25735, ZN => n7290);
   U22871 : OAI22_X1 port map( A1 => n9286, A2 => n25583, B1 => n25782, B2 => 
                           n25577, ZN => n6463);
   U22872 : OAI22_X1 port map( A1 => n9285, A2 => n25583, B1 => n25785, B2 => 
                           n25577, ZN => n6464);
   U22873 : OAI22_X1 port map( A1 => n9284, A2 => n25583, B1 => n25788, B2 => 
                           n25577, ZN => n6465);
   U22874 : OAI22_X1 port map( A1 => n9283, A2 => n25583, B1 => n25791, B2 => 
                           n25577, ZN => n6466);
   U22875 : OAI22_X1 port map( A1 => n9282, A2 => n25583, B1 => n25794, B2 => 
                           n25577, ZN => n6467);
   U22876 : OAI22_X1 port map( A1 => n9281, A2 => n25583, B1 => n25797, B2 => 
                           n25577, ZN => n6468);
   U22877 : OAI22_X1 port map( A1 => n9280, A2 => n25583, B1 => n25800, B2 => 
                           n25577, ZN => n6469);
   U22878 : OAI22_X1 port map( A1 => n9279, A2 => n25583, B1 => n25803, B2 => 
                           n25577, ZN => n6470);
   U22879 : OAI22_X1 port map( A1 => n9278, A2 => n25583, B1 => n25806, B2 => 
                           n25577, ZN => n6471);
   U22880 : OAI22_X1 port map( A1 => n9277, A2 => n25583, B1 => n25809, B2 => 
                           n25577, ZN => n6472);
   U22881 : OAI22_X1 port map( A1 => n9276, A2 => n25583, B1 => n25812, B2 => 
                           n25577, ZN => n6473);
   U22882 : OAI22_X1 port map( A1 => n9275, A2 => n25584, B1 => n25815, B2 => 
                           n25577, ZN => n6474);
   U22883 : OAI22_X1 port map( A1 => n9274, A2 => n25584, B1 => n25818, B2 => 
                           n25578, ZN => n6475);
   U22884 : OAI22_X1 port map( A1 => n9273, A2 => n25584, B1 => n25821, B2 => 
                           n25578, ZN => n6476);
   U22885 : OAI22_X1 port map( A1 => n9272, A2 => n25584, B1 => n25824, B2 => 
                           n25578, ZN => n6477);
   U22886 : OAI22_X1 port map( A1 => n9271, A2 => n25584, B1 => n25827, B2 => 
                           n25578, ZN => n6478);
   U22887 : OAI22_X1 port map( A1 => n9270, A2 => n25584, B1 => n25830, B2 => 
                           n25578, ZN => n6479);
   U22888 : OAI22_X1 port map( A1 => n9269, A2 => n25584, B1 => n25833, B2 => 
                           n25578, ZN => n6480);
   U22889 : OAI22_X1 port map( A1 => n9268, A2 => n25584, B1 => n25836, B2 => 
                           n25578, ZN => n6481);
   U22890 : OAI22_X1 port map( A1 => n9267, A2 => n25584, B1 => n25839, B2 => 
                           n25578, ZN => n6482);
   U22891 : OAI22_X1 port map( A1 => n9266, A2 => n25584, B1 => n25842, B2 => 
                           n25578, ZN => n6483);
   U22892 : OAI22_X1 port map( A1 => n9265, A2 => n25584, B1 => n25845, B2 => 
                           n25578, ZN => n6484);
   U22893 : OAI22_X1 port map( A1 => n9264, A2 => n25584, B1 => n25848, B2 => 
                           n25578, ZN => n6485);
   U22894 : OAI22_X1 port map( A1 => n9263, A2 => n25585, B1 => n25851, B2 => 
                           n25578, ZN => n6486);
   U22895 : OAI22_X1 port map( A1 => n9262, A2 => n25585, B1 => n25854, B2 => 
                           n25579, ZN => n6487);
   U22896 : OAI22_X1 port map( A1 => n9261, A2 => n25585, B1 => n25857, B2 => 
                           n25579, ZN => n6488);
   U22897 : OAI22_X1 port map( A1 => n9260, A2 => n25585, B1 => n25860, B2 => 
                           n25579, ZN => n6489);
   U22898 : OAI22_X1 port map( A1 => n9259, A2 => n25585, B1 => n25863, B2 => 
                           n25579, ZN => n6490);
   U22899 : OAI22_X1 port map( A1 => n9258, A2 => n25585, B1 => n25866, B2 => 
                           n25579, ZN => n6491);
   U22900 : OAI22_X1 port map( A1 => n9257, A2 => n25585, B1 => n25869, B2 => 
                           n25579, ZN => n6492);
   U22901 : OAI22_X1 port map( A1 => n9256, A2 => n25585, B1 => n25872, B2 => 
                           n25579, ZN => n6493);
   U22902 : OAI22_X1 port map( A1 => n9255, A2 => n25585, B1 => n25875, B2 => 
                           n25579, ZN => n6494);
   U22903 : OAI22_X1 port map( A1 => n9254, A2 => n25585, B1 => n25878, B2 => 
                           n25579, ZN => n6495);
   U22904 : OAI22_X1 port map( A1 => n9253, A2 => n25585, B1 => n25881, B2 => 
                           n25579, ZN => n6496);
   U22905 : OAI22_X1 port map( A1 => n9252, A2 => n25585, B1 => n25884, B2 => 
                           n25579, ZN => n6497);
   U22906 : OAI22_X1 port map( A1 => n9251, A2 => n25586, B1 => n25887, B2 => 
                           n25579, ZN => n6498);
   U22907 : OAI22_X1 port map( A1 => n9250, A2 => n25586, B1 => n25890, B2 => 
                           n25580, ZN => n6499);
   U22908 : OAI22_X1 port map( A1 => n9249, A2 => n25586, B1 => n25893, B2 => 
                           n25580, ZN => n6500);
   U22909 : OAI22_X1 port map( A1 => n9248, A2 => n25586, B1 => n25896, B2 => 
                           n25580, ZN => n6501);
   U22910 : OAI22_X1 port map( A1 => n9247, A2 => n25586, B1 => n25899, B2 => 
                           n25580, ZN => n6502);
   U22911 : OAI22_X1 port map( A1 => n9246, A2 => n25586, B1 => n25902, B2 => 
                           n25580, ZN => n6503);
   U22912 : OAI22_X1 port map( A1 => n9245, A2 => n25586, B1 => n25905, B2 => 
                           n25580, ZN => n6504);
   U22913 : OAI22_X1 port map( A1 => n9244, A2 => n25586, B1 => n25908, B2 => 
                           n25580, ZN => n6505);
   U22914 : OAI22_X1 port map( A1 => n9243, A2 => n25586, B1 => n25911, B2 => 
                           n25580, ZN => n6506);
   U22915 : OAI22_X1 port map( A1 => n9242, A2 => n25586, B1 => n25914, B2 => 
                           n25580, ZN => n6507);
   U22916 : OAI22_X1 port map( A1 => n9241, A2 => n25586, B1 => n25917, B2 => 
                           n25580, ZN => n6508);
   U22917 : OAI22_X1 port map( A1 => n9240, A2 => n25586, B1 => n25920, B2 => 
                           n25580, ZN => n6509);
   U22918 : OAI22_X1 port map( A1 => n9239, A2 => n25587, B1 => n25923, B2 => 
                           n25580, ZN => n6510);
   U22919 : OAI22_X1 port map( A1 => n9238, A2 => n25587, B1 => n25926, B2 => 
                           n25581, ZN => n6511);
   U22920 : OAI22_X1 port map( A1 => n9237, A2 => n25587, B1 => n25929, B2 => 
                           n25581, ZN => n6512);
   U22921 : OAI22_X1 port map( A1 => n9236, A2 => n25587, B1 => n25932, B2 => 
                           n25581, ZN => n6513);
   U22922 : OAI22_X1 port map( A1 => n9235, A2 => n25587, B1 => n25935, B2 => 
                           n25581, ZN => n6514);
   U22923 : OAI22_X1 port map( A1 => n9234, A2 => n25587, B1 => n25938, B2 => 
                           n25581, ZN => n6515);
   U22924 : OAI22_X1 port map( A1 => n9233, A2 => n25587, B1 => n25941, B2 => 
                           n25581, ZN => n6516);
   U22925 : OAI22_X1 port map( A1 => n9232, A2 => n25587, B1 => n25944, B2 => 
                           n25581, ZN => n6517);
   U22926 : OAI22_X1 port map( A1 => n9231, A2 => n25587, B1 => n25947, B2 => 
                           n25581, ZN => n6518);
   U22927 : OAI22_X1 port map( A1 => n9230, A2 => n25587, B1 => n25950, B2 => 
                           n25581, ZN => n6519);
   U22928 : OAI22_X1 port map( A1 => n9229, A2 => n25587, B1 => n25953, B2 => 
                           n25581, ZN => n6520);
   U22929 : OAI22_X1 port map( A1 => n9228, A2 => n25587, B1 => n25956, B2 => 
                           n25581, ZN => n6521);
   U22930 : OAI22_X1 port map( A1 => n9227, A2 => n25588, B1 => n25959, B2 => 
                           n25581, ZN => n6522);
   U22931 : OAI22_X1 port map( A1 => n9030, A2 => n25506, B1 => n25782, B2 => 
                           n25500, ZN => n6079);
   U22932 : OAI22_X1 port map( A1 => n9029, A2 => n25506, B1 => n25785, B2 => 
                           n25500, ZN => n6080);
   U22933 : OAI22_X1 port map( A1 => n9028, A2 => n25506, B1 => n25788, B2 => 
                           n25500, ZN => n6081);
   U22934 : OAI22_X1 port map( A1 => n9027, A2 => n25506, B1 => n25791, B2 => 
                           n25500, ZN => n6082);
   U22935 : OAI22_X1 port map( A1 => n9026, A2 => n25506, B1 => n25794, B2 => 
                           n25500, ZN => n6083);
   U22936 : OAI22_X1 port map( A1 => n9025, A2 => n25506, B1 => n25797, B2 => 
                           n25500, ZN => n6084);
   U22937 : OAI22_X1 port map( A1 => n9024, A2 => n25506, B1 => n25800, B2 => 
                           n25500, ZN => n6085);
   U22938 : OAI22_X1 port map( A1 => n9023, A2 => n25506, B1 => n25803, B2 => 
                           n25500, ZN => n6086);
   U22939 : OAI22_X1 port map( A1 => n9022, A2 => n25506, B1 => n25806, B2 => 
                           n25500, ZN => n6087);
   U22940 : OAI22_X1 port map( A1 => n9021, A2 => n25506, B1 => n25809, B2 => 
                           n25500, ZN => n6088);
   U22941 : OAI22_X1 port map( A1 => n9020, A2 => n25506, B1 => n25812, B2 => 
                           n25500, ZN => n6089);
   U22942 : OAI22_X1 port map( A1 => n9019, A2 => n25507, B1 => n25815, B2 => 
                           n25500, ZN => n6090);
   U22943 : OAI22_X1 port map( A1 => n9018, A2 => n25507, B1 => n25818, B2 => 
                           n25501, ZN => n6091);
   U22944 : OAI22_X1 port map( A1 => n9017, A2 => n25507, B1 => n25821, B2 => 
                           n25501, ZN => n6092);
   U22945 : OAI22_X1 port map( A1 => n9016, A2 => n25507, B1 => n25824, B2 => 
                           n25501, ZN => n6093);
   U22946 : OAI22_X1 port map( A1 => n9015, A2 => n25507, B1 => n25827, B2 => 
                           n25501, ZN => n6094);
   U22947 : OAI22_X1 port map( A1 => n9014, A2 => n25507, B1 => n25830, B2 => 
                           n25501, ZN => n6095);
   U22948 : OAI22_X1 port map( A1 => n9013, A2 => n25507, B1 => n25833, B2 => 
                           n25501, ZN => n6096);
   U22949 : OAI22_X1 port map( A1 => n9012, A2 => n25507, B1 => n25836, B2 => 
                           n25501, ZN => n6097);
   U22950 : OAI22_X1 port map( A1 => n9011, A2 => n25507, B1 => n25839, B2 => 
                           n25501, ZN => n6098);
   U22951 : OAI22_X1 port map( A1 => n9010, A2 => n25507, B1 => n25842, B2 => 
                           n25501, ZN => n6099);
   U22952 : OAI22_X1 port map( A1 => n9009, A2 => n25507, B1 => n25845, B2 => 
                           n25501, ZN => n6100);
   U22953 : OAI22_X1 port map( A1 => n9008, A2 => n25507, B1 => n25848, B2 => 
                           n25501, ZN => n6101);
   U22954 : OAI22_X1 port map( A1 => n9007, A2 => n25508, B1 => n25851, B2 => 
                           n25501, ZN => n6102);
   U22955 : OAI22_X1 port map( A1 => n9006, A2 => n25508, B1 => n25854, B2 => 
                           n25502, ZN => n6103);
   U22956 : OAI22_X1 port map( A1 => n9005, A2 => n25508, B1 => n25857, B2 => 
                           n25502, ZN => n6104);
   U22957 : OAI22_X1 port map( A1 => n9004, A2 => n25508, B1 => n25860, B2 => 
                           n25502, ZN => n6105);
   U22958 : OAI22_X1 port map( A1 => n9003, A2 => n25508, B1 => n25863, B2 => 
                           n25502, ZN => n6106);
   U22959 : OAI22_X1 port map( A1 => n9002, A2 => n25508, B1 => n25866, B2 => 
                           n25502, ZN => n6107);
   U22960 : OAI22_X1 port map( A1 => n9001, A2 => n25508, B1 => n25869, B2 => 
                           n25502, ZN => n6108);
   U22961 : OAI22_X1 port map( A1 => n9000, A2 => n25508, B1 => n25872, B2 => 
                           n25502, ZN => n6109);
   U22962 : OAI22_X1 port map( A1 => n8999, A2 => n25508, B1 => n25875, B2 => 
                           n25502, ZN => n6110);
   U22963 : OAI22_X1 port map( A1 => n8998, A2 => n25508, B1 => n25878, B2 => 
                           n25502, ZN => n6111);
   U22964 : OAI22_X1 port map( A1 => n8997, A2 => n25508, B1 => n25881, B2 => 
                           n25502, ZN => n6112);
   U22965 : OAI22_X1 port map( A1 => n8996, A2 => n25508, B1 => n25884, B2 => 
                           n25502, ZN => n6113);
   U22966 : OAI22_X1 port map( A1 => n8995, A2 => n25509, B1 => n25887, B2 => 
                           n25502, ZN => n6114);
   U22967 : OAI22_X1 port map( A1 => n8994, A2 => n25509, B1 => n25890, B2 => 
                           n25503, ZN => n6115);
   U22968 : OAI22_X1 port map( A1 => n8993, A2 => n25509, B1 => n25893, B2 => 
                           n25503, ZN => n6116);
   U22969 : OAI22_X1 port map( A1 => n8992, A2 => n25509, B1 => n25896, B2 => 
                           n25503, ZN => n6117);
   U22970 : OAI22_X1 port map( A1 => n8991, A2 => n25509, B1 => n25899, B2 => 
                           n25503, ZN => n6118);
   U22971 : OAI22_X1 port map( A1 => n8990, A2 => n25509, B1 => n25902, B2 => 
                           n25503, ZN => n6119);
   U22972 : OAI22_X1 port map( A1 => n8989, A2 => n25509, B1 => n25905, B2 => 
                           n25503, ZN => n6120);
   U22973 : OAI22_X1 port map( A1 => n8988, A2 => n25509, B1 => n25908, B2 => 
                           n25503, ZN => n6121);
   U22974 : OAI22_X1 port map( A1 => n8987, A2 => n25509, B1 => n25911, B2 => 
                           n25503, ZN => n6122);
   U22975 : OAI22_X1 port map( A1 => n8986, A2 => n25509, B1 => n25914, B2 => 
                           n25503, ZN => n6123);
   U22976 : OAI22_X1 port map( A1 => n8985, A2 => n25509, B1 => n25917, B2 => 
                           n25503, ZN => n6124);
   U22977 : OAI22_X1 port map( A1 => n8984, A2 => n25509, B1 => n25920, B2 => 
                           n25503, ZN => n6125);
   U22978 : OAI22_X1 port map( A1 => n8983, A2 => n25510, B1 => n25923, B2 => 
                           n25503, ZN => n6126);
   U22979 : OAI22_X1 port map( A1 => n8982, A2 => n25510, B1 => n25926, B2 => 
                           n25504, ZN => n6127);
   U22980 : OAI22_X1 port map( A1 => n8981, A2 => n25510, B1 => n25929, B2 => 
                           n25504, ZN => n6128);
   U22981 : OAI22_X1 port map( A1 => n8980, A2 => n25510, B1 => n25932, B2 => 
                           n25504, ZN => n6129);
   U22982 : OAI22_X1 port map( A1 => n8979, A2 => n25510, B1 => n25935, B2 => 
                           n25504, ZN => n6130);
   U22983 : OAI22_X1 port map( A1 => n8978, A2 => n25510, B1 => n25938, B2 => 
                           n25504, ZN => n6131);
   U22984 : OAI22_X1 port map( A1 => n8977, A2 => n25510, B1 => n25941, B2 => 
                           n25504, ZN => n6132);
   U22985 : OAI22_X1 port map( A1 => n8976, A2 => n25510, B1 => n25944, B2 => 
                           n25504, ZN => n6133);
   U22986 : OAI22_X1 port map( A1 => n8975, A2 => n25510, B1 => n25947, B2 => 
                           n25504, ZN => n6134);
   U22987 : OAI22_X1 port map( A1 => n8974, A2 => n25510, B1 => n25950, B2 => 
                           n25504, ZN => n6135);
   U22988 : OAI22_X1 port map( A1 => n8973, A2 => n25510, B1 => n25953, B2 => 
                           n25504, ZN => n6136);
   U22989 : OAI22_X1 port map( A1 => n8972, A2 => n25510, B1 => n25956, B2 => 
                           n25504, ZN => n6137);
   U22990 : OAI22_X1 port map( A1 => n8971, A2 => n25511, B1 => n25959, B2 => 
                           n25504, ZN => n6138);
   U22991 : OAI22_X1 port map( A1 => n9478, A2 => n25775, B1 => n25769, B2 => 
                           n25781, ZN => n7423);
   U22992 : OAI22_X1 port map( A1 => n9477, A2 => n25775, B1 => n25769, B2 => 
                           n25784, ZN => n7424);
   U22993 : OAI22_X1 port map( A1 => n9476, A2 => n25775, B1 => n25769, B2 => 
                           n25787, ZN => n7425);
   U22994 : OAI22_X1 port map( A1 => n9475, A2 => n25775, B1 => n25769, B2 => 
                           n25790, ZN => n7426);
   U22995 : OAI22_X1 port map( A1 => n9474, A2 => n25775, B1 => n25769, B2 => 
                           n25793, ZN => n7427);
   U22996 : OAI22_X1 port map( A1 => n9473, A2 => n25775, B1 => n25769, B2 => 
                           n25796, ZN => n7428);
   U22997 : OAI22_X1 port map( A1 => n9472, A2 => n25775, B1 => n25769, B2 => 
                           n25799, ZN => n7429);
   U22998 : OAI22_X1 port map( A1 => n9471, A2 => n25775, B1 => n25769, B2 => 
                           n25802, ZN => n7430);
   U22999 : OAI22_X1 port map( A1 => n9470, A2 => n25775, B1 => n25769, B2 => 
                           n25805, ZN => n7431);
   U23000 : OAI22_X1 port map( A1 => n9469, A2 => n25775, B1 => n25769, B2 => 
                           n25808, ZN => n7432);
   U23001 : OAI22_X1 port map( A1 => n9468, A2 => n25775, B1 => n25769, B2 => 
                           n25811, ZN => n7433);
   U23002 : OAI22_X1 port map( A1 => n9467, A2 => n25776, B1 => n25769, B2 => 
                           n25814, ZN => n7434);
   U23003 : OAI22_X1 port map( A1 => n9094, A2 => n25750, B1 => n25781, B2 => 
                           n25744, ZN => n7295);
   U23004 : OAI22_X1 port map( A1 => n9093, A2 => n25750, B1 => n25784, B2 => 
                           n25744, ZN => n7296);
   U23005 : OAI22_X1 port map( A1 => n9092, A2 => n25750, B1 => n25787, B2 => 
                           n25744, ZN => n7297);
   U23006 : OAI22_X1 port map( A1 => n9091, A2 => n25750, B1 => n25790, B2 => 
                           n25744, ZN => n7298);
   U23007 : OAI22_X1 port map( A1 => n9090, A2 => n25750, B1 => n25793, B2 => 
                           n25744, ZN => n7299);
   U23008 : OAI22_X1 port map( A1 => n9089, A2 => n25750, B1 => n25796, B2 => 
                           n25744, ZN => n7300);
   U23009 : OAI22_X1 port map( A1 => n9088, A2 => n25750, B1 => n25799, B2 => 
                           n25744, ZN => n7301);
   U23010 : OAI22_X1 port map( A1 => n9087, A2 => n25750, B1 => n25802, B2 => 
                           n25744, ZN => n7302);
   U23011 : OAI22_X1 port map( A1 => n9086, A2 => n25750, B1 => n25805, B2 => 
                           n25744, ZN => n7303);
   U23012 : OAI22_X1 port map( A1 => n9085, A2 => n25750, B1 => n25808, B2 => 
                           n25744, ZN => n7304);
   U23013 : OAI22_X1 port map( A1 => n9084, A2 => n25750, B1 => n25811, B2 => 
                           n25744, ZN => n7305);
   U23014 : OAI22_X1 port map( A1 => n9083, A2 => n25751, B1 => n25814, B2 => 
                           n25744, ZN => n7306);
   U23015 : OAI22_X1 port map( A1 => n9082, A2 => n25751, B1 => n25817, B2 => 
                           n25745, ZN => n7307);
   U23016 : OAI22_X1 port map( A1 => n9081, A2 => n25751, B1 => n25820, B2 => 
                           n25745, ZN => n7308);
   U23017 : OAI22_X1 port map( A1 => n9080, A2 => n25751, B1 => n25823, B2 => 
                           n25745, ZN => n7309);
   U23018 : OAI22_X1 port map( A1 => n9079, A2 => n25751, B1 => n25826, B2 => 
                           n25745, ZN => n7310);
   U23019 : OAI22_X1 port map( A1 => n9078, A2 => n25751, B1 => n25829, B2 => 
                           n25745, ZN => n7311);
   U23020 : OAI22_X1 port map( A1 => n9077, A2 => n25751, B1 => n25832, B2 => 
                           n25745, ZN => n7312);
   U23021 : OAI22_X1 port map( A1 => n9076, A2 => n25751, B1 => n25835, B2 => 
                           n25745, ZN => n7313);
   U23022 : OAI22_X1 port map( A1 => n9075, A2 => n25751, B1 => n25838, B2 => 
                           n25745, ZN => n7314);
   U23023 : OAI22_X1 port map( A1 => n9074, A2 => n25751, B1 => n25841, B2 => 
                           n25745, ZN => n7315);
   U23024 : OAI22_X1 port map( A1 => n9073, A2 => n25751, B1 => n25844, B2 => 
                           n25745, ZN => n7316);
   U23025 : OAI22_X1 port map( A1 => n9072, A2 => n25751, B1 => n25847, B2 => 
                           n25745, ZN => n7317);
   U23026 : OAI22_X1 port map( A1 => n9071, A2 => n25752, B1 => n25850, B2 => 
                           n25745, ZN => n7318);
   U23027 : OAI22_X1 port map( A1 => n9070, A2 => n25752, B1 => n25853, B2 => 
                           n25746, ZN => n7319);
   U23028 : OAI22_X1 port map( A1 => n9069, A2 => n25752, B1 => n25856, B2 => 
                           n25746, ZN => n7320);
   U23029 : OAI22_X1 port map( A1 => n9068, A2 => n25752, B1 => n25859, B2 => 
                           n25746, ZN => n7321);
   U23030 : OAI22_X1 port map( A1 => n9067, A2 => n25752, B1 => n25862, B2 => 
                           n25746, ZN => n7322);
   U23031 : OAI22_X1 port map( A1 => n9066, A2 => n25752, B1 => n25865, B2 => 
                           n25746, ZN => n7323);
   U23032 : OAI22_X1 port map( A1 => n9065, A2 => n25752, B1 => n25868, B2 => 
                           n25746, ZN => n7324);
   U23033 : OAI22_X1 port map( A1 => n9064, A2 => n25752, B1 => n25871, B2 => 
                           n25746, ZN => n7325);
   U23034 : OAI22_X1 port map( A1 => n9063, A2 => n25752, B1 => n25874, B2 => 
                           n25746, ZN => n7326);
   U23035 : OAI22_X1 port map( A1 => n9062, A2 => n25752, B1 => n25877, B2 => 
                           n25746, ZN => n7327);
   U23036 : OAI22_X1 port map( A1 => n9061, A2 => n25752, B1 => n25880, B2 => 
                           n25746, ZN => n7328);
   U23037 : OAI22_X1 port map( A1 => n9060, A2 => n25752, B1 => n25883, B2 => 
                           n25746, ZN => n7329);
   U23038 : OAI22_X1 port map( A1 => n9059, A2 => n25753, B1 => n25886, B2 => 
                           n25746, ZN => n7330);
   U23039 : OAI22_X1 port map( A1 => n9058, A2 => n25753, B1 => n25889, B2 => 
                           n25747, ZN => n7331);
   U23040 : OAI22_X1 port map( A1 => n9057, A2 => n25753, B1 => n25892, B2 => 
                           n25747, ZN => n7332);
   U23041 : OAI22_X1 port map( A1 => n9056, A2 => n25753, B1 => n25895, B2 => 
                           n25747, ZN => n7333);
   U23042 : OAI22_X1 port map( A1 => n9055, A2 => n25753, B1 => n25898, B2 => 
                           n25747, ZN => n7334);
   U23043 : OAI22_X1 port map( A1 => n9054, A2 => n25753, B1 => n25901, B2 => 
                           n25747, ZN => n7335);
   U23044 : OAI22_X1 port map( A1 => n9053, A2 => n25753, B1 => n25904, B2 => 
                           n25747, ZN => n7336);
   U23045 : OAI22_X1 port map( A1 => n9052, A2 => n25753, B1 => n25907, B2 => 
                           n25747, ZN => n7337);
   U23046 : OAI22_X1 port map( A1 => n9051, A2 => n25753, B1 => n25910, B2 => 
                           n25747, ZN => n7338);
   U23047 : OAI22_X1 port map( A1 => n9050, A2 => n25753, B1 => n25913, B2 => 
                           n25747, ZN => n7339);
   U23048 : OAI22_X1 port map( A1 => n9049, A2 => n25753, B1 => n25916, B2 => 
                           n25747, ZN => n7340);
   U23049 : OAI22_X1 port map( A1 => n9048, A2 => n25753, B1 => n25919, B2 => 
                           n25747, ZN => n7341);
   U23050 : OAI22_X1 port map( A1 => n9047, A2 => n25754, B1 => n25922, B2 => 
                           n25747, ZN => n7342);
   U23051 : OAI22_X1 port map( A1 => n9046, A2 => n25754, B1 => n25925, B2 => 
                           n25748, ZN => n7343);
   U23052 : OAI22_X1 port map( A1 => n9045, A2 => n25754, B1 => n25928, B2 => 
                           n25748, ZN => n7344);
   U23053 : OAI22_X1 port map( A1 => n9044, A2 => n25754, B1 => n25931, B2 => 
                           n25748, ZN => n7345);
   U23054 : OAI22_X1 port map( A1 => n9043, A2 => n25754, B1 => n25934, B2 => 
                           n25748, ZN => n7346);
   U23055 : OAI22_X1 port map( A1 => n9042, A2 => n25754, B1 => n25937, B2 => 
                           n25748, ZN => n7347);
   U23056 : OAI22_X1 port map( A1 => n9041, A2 => n25754, B1 => n25940, B2 => 
                           n25748, ZN => n7348);
   U23057 : OAI22_X1 port map( A1 => n9040, A2 => n25754, B1 => n25943, B2 => 
                           n25748, ZN => n7349);
   U23058 : OAI22_X1 port map( A1 => n9039, A2 => n25754, B1 => n25946, B2 => 
                           n25748, ZN => n7350);
   U23059 : OAI22_X1 port map( A1 => n9038, A2 => n25754, B1 => n25949, B2 => 
                           n25748, ZN => n7351);
   U23060 : OAI22_X1 port map( A1 => n9037, A2 => n25754, B1 => n25952, B2 => 
                           n25748, ZN => n7352);
   U23061 : OAI22_X1 port map( A1 => n9036, A2 => n25754, B1 => n25955, B2 => 
                           n25748, ZN => n7353);
   U23062 : OAI22_X1 port map( A1 => n9035, A2 => n25755, B1 => n25958, B2 => 
                           n25748, ZN => n7354);
   U23063 : OAI22_X1 port map( A1 => n9350, A2 => n25686, B1 => n25781, B2 => 
                           n25680, ZN => n6975);
   U23064 : OAI22_X1 port map( A1 => n9349, A2 => n25686, B1 => n25784, B2 => 
                           n25680, ZN => n6976);
   U23065 : OAI22_X1 port map( A1 => n9348, A2 => n25686, B1 => n25787, B2 => 
                           n25680, ZN => n6977);
   U23066 : OAI22_X1 port map( A1 => n9347, A2 => n25686, B1 => n25790, B2 => 
                           n25680, ZN => n6978);
   U23067 : OAI22_X1 port map( A1 => n9346, A2 => n25686, B1 => n25793, B2 => 
                           n25680, ZN => n6979);
   U23068 : OAI22_X1 port map( A1 => n9345, A2 => n25686, B1 => n25796, B2 => 
                           n25680, ZN => n6980);
   U23069 : OAI22_X1 port map( A1 => n9344, A2 => n25686, B1 => n25799, B2 => 
                           n25680, ZN => n6981);
   U23070 : OAI22_X1 port map( A1 => n9343, A2 => n25686, B1 => n25802, B2 => 
                           n25680, ZN => n6982);
   U23071 : OAI22_X1 port map( A1 => n9342, A2 => n25686, B1 => n25805, B2 => 
                           n25680, ZN => n6983);
   U23072 : OAI22_X1 port map( A1 => n9341, A2 => n25686, B1 => n25808, B2 => 
                           n25680, ZN => n6984);
   U23073 : OAI22_X1 port map( A1 => n9340, A2 => n25686, B1 => n25811, B2 => 
                           n25680, ZN => n6985);
   U23074 : OAI22_X1 port map( A1 => n9339, A2 => n25687, B1 => n25814, B2 => 
                           n25680, ZN => n6986);
   U23075 : OAI22_X1 port map( A1 => n9338, A2 => n25687, B1 => n25817, B2 => 
                           n25681, ZN => n6987);
   U23076 : OAI22_X1 port map( A1 => n9337, A2 => n25687, B1 => n25820, B2 => 
                           n25681, ZN => n6988);
   U23077 : OAI22_X1 port map( A1 => n9336, A2 => n25687, B1 => n25823, B2 => 
                           n25681, ZN => n6989);
   U23078 : OAI22_X1 port map( A1 => n9335, A2 => n25687, B1 => n25826, B2 => 
                           n25681, ZN => n6990);
   U23079 : OAI22_X1 port map( A1 => n9334, A2 => n25687, B1 => n25829, B2 => 
                           n25681, ZN => n6991);
   U23080 : OAI22_X1 port map( A1 => n9333, A2 => n25687, B1 => n25832, B2 => 
                           n25681, ZN => n6992);
   U23081 : OAI22_X1 port map( A1 => n9332, A2 => n25687, B1 => n25835, B2 => 
                           n25681, ZN => n6993);
   U23082 : OAI22_X1 port map( A1 => n9331, A2 => n25687, B1 => n25838, B2 => 
                           n25681, ZN => n6994);
   U23083 : OAI22_X1 port map( A1 => n9330, A2 => n25687, B1 => n25841, B2 => 
                           n25681, ZN => n6995);
   U23084 : OAI22_X1 port map( A1 => n9329, A2 => n25687, B1 => n25844, B2 => 
                           n25681, ZN => n6996);
   U23085 : OAI22_X1 port map( A1 => n9328, A2 => n25687, B1 => n25847, B2 => 
                           n25681, ZN => n6997);
   U23086 : OAI22_X1 port map( A1 => n9327, A2 => n25688, B1 => n25850, B2 => 
                           n25681, ZN => n6998);
   U23087 : OAI22_X1 port map( A1 => n9326, A2 => n25688, B1 => n25853, B2 => 
                           n25682, ZN => n6999);
   U23088 : OAI22_X1 port map( A1 => n9325, A2 => n25688, B1 => n25856, B2 => 
                           n25682, ZN => n7000);
   U23089 : OAI22_X1 port map( A1 => n9324, A2 => n25688, B1 => n25859, B2 => 
                           n25682, ZN => n7001);
   U23090 : OAI22_X1 port map( A1 => n9323, A2 => n25688, B1 => n25862, B2 => 
                           n25682, ZN => n7002);
   U23091 : OAI22_X1 port map( A1 => n9322, A2 => n25688, B1 => n25865, B2 => 
                           n25682, ZN => n7003);
   U23092 : OAI22_X1 port map( A1 => n9321, A2 => n25688, B1 => n25868, B2 => 
                           n25682, ZN => n7004);
   U23093 : OAI22_X1 port map( A1 => n9320, A2 => n25688, B1 => n25871, B2 => 
                           n25682, ZN => n7005);
   U23094 : OAI22_X1 port map( A1 => n9319, A2 => n25688, B1 => n25874, B2 => 
                           n25682, ZN => n7006);
   U23095 : OAI22_X1 port map( A1 => n9318, A2 => n25688, B1 => n25877, B2 => 
                           n25682, ZN => n7007);
   U23096 : OAI22_X1 port map( A1 => n9317, A2 => n25688, B1 => n25880, B2 => 
                           n25682, ZN => n7008);
   U23097 : OAI22_X1 port map( A1 => n9316, A2 => n25688, B1 => n25883, B2 => 
                           n25682, ZN => n7009);
   U23098 : OAI22_X1 port map( A1 => n9315, A2 => n25689, B1 => n25886, B2 => 
                           n25682, ZN => n7010);
   U23099 : OAI22_X1 port map( A1 => n9314, A2 => n25689, B1 => n25889, B2 => 
                           n25683, ZN => n7011);
   U23100 : OAI22_X1 port map( A1 => n9313, A2 => n25689, B1 => n25892, B2 => 
                           n25683, ZN => n7012);
   U23101 : OAI22_X1 port map( A1 => n9312, A2 => n25689, B1 => n25895, B2 => 
                           n25683, ZN => n7013);
   U23102 : OAI22_X1 port map( A1 => n9311, A2 => n25689, B1 => n25898, B2 => 
                           n25683, ZN => n7014);
   U23103 : OAI22_X1 port map( A1 => n9310, A2 => n25689, B1 => n25901, B2 => 
                           n25683, ZN => n7015);
   U23104 : OAI22_X1 port map( A1 => n9309, A2 => n25689, B1 => n25904, B2 => 
                           n25683, ZN => n7016);
   U23105 : OAI22_X1 port map( A1 => n9308, A2 => n25689, B1 => n25907, B2 => 
                           n25683, ZN => n7017);
   U23106 : OAI22_X1 port map( A1 => n9307, A2 => n25689, B1 => n25910, B2 => 
                           n25683, ZN => n7018);
   U23107 : OAI22_X1 port map( A1 => n9306, A2 => n25689, B1 => n25913, B2 => 
                           n25683, ZN => n7019);
   U23108 : OAI22_X1 port map( A1 => n9305, A2 => n25689, B1 => n25916, B2 => 
                           n25683, ZN => n7020);
   U23109 : OAI22_X1 port map( A1 => n9304, A2 => n25689, B1 => n25919, B2 => 
                           n25683, ZN => n7021);
   U23110 : OAI22_X1 port map( A1 => n9303, A2 => n25690, B1 => n25922, B2 => 
                           n25683, ZN => n7022);
   U23111 : OAI22_X1 port map( A1 => n9302, A2 => n25690, B1 => n25925, B2 => 
                           n25684, ZN => n7023);
   U23112 : OAI22_X1 port map( A1 => n9301, A2 => n25690, B1 => n25928, B2 => 
                           n25684, ZN => n7024);
   U23113 : OAI22_X1 port map( A1 => n9300, A2 => n25690, B1 => n25931, B2 => 
                           n25684, ZN => n7025);
   U23114 : OAI22_X1 port map( A1 => n9299, A2 => n25690, B1 => n25934, B2 => 
                           n25684, ZN => n7026);
   U23115 : OAI22_X1 port map( A1 => n9298, A2 => n25690, B1 => n25937, B2 => 
                           n25684, ZN => n7027);
   U23116 : OAI22_X1 port map( A1 => n9297, A2 => n25690, B1 => n25940, B2 => 
                           n25684, ZN => n7028);
   U23117 : OAI22_X1 port map( A1 => n9296, A2 => n25690, B1 => n25943, B2 => 
                           n25684, ZN => n7029);
   U23118 : OAI22_X1 port map( A1 => n9295, A2 => n25690, B1 => n25946, B2 => 
                           n25684, ZN => n7030);
   U23119 : OAI22_X1 port map( A1 => n9294, A2 => n25690, B1 => n25949, B2 => 
                           n25684, ZN => n7031);
   U23120 : OAI22_X1 port map( A1 => n9293, A2 => n25690, B1 => n25952, B2 => 
                           n25684, ZN => n7032);
   U23121 : OAI22_X1 port map( A1 => n9292, A2 => n25690, B1 => n25955, B2 => 
                           n25684, ZN => n7033);
   U23122 : OAI22_X1 port map( A1 => n9291, A2 => n25691, B1 => n25958, B2 => 
                           n25684, ZN => n7034);
   U23123 : OAI22_X1 port map( A1 => n25495, A2 => n19940, B1 => n25782, B2 => 
                           n25487, ZN => n6015);
   U23124 : OAI22_X1 port map( A1 => n25495, A2 => n19939, B1 => n25785, B2 => 
                           n25487, ZN => n6016);
   U23125 : OAI22_X1 port map( A1 => n25495, A2 => n19938, B1 => n25788, B2 => 
                           n25487, ZN => n6017);
   U23126 : OAI22_X1 port map( A1 => n25495, A2 => n19937, B1 => n25791, B2 => 
                           n25487, ZN => n6018);
   U23127 : OAI22_X1 port map( A1 => n25495, A2 => n19936, B1 => n25794, B2 => 
                           n25487, ZN => n6019);
   U23128 : OAI22_X1 port map( A1 => n25495, A2 => n19935, B1 => n25797, B2 => 
                           n25487, ZN => n6020);
   U23129 : OAI22_X1 port map( A1 => n25495, A2 => n19934, B1 => n25800, B2 => 
                           n25487, ZN => n6021);
   U23130 : OAI22_X1 port map( A1 => n25495, A2 => n19933, B1 => n25803, B2 => 
                           n25487, ZN => n6022);
   U23131 : OAI22_X1 port map( A1 => n25495, A2 => n19932, B1 => n25806, B2 => 
                           n25487, ZN => n6023);
   U23132 : OAI22_X1 port map( A1 => n25495, A2 => n19931, B1 => n25809, B2 => 
                           n25487, ZN => n6024);
   U23133 : OAI22_X1 port map( A1 => n25495, A2 => n19930, B1 => n25812, B2 => 
                           n25487, ZN => n6025);
   U23134 : OAI22_X1 port map( A1 => n25495, A2 => n19929, B1 => n25815, B2 => 
                           n25487, ZN => n6026);
   U23135 : OAI22_X1 port map( A1 => n25496, A2 => n19928, B1 => n25818, B2 => 
                           n25488, ZN => n6027);
   U23136 : OAI22_X1 port map( A1 => n25496, A2 => n19927, B1 => n25821, B2 => 
                           n25488, ZN => n6028);
   U23137 : OAI22_X1 port map( A1 => n25496, A2 => n19926, B1 => n25824, B2 => 
                           n25488, ZN => n6029);
   U23138 : OAI22_X1 port map( A1 => n25496, A2 => n19925, B1 => n25827, B2 => 
                           n25488, ZN => n6030);
   U23139 : OAI22_X1 port map( A1 => n25496, A2 => n19924, B1 => n25830, B2 => 
                           n25488, ZN => n6031);
   U23140 : OAI22_X1 port map( A1 => n25496, A2 => n19923, B1 => n25833, B2 => 
                           n25488, ZN => n6032);
   U23141 : OAI22_X1 port map( A1 => n25496, A2 => n19922, B1 => n25836, B2 => 
                           n25488, ZN => n6033);
   U23142 : OAI22_X1 port map( A1 => n25496, A2 => n19921, B1 => n25839, B2 => 
                           n25488, ZN => n6034);
   U23143 : OAI22_X1 port map( A1 => n25496, A2 => n19920, B1 => n25842, B2 => 
                           n25488, ZN => n6035);
   U23144 : OAI22_X1 port map( A1 => n25496, A2 => n19919, B1 => n25845, B2 => 
                           n25488, ZN => n6036);
   U23145 : OAI22_X1 port map( A1 => n25496, A2 => n19918, B1 => n25848, B2 => 
                           n25488, ZN => n6037);
   U23146 : OAI22_X1 port map( A1 => n25496, A2 => n19917, B1 => n25851, B2 => 
                           n25488, ZN => n6038);
   U23147 : OAI22_X1 port map( A1 => n25496, A2 => n19916, B1 => n25854, B2 => 
                           n25489, ZN => n6039);
   U23148 : OAI22_X1 port map( A1 => n25497, A2 => n19915, B1 => n25857, B2 => 
                           n25489, ZN => n6040);
   U23149 : OAI22_X1 port map( A1 => n25497, A2 => n19914, B1 => n25860, B2 => 
                           n25489, ZN => n6041);
   U23150 : OAI22_X1 port map( A1 => n25497, A2 => n19913, B1 => n25863, B2 => 
                           n25489, ZN => n6042);
   U23151 : OAI22_X1 port map( A1 => n25497, A2 => n19912, B1 => n25866, B2 => 
                           n25489, ZN => n6043);
   U23152 : OAI22_X1 port map( A1 => n25497, A2 => n19911, B1 => n25869, B2 => 
                           n25489, ZN => n6044);
   U23153 : OAI22_X1 port map( A1 => n25497, A2 => n19910, B1 => n25872, B2 => 
                           n25489, ZN => n6045);
   U23154 : OAI22_X1 port map( A1 => n25497, A2 => n19909, B1 => n25875, B2 => 
                           n25489, ZN => n6046);
   U23155 : OAI22_X1 port map( A1 => n25497, A2 => n19908, B1 => n25878, B2 => 
                           n25489, ZN => n6047);
   U23156 : OAI22_X1 port map( A1 => n25497, A2 => n19907, B1 => n25881, B2 => 
                           n25489, ZN => n6048);
   U23157 : OAI22_X1 port map( A1 => n25497, A2 => n19906, B1 => n25884, B2 => 
                           n25489, ZN => n6049);
   U23158 : OAI22_X1 port map( A1 => n25497, A2 => n19905, B1 => n25887, B2 => 
                           n25489, ZN => n6050);
   U23159 : OAI22_X1 port map( A1 => n25497, A2 => n19904, B1 => n25890, B2 => 
                           n25490, ZN => n6051);
   U23160 : OAI22_X1 port map( A1 => n25497, A2 => n19903, B1 => n25893, B2 => 
                           n25490, ZN => n6052);
   U23161 : OAI22_X1 port map( A1 => n25498, A2 => n19902, B1 => n25896, B2 => 
                           n25490, ZN => n6053);
   U23162 : OAI22_X1 port map( A1 => n25498, A2 => n19901, B1 => n25899, B2 => 
                           n25490, ZN => n6054);
   U23163 : OAI22_X1 port map( A1 => n25498, A2 => n19900, B1 => n25902, B2 => 
                           n25490, ZN => n6055);
   U23164 : OAI22_X1 port map( A1 => n25498, A2 => n19899, B1 => n25905, B2 => 
                           n25490, ZN => n6056);
   U23165 : OAI22_X1 port map( A1 => n25498, A2 => n19898, B1 => n25908, B2 => 
                           n25490, ZN => n6057);
   U23166 : OAI22_X1 port map( A1 => n25498, A2 => n19897, B1 => n25911, B2 => 
                           n25490, ZN => n6058);
   U23167 : OAI22_X1 port map( A1 => n25498, A2 => n19896, B1 => n25914, B2 => 
                           n25490, ZN => n6059);
   U23168 : OAI22_X1 port map( A1 => n25498, A2 => n19895, B1 => n25917, B2 => 
                           n25490, ZN => n6060);
   U23169 : OAI22_X1 port map( A1 => n25498, A2 => n19894, B1 => n25920, B2 => 
                           n25490, ZN => n6061);
   U23170 : OAI22_X1 port map( A1 => n25498, A2 => n19893, B1 => n25923, B2 => 
                           n25490, ZN => n6062);
   U23171 : OAI22_X1 port map( A1 => n25498, A2 => n19892, B1 => n25926, B2 => 
                           n25491, ZN => n6063);
   U23172 : OAI22_X1 port map( A1 => n25498, A2 => n19891, B1 => n25929, B2 => 
                           n25491, ZN => n6064);
   U23173 : OAI22_X1 port map( A1 => n25498, A2 => n19890, B1 => n25932, B2 => 
                           n25491, ZN => n6065);
   U23174 : OAI22_X1 port map( A1 => n25499, A2 => n19889, B1 => n25935, B2 => 
                           n25491, ZN => n6066);
   U23175 : OAI22_X1 port map( A1 => n25499, A2 => n19888, B1 => n25938, B2 => 
                           n25491, ZN => n6067);
   U23176 : OAI22_X1 port map( A1 => n25499, A2 => n19887, B1 => n25941, B2 => 
                           n25491, ZN => n6068);
   U23177 : OAI22_X1 port map( A1 => n25499, A2 => n19886, B1 => n25944, B2 => 
                           n25491, ZN => n6069);
   U23178 : OAI22_X1 port map( A1 => n25499, A2 => n19885, B1 => n25947, B2 => 
                           n25491, ZN => n6070);
   U23179 : OAI22_X1 port map( A1 => n25499, A2 => n19884, B1 => n25950, B2 => 
                           n25491, ZN => n6071);
   U23180 : OAI22_X1 port map( A1 => n25499, A2 => n19883, B1 => n25953, B2 => 
                           n25491, ZN => n6072);
   U23181 : OAI22_X1 port map( A1 => n25499, A2 => n19882, B1 => n25956, B2 => 
                           n25491, ZN => n6073);
   U23182 : OAI22_X1 port map( A1 => n25499, A2 => n19881, B1 => n25959, B2 => 
                           n25491, ZN => n6074);
   U23183 : OAI22_X1 port map( A1 => n25700, A2 => n19685, B1 => n25781, B2 => 
                           n25692, ZN => n7039);
   U23184 : OAI22_X1 port map( A1 => n25700, A2 => n19684, B1 => n25784, B2 => 
                           n25692, ZN => n7040);
   U23185 : OAI22_X1 port map( A1 => n25700, A2 => n19683, B1 => n25787, B2 => 
                           n25692, ZN => n7041);
   U23186 : OAI22_X1 port map( A1 => n25700, A2 => n19682, B1 => n25790, B2 => 
                           n25692, ZN => n7042);
   U23187 : OAI22_X1 port map( A1 => n25700, A2 => n19681, B1 => n25793, B2 => 
                           n25692, ZN => n7043);
   U23188 : OAI22_X1 port map( A1 => n25700, A2 => n19680, B1 => n25796, B2 => 
                           n25692, ZN => n7044);
   U23189 : OAI22_X1 port map( A1 => n25700, A2 => n19679, B1 => n25799, B2 => 
                           n25692, ZN => n7045);
   U23190 : OAI22_X1 port map( A1 => n25700, A2 => n19678, B1 => n25802, B2 => 
                           n25692, ZN => n7046);
   U23191 : OAI22_X1 port map( A1 => n25700, A2 => n19677, B1 => n25805, B2 => 
                           n25692, ZN => n7047);
   U23192 : OAI22_X1 port map( A1 => n25700, A2 => n19676, B1 => n25808, B2 => 
                           n25692, ZN => n7048);
   U23193 : OAI22_X1 port map( A1 => n25700, A2 => n19675, B1 => n25811, B2 => 
                           n25692, ZN => n7049);
   U23194 : OAI22_X1 port map( A1 => n25700, A2 => n19674, B1 => n25814, B2 => 
                           n25692, ZN => n7050);
   U23195 : OAI22_X1 port map( A1 => n25701, A2 => n19673, B1 => n25817, B2 => 
                           n25693, ZN => n7051);
   U23196 : OAI22_X1 port map( A1 => n25701, A2 => n19672, B1 => n25820, B2 => 
                           n25693, ZN => n7052);
   U23197 : OAI22_X1 port map( A1 => n25701, A2 => n19671, B1 => n25823, B2 => 
                           n25693, ZN => n7053);
   U23198 : OAI22_X1 port map( A1 => n25701, A2 => n19670, B1 => n25826, B2 => 
                           n25693, ZN => n7054);
   U23199 : OAI22_X1 port map( A1 => n25701, A2 => n19669, B1 => n25829, B2 => 
                           n25693, ZN => n7055);
   U23200 : OAI22_X1 port map( A1 => n25701, A2 => n19668, B1 => n25832, B2 => 
                           n25693, ZN => n7056);
   U23201 : OAI22_X1 port map( A1 => n25701, A2 => n19667, B1 => n25835, B2 => 
                           n25693, ZN => n7057);
   U23202 : OAI22_X1 port map( A1 => n25701, A2 => n19666, B1 => n25838, B2 => 
                           n25693, ZN => n7058);
   U23203 : OAI22_X1 port map( A1 => n25701, A2 => n19665, B1 => n25841, B2 => 
                           n25693, ZN => n7059);
   U23204 : OAI22_X1 port map( A1 => n25701, A2 => n19664, B1 => n25844, B2 => 
                           n25693, ZN => n7060);
   U23205 : OAI22_X1 port map( A1 => n25701, A2 => n19663, B1 => n25847, B2 => 
                           n25693, ZN => n7061);
   U23206 : OAI22_X1 port map( A1 => n25701, A2 => n19662, B1 => n25850, B2 => 
                           n25693, ZN => n7062);
   U23207 : OAI22_X1 port map( A1 => n25701, A2 => n19661, B1 => n25853, B2 => 
                           n25694, ZN => n7063);
   U23208 : OAI22_X1 port map( A1 => n25702, A2 => n19660, B1 => n25856, B2 => 
                           n25694, ZN => n7064);
   U23209 : OAI22_X1 port map( A1 => n25702, A2 => n19659, B1 => n25859, B2 => 
                           n25694, ZN => n7065);
   U23210 : OAI22_X1 port map( A1 => n25702, A2 => n19658, B1 => n25862, B2 => 
                           n25694, ZN => n7066);
   U23211 : OAI22_X1 port map( A1 => n25702, A2 => n19657, B1 => n25865, B2 => 
                           n25694, ZN => n7067);
   U23212 : OAI22_X1 port map( A1 => n25702, A2 => n19656, B1 => n25868, B2 => 
                           n25694, ZN => n7068);
   U23213 : OAI22_X1 port map( A1 => n25702, A2 => n19655, B1 => n25871, B2 => 
                           n25694, ZN => n7069);
   U23214 : OAI22_X1 port map( A1 => n25702, A2 => n19654, B1 => n25874, B2 => 
                           n25694, ZN => n7070);
   U23215 : OAI22_X1 port map( A1 => n25702, A2 => n19653, B1 => n25877, B2 => 
                           n25694, ZN => n7071);
   U23216 : OAI22_X1 port map( A1 => n25702, A2 => n19652, B1 => n25880, B2 => 
                           n25694, ZN => n7072);
   U23217 : OAI22_X1 port map( A1 => n25702, A2 => n19651, B1 => n25883, B2 => 
                           n25694, ZN => n7073);
   U23218 : OAI22_X1 port map( A1 => n25702, A2 => n19650, B1 => n25886, B2 => 
                           n25694, ZN => n7074);
   U23219 : OAI22_X1 port map( A1 => n25702, A2 => n19649, B1 => n25889, B2 => 
                           n25695, ZN => n7075);
   U23220 : OAI22_X1 port map( A1 => n25702, A2 => n19648, B1 => n25892, B2 => 
                           n25695, ZN => n7076);
   U23221 : OAI22_X1 port map( A1 => n25703, A2 => n19647, B1 => n25895, B2 => 
                           n25695, ZN => n7077);
   U23222 : OAI22_X1 port map( A1 => n25703, A2 => n19646, B1 => n25898, B2 => 
                           n25695, ZN => n7078);
   U23223 : OAI22_X1 port map( A1 => n25703, A2 => n19645, B1 => n25901, B2 => 
                           n25695, ZN => n7079);
   U23224 : OAI22_X1 port map( A1 => n25703, A2 => n19644, B1 => n25904, B2 => 
                           n25695, ZN => n7080);
   U23225 : OAI22_X1 port map( A1 => n25703, A2 => n19643, B1 => n25907, B2 => 
                           n25695, ZN => n7081);
   U23226 : OAI22_X1 port map( A1 => n25703, A2 => n19642, B1 => n25910, B2 => 
                           n25695, ZN => n7082);
   U23227 : OAI22_X1 port map( A1 => n25703, A2 => n19641, B1 => n25913, B2 => 
                           n25695, ZN => n7083);
   U23228 : OAI22_X1 port map( A1 => n25703, A2 => n19640, B1 => n25916, B2 => 
                           n25695, ZN => n7084);
   U23229 : OAI22_X1 port map( A1 => n25703, A2 => n19639, B1 => n25919, B2 => 
                           n25695, ZN => n7085);
   U23230 : OAI22_X1 port map( A1 => n25703, A2 => n19638, B1 => n25922, B2 => 
                           n25695, ZN => n7086);
   U23231 : OAI22_X1 port map( A1 => n25703, A2 => n19637, B1 => n25925, B2 => 
                           n25696, ZN => n7087);
   U23232 : OAI22_X1 port map( A1 => n25703, A2 => n19636, B1 => n25928, B2 => 
                           n25696, ZN => n7088);
   U23233 : OAI22_X1 port map( A1 => n25703, A2 => n19635, B1 => n25931, B2 => 
                           n25696, ZN => n7089);
   U23234 : OAI22_X1 port map( A1 => n25704, A2 => n19634, B1 => n25934, B2 => 
                           n25696, ZN => n7090);
   U23235 : OAI22_X1 port map( A1 => n25704, A2 => n19633, B1 => n25937, B2 => 
                           n25696, ZN => n7091);
   U23236 : OAI22_X1 port map( A1 => n25704, A2 => n19632, B1 => n25940, B2 => 
                           n25696, ZN => n7092);
   U23237 : OAI22_X1 port map( A1 => n25704, A2 => n19631, B1 => n25943, B2 => 
                           n25696, ZN => n7093);
   U23238 : OAI22_X1 port map( A1 => n25704, A2 => n19630, B1 => n25946, B2 => 
                           n25696, ZN => n7094);
   U23239 : OAI22_X1 port map( A1 => n25704, A2 => n19629, B1 => n25949, B2 => 
                           n25696, ZN => n7095);
   U23240 : OAI22_X1 port map( A1 => n25704, A2 => n19628, B1 => n25952, B2 => 
                           n25696, ZN => n7096);
   U23241 : OAI22_X1 port map( A1 => n25704, A2 => n19627, B1 => n25955, B2 => 
                           n25696, ZN => n7097);
   U23242 : OAI22_X1 port map( A1 => n25704, A2 => n19626, B1 => n25958, B2 => 
                           n25696, ZN => n7098);
   U23243 : NAND2_X1 port map( A1 => n22753, A2 => n22754, ZN => n5374);
   U23244 : NOR4_X1 port map( A1 => n22780, A2 => n22781, A3 => n22782, A4 => 
                           n22783, ZN => n22753);
   U23245 : NOR4_X1 port map( A1 => n22755, A2 => n22756, A3 => n22757, A4 => 
                           n22758, ZN => n22754);
   U23246 : OAI221_X1 port map( B1 => n20710, B2 => n24997, C1 => n8967, C2 => 
                           n24991, A => n22801, ZN => n22780);
   U23247 : NAND2_X1 port map( A1 => n22840, A2 => n22841, ZN => n5371);
   U23248 : NOR4_X1 port map( A1 => n22850, A2 => n22851, A3 => n22852, A4 => 
                           n22853, ZN => n22840);
   U23249 : NOR4_X1 port map( A1 => n22842, A2 => n22843, A3 => n22844, A4 => 
                           n22845, ZN => n22841);
   U23250 : OAI221_X1 port map( B1 => n20713, B2 => n24997, C1 => n8970, C2 => 
                           n24991, A => n22857, ZN => n22850);
   U23251 : NAND2_X1 port map( A1 => n22822, A2 => n22823, ZN => n5372);
   U23252 : NOR4_X1 port map( A1 => n22832, A2 => n22833, A3 => n22834, A4 => 
                           n22835, ZN => n22822);
   U23253 : NOR4_X1 port map( A1 => n22824, A2 => n22825, A3 => n22826, A4 => 
                           n22827, ZN => n22823);
   U23254 : OAI221_X1 port map( B1 => n20712, B2 => n24997, C1 => n8969, C2 => 
                           n24991, A => n22839, ZN => n22832);
   U23255 : NAND2_X1 port map( A1 => n22804, A2 => n22805, ZN => n5373);
   U23256 : NOR4_X1 port map( A1 => n22814, A2 => n22815, A3 => n22816, A4 => 
                           n22817, ZN => n22804);
   U23257 : NOR4_X1 port map( A1 => n22806, A2 => n22807, A3 => n22808, A4 => 
                           n22809, ZN => n22805);
   U23258 : OAI221_X1 port map( B1 => n20711, B2 => n24997, C1 => n8968, C2 => 
                           n24991, A => n22821, ZN => n22814);
   U23259 : NAND2_X1 port map( A1 => n21643, A2 => n21644, ZN => n5435);
   U23260 : NOR4_X1 port map( A1 => n21653, A2 => n21654, A3 => n21655, A4 => 
                           n21656, ZN => n21643);
   U23261 : NOR4_X1 port map( A1 => n21645, A2 => n21646, A3 => n21647, A4 => 
                           n21648, ZN => n21644);
   U23262 : OAI221_X1 port map( B1 => n20713, B2 => n25195, C1 => n8970, C2 => 
                           n25189, A => n21660, ZN => n21653);
   U23263 : NAND2_X1 port map( A1 => n21625, A2 => n21626, ZN => n5436);
   U23264 : NOR4_X1 port map( A1 => n21635, A2 => n21636, A3 => n21637, A4 => 
                           n21638, ZN => n21625);
   U23265 : NOR4_X1 port map( A1 => n21627, A2 => n21628, A3 => n21629, A4 => 
                           n21630, ZN => n21626);
   U23266 : OAI221_X1 port map( B1 => n20712, B2 => n25195, C1 => n8969, C2 => 
                           n25189, A => n21642, ZN => n21635);
   U23267 : NAND2_X1 port map( A1 => n21607, A2 => n21608, ZN => n5437);
   U23268 : NOR4_X1 port map( A1 => n21617, A2 => n21618, A3 => n21619, A4 => 
                           n21620, ZN => n21607);
   U23269 : NOR4_X1 port map( A1 => n21609, A2 => n21610, A3 => n21611, A4 => 
                           n21612, ZN => n21608);
   U23270 : OAI221_X1 port map( B1 => n20711, B2 => n25195, C1 => n8968, C2 => 
                           n25189, A => n21624, ZN => n21617);
   U23271 : NAND2_X1 port map( A1 => n21556, A2 => n21557, ZN => n5438);
   U23272 : NOR4_X1 port map( A1 => n21583, A2 => n21584, A3 => n21585, A4 => 
                           n21586, ZN => n21556);
   U23273 : NOR4_X1 port map( A1 => n21558, A2 => n21559, A3 => n21560, A4 => 
                           n21561, ZN => n21557);
   U23274 : OAI221_X1 port map( B1 => n20710, B2 => n25195, C1 => n8967, C2 => 
                           n25189, A => n21604, ZN => n21583);
   U23275 : NAND2_X1 port map( A1 => n23920, A2 => n23921, ZN => n5311);
   U23276 : NOR4_X1 port map( A1 => n23941, A2 => n23942, A3 => n23943, A4 => 
                           n23944, ZN => n23920);
   U23277 : NOR4_X1 port map( A1 => n23922, A2 => n23923, A3 => n23924, A4 => 
                           n23925, ZN => n23921);
   U23278 : OAI221_X1 port map( B1 => n20773, B2 => n24992, C1 => n9030, C2 => 
                           n24986, A => n23949, ZN => n23941);
   U23279 : NAND2_X1 port map( A1 => n23902, A2 => n23903, ZN => n5312);
   U23280 : NOR4_X1 port map( A1 => n23912, A2 => n23913, A3 => n23914, A4 => 
                           n23915, ZN => n23902);
   U23281 : NOR4_X1 port map( A1 => n23904, A2 => n23905, A3 => n23906, A4 => 
                           n23907, ZN => n23903);
   U23282 : OAI221_X1 port map( B1 => n20772, B2 => n24992, C1 => n9029, C2 => 
                           n24986, A => n23919, ZN => n23912);
   U23283 : NAND2_X1 port map( A1 => n23884, A2 => n23885, ZN => n5313);
   U23284 : NOR4_X1 port map( A1 => n23894, A2 => n23895, A3 => n23896, A4 => 
                           n23897, ZN => n23884);
   U23285 : NOR4_X1 port map( A1 => n23886, A2 => n23887, A3 => n23888, A4 => 
                           n23889, ZN => n23885);
   U23286 : OAI221_X1 port map( B1 => n20771, B2 => n24992, C1 => n9028, C2 => 
                           n24986, A => n23901, ZN => n23894);
   U23287 : NAND2_X1 port map( A1 => n23866, A2 => n23867, ZN => n5314);
   U23288 : NOR4_X1 port map( A1 => n23876, A2 => n23877, A3 => n23878, A4 => 
                           n23879, ZN => n23866);
   U23289 : NOR4_X1 port map( A1 => n23868, A2 => n23869, A3 => n23870, A4 => 
                           n23871, ZN => n23867);
   U23290 : OAI221_X1 port map( B1 => n20770, B2 => n24992, C1 => n9027, C2 => 
                           n24986, A => n23883, ZN => n23876);
   U23291 : NAND2_X1 port map( A1 => n23848, A2 => n23849, ZN => n5315);
   U23292 : NOR4_X1 port map( A1 => n23858, A2 => n23859, A3 => n23860, A4 => 
                           n23861, ZN => n23848);
   U23293 : NOR4_X1 port map( A1 => n23850, A2 => n23851, A3 => n23852, A4 => 
                           n23853, ZN => n23849);
   U23294 : OAI221_X1 port map( B1 => n20769, B2 => n24992, C1 => n9026, C2 => 
                           n24986, A => n23865, ZN => n23858);
   U23295 : NAND2_X1 port map( A1 => n23830, A2 => n23831, ZN => n5316);
   U23296 : NOR4_X1 port map( A1 => n23840, A2 => n23841, A3 => n23842, A4 => 
                           n23843, ZN => n23830);
   U23297 : NOR4_X1 port map( A1 => n23832, A2 => n23833, A3 => n23834, A4 => 
                           n23835, ZN => n23831);
   U23298 : OAI221_X1 port map( B1 => n20768, B2 => n24992, C1 => n9025, C2 => 
                           n24986, A => n23847, ZN => n23840);
   U23299 : NAND2_X1 port map( A1 => n23812, A2 => n23813, ZN => n5317);
   U23300 : NOR4_X1 port map( A1 => n23822, A2 => n23823, A3 => n23824, A4 => 
                           n23825, ZN => n23812);
   U23301 : NOR4_X1 port map( A1 => n23814, A2 => n23815, A3 => n23816, A4 => 
                           n23817, ZN => n23813);
   U23302 : OAI221_X1 port map( B1 => n20767, B2 => n24992, C1 => n9024, C2 => 
                           n24986, A => n23829, ZN => n23822);
   U23303 : NAND2_X1 port map( A1 => n23794, A2 => n23795, ZN => n5318);
   U23304 : NOR4_X1 port map( A1 => n23804, A2 => n23805, A3 => n23806, A4 => 
                           n23807, ZN => n23794);
   U23305 : NOR4_X1 port map( A1 => n23796, A2 => n23797, A3 => n23798, A4 => 
                           n23799, ZN => n23795);
   U23306 : OAI221_X1 port map( B1 => n20766, B2 => n24992, C1 => n9023, C2 => 
                           n24986, A => n23811, ZN => n23804);
   U23307 : NAND2_X1 port map( A1 => n23776, A2 => n23777, ZN => n5319);
   U23308 : NOR4_X1 port map( A1 => n23786, A2 => n23787, A3 => n23788, A4 => 
                           n23789, ZN => n23776);
   U23309 : NOR4_X1 port map( A1 => n23778, A2 => n23779, A3 => n23780, A4 => 
                           n23781, ZN => n23777);
   U23310 : OAI221_X1 port map( B1 => n20765, B2 => n24992, C1 => n9022, C2 => 
                           n24986, A => n23793, ZN => n23786);
   U23311 : NAND2_X1 port map( A1 => n23758, A2 => n23759, ZN => n5320);
   U23312 : NOR4_X1 port map( A1 => n23768, A2 => n23769, A3 => n23770, A4 => 
                           n23771, ZN => n23758);
   U23313 : NOR4_X1 port map( A1 => n23760, A2 => n23761, A3 => n23762, A4 => 
                           n23763, ZN => n23759);
   U23314 : OAI221_X1 port map( B1 => n20764, B2 => n24992, C1 => n9021, C2 => 
                           n24986, A => n23775, ZN => n23768);
   U23315 : NAND2_X1 port map( A1 => n23740, A2 => n23741, ZN => n5321);
   U23316 : NOR4_X1 port map( A1 => n23750, A2 => n23751, A3 => n23752, A4 => 
                           n23753, ZN => n23740);
   U23317 : NOR4_X1 port map( A1 => n23742, A2 => n23743, A3 => n23744, A4 => 
                           n23745, ZN => n23741);
   U23318 : OAI221_X1 port map( B1 => n20763, B2 => n24992, C1 => n9020, C2 => 
                           n24986, A => n23757, ZN => n23750);
   U23319 : NAND2_X1 port map( A1 => n23722, A2 => n23723, ZN => n5322);
   U23320 : NOR4_X1 port map( A1 => n23732, A2 => n23733, A3 => n23734, A4 => 
                           n23735, ZN => n23722);
   U23321 : NOR4_X1 port map( A1 => n23724, A2 => n23725, A3 => n23726, A4 => 
                           n23727, ZN => n23723);
   U23322 : OAI221_X1 port map( B1 => n20762, B2 => n24992, C1 => n9019, C2 => 
                           n24986, A => n23739, ZN => n23732);
   U23323 : NAND2_X1 port map( A1 => n23704, A2 => n23705, ZN => n5323);
   U23324 : NOR4_X1 port map( A1 => n23714, A2 => n23715, A3 => n23716, A4 => 
                           n23717, ZN => n23704);
   U23325 : NOR4_X1 port map( A1 => n23706, A2 => n23707, A3 => n23708, A4 => 
                           n23709, ZN => n23705);
   U23326 : OAI221_X1 port map( B1 => n20761, B2 => n24993, C1 => n9018, C2 => 
                           n24987, A => n23721, ZN => n23714);
   U23327 : NAND2_X1 port map( A1 => n23686, A2 => n23687, ZN => n5324);
   U23328 : NOR4_X1 port map( A1 => n23696, A2 => n23697, A3 => n23698, A4 => 
                           n23699, ZN => n23686);
   U23329 : NOR4_X1 port map( A1 => n23688, A2 => n23689, A3 => n23690, A4 => 
                           n23691, ZN => n23687);
   U23330 : OAI221_X1 port map( B1 => n20760, B2 => n24993, C1 => n9017, C2 => 
                           n24987, A => n23703, ZN => n23696);
   U23331 : NAND2_X1 port map( A1 => n23668, A2 => n23669, ZN => n5325);
   U23332 : NOR4_X1 port map( A1 => n23678, A2 => n23679, A3 => n23680, A4 => 
                           n23681, ZN => n23668);
   U23333 : NOR4_X1 port map( A1 => n23670, A2 => n23671, A3 => n23672, A4 => 
                           n23673, ZN => n23669);
   U23334 : OAI221_X1 port map( B1 => n20759, B2 => n24993, C1 => n9016, C2 => 
                           n24987, A => n23685, ZN => n23678);
   U23335 : NAND2_X1 port map( A1 => n23650, A2 => n23651, ZN => n5326);
   U23336 : NOR4_X1 port map( A1 => n23660, A2 => n23661, A3 => n23662, A4 => 
                           n23663, ZN => n23650);
   U23337 : NOR4_X1 port map( A1 => n23652, A2 => n23653, A3 => n23654, A4 => 
                           n23655, ZN => n23651);
   U23338 : OAI221_X1 port map( B1 => n20758, B2 => n24993, C1 => n9015, C2 => 
                           n24987, A => n23667, ZN => n23660);
   U23339 : NAND2_X1 port map( A1 => n23632, A2 => n23633, ZN => n5327);
   U23340 : NOR4_X1 port map( A1 => n23642, A2 => n23643, A3 => n23644, A4 => 
                           n23645, ZN => n23632);
   U23341 : NOR4_X1 port map( A1 => n23634, A2 => n23635, A3 => n23636, A4 => 
                           n23637, ZN => n23633);
   U23342 : OAI221_X1 port map( B1 => n20757, B2 => n24993, C1 => n9014, C2 => 
                           n24987, A => n23649, ZN => n23642);
   U23343 : NAND2_X1 port map( A1 => n23614, A2 => n23615, ZN => n5328);
   U23344 : NOR4_X1 port map( A1 => n23624, A2 => n23625, A3 => n23626, A4 => 
                           n23627, ZN => n23614);
   U23345 : NOR4_X1 port map( A1 => n23616, A2 => n23617, A3 => n23618, A4 => 
                           n23619, ZN => n23615);
   U23346 : OAI221_X1 port map( B1 => n20756, B2 => n24993, C1 => n9013, C2 => 
                           n24987, A => n23631, ZN => n23624);
   U23347 : NAND2_X1 port map( A1 => n23596, A2 => n23597, ZN => n5329);
   U23348 : NOR4_X1 port map( A1 => n23606, A2 => n23607, A3 => n23608, A4 => 
                           n23609, ZN => n23596);
   U23349 : NOR4_X1 port map( A1 => n23598, A2 => n23599, A3 => n23600, A4 => 
                           n23601, ZN => n23597);
   U23350 : OAI221_X1 port map( B1 => n20755, B2 => n24993, C1 => n9012, C2 => 
                           n24987, A => n23613, ZN => n23606);
   U23351 : NAND2_X1 port map( A1 => n23578, A2 => n23579, ZN => n5330);
   U23352 : NOR4_X1 port map( A1 => n23588, A2 => n23589, A3 => n23590, A4 => 
                           n23591, ZN => n23578);
   U23353 : NOR4_X1 port map( A1 => n23580, A2 => n23581, A3 => n23582, A4 => 
                           n23583, ZN => n23579);
   U23354 : OAI221_X1 port map( B1 => n20754, B2 => n24993, C1 => n9011, C2 => 
                           n24987, A => n23595, ZN => n23588);
   U23355 : NAND2_X1 port map( A1 => n23560, A2 => n23561, ZN => n5331);
   U23356 : NOR4_X1 port map( A1 => n23570, A2 => n23571, A3 => n23572, A4 => 
                           n23573, ZN => n23560);
   U23357 : NOR4_X1 port map( A1 => n23562, A2 => n23563, A3 => n23564, A4 => 
                           n23565, ZN => n23561);
   U23358 : OAI221_X1 port map( B1 => n20753, B2 => n24993, C1 => n9010, C2 => 
                           n24987, A => n23577, ZN => n23570);
   U23359 : NAND2_X1 port map( A1 => n23542, A2 => n23543, ZN => n5332);
   U23360 : NOR4_X1 port map( A1 => n23552, A2 => n23553, A3 => n23554, A4 => 
                           n23555, ZN => n23542);
   U23361 : NOR4_X1 port map( A1 => n23544, A2 => n23545, A3 => n23546, A4 => 
                           n23547, ZN => n23543);
   U23362 : OAI221_X1 port map( B1 => n20752, B2 => n24993, C1 => n9009, C2 => 
                           n24987, A => n23559, ZN => n23552);
   U23363 : NAND2_X1 port map( A1 => n23524, A2 => n23525, ZN => n5333);
   U23364 : NOR4_X1 port map( A1 => n23534, A2 => n23535, A3 => n23536, A4 => 
                           n23537, ZN => n23524);
   U23365 : NOR4_X1 port map( A1 => n23526, A2 => n23527, A3 => n23528, A4 => 
                           n23529, ZN => n23525);
   U23366 : OAI221_X1 port map( B1 => n20751, B2 => n24993, C1 => n9008, C2 => 
                           n24987, A => n23541, ZN => n23534);
   U23367 : NAND2_X1 port map( A1 => n23506, A2 => n23507, ZN => n5334);
   U23368 : NOR4_X1 port map( A1 => n23516, A2 => n23517, A3 => n23518, A4 => 
                           n23519, ZN => n23506);
   U23369 : NOR4_X1 port map( A1 => n23508, A2 => n23509, A3 => n23510, A4 => 
                           n23511, ZN => n23507);
   U23370 : OAI221_X1 port map( B1 => n20750, B2 => n24993, C1 => n9007, C2 => 
                           n24987, A => n23523, ZN => n23516);
   U23371 : NAND2_X1 port map( A1 => n23488, A2 => n23489, ZN => n5335);
   U23372 : NOR4_X1 port map( A1 => n23498, A2 => n23499, A3 => n23500, A4 => 
                           n23501, ZN => n23488);
   U23373 : NOR4_X1 port map( A1 => n23490, A2 => n23491, A3 => n23492, A4 => 
                           n23493, ZN => n23489);
   U23374 : OAI221_X1 port map( B1 => n20749, B2 => n24994, C1 => n9006, C2 => 
                           n24988, A => n23505, ZN => n23498);
   U23375 : NAND2_X1 port map( A1 => n23470, A2 => n23471, ZN => n5336);
   U23376 : NOR4_X1 port map( A1 => n23480, A2 => n23481, A3 => n23482, A4 => 
                           n23483, ZN => n23470);
   U23377 : NOR4_X1 port map( A1 => n23472, A2 => n23473, A3 => n23474, A4 => 
                           n23475, ZN => n23471);
   U23378 : OAI221_X1 port map( B1 => n20748, B2 => n24994, C1 => n9005, C2 => 
                           n24988, A => n23487, ZN => n23480);
   U23379 : NAND2_X1 port map( A1 => n23452, A2 => n23453, ZN => n5337);
   U23380 : NOR4_X1 port map( A1 => n23462, A2 => n23463, A3 => n23464, A4 => 
                           n23465, ZN => n23452);
   U23381 : NOR4_X1 port map( A1 => n23454, A2 => n23455, A3 => n23456, A4 => 
                           n23457, ZN => n23453);
   U23382 : OAI221_X1 port map( B1 => n20747, B2 => n24994, C1 => n9004, C2 => 
                           n24988, A => n23469, ZN => n23462);
   U23383 : NAND2_X1 port map( A1 => n23434, A2 => n23435, ZN => n5338);
   U23384 : NOR4_X1 port map( A1 => n23444, A2 => n23445, A3 => n23446, A4 => 
                           n23447, ZN => n23434);
   U23385 : NOR4_X1 port map( A1 => n23436, A2 => n23437, A3 => n23438, A4 => 
                           n23439, ZN => n23435);
   U23386 : OAI221_X1 port map( B1 => n20746, B2 => n24994, C1 => n9003, C2 => 
                           n24988, A => n23451, ZN => n23444);
   U23387 : NAND2_X1 port map( A1 => n23416, A2 => n23417, ZN => n5339);
   U23388 : NOR4_X1 port map( A1 => n23426, A2 => n23427, A3 => n23428, A4 => 
                           n23429, ZN => n23416);
   U23389 : NOR4_X1 port map( A1 => n23418, A2 => n23419, A3 => n23420, A4 => 
                           n23421, ZN => n23417);
   U23390 : OAI221_X1 port map( B1 => n20745, B2 => n24994, C1 => n9002, C2 => 
                           n24988, A => n23433, ZN => n23426);
   U23391 : NAND2_X1 port map( A1 => n23398, A2 => n23399, ZN => n5340);
   U23392 : NOR4_X1 port map( A1 => n23408, A2 => n23409, A3 => n23410, A4 => 
                           n23411, ZN => n23398);
   U23393 : NOR4_X1 port map( A1 => n23400, A2 => n23401, A3 => n23402, A4 => 
                           n23403, ZN => n23399);
   U23394 : OAI221_X1 port map( B1 => n20744, B2 => n24994, C1 => n9001, C2 => 
                           n24988, A => n23415, ZN => n23408);
   U23395 : NAND2_X1 port map( A1 => n23380, A2 => n23381, ZN => n5341);
   U23396 : NOR4_X1 port map( A1 => n23390, A2 => n23391, A3 => n23392, A4 => 
                           n23393, ZN => n23380);
   U23397 : NOR4_X1 port map( A1 => n23382, A2 => n23383, A3 => n23384, A4 => 
                           n23385, ZN => n23381);
   U23398 : OAI221_X1 port map( B1 => n20743, B2 => n24994, C1 => n9000, C2 => 
                           n24988, A => n23397, ZN => n23390);
   U23399 : NAND2_X1 port map( A1 => n23362, A2 => n23363, ZN => n5342);
   U23400 : NOR4_X1 port map( A1 => n23372, A2 => n23373, A3 => n23374, A4 => 
                           n23375, ZN => n23362);
   U23401 : NOR4_X1 port map( A1 => n23364, A2 => n23365, A3 => n23366, A4 => 
                           n23367, ZN => n23363);
   U23402 : OAI221_X1 port map( B1 => n20742, B2 => n24994, C1 => n8999, C2 => 
                           n24988, A => n23379, ZN => n23372);
   U23403 : NAND2_X1 port map( A1 => n23344, A2 => n23345, ZN => n5343);
   U23404 : NOR4_X1 port map( A1 => n23354, A2 => n23355, A3 => n23356, A4 => 
                           n23357, ZN => n23344);
   U23405 : NOR4_X1 port map( A1 => n23346, A2 => n23347, A3 => n23348, A4 => 
                           n23349, ZN => n23345);
   U23406 : OAI221_X1 port map( B1 => n20741, B2 => n24994, C1 => n8998, C2 => 
                           n24988, A => n23361, ZN => n23354);
   U23407 : NAND2_X1 port map( A1 => n23326, A2 => n23327, ZN => n5344);
   U23408 : NOR4_X1 port map( A1 => n23336, A2 => n23337, A3 => n23338, A4 => 
                           n23339, ZN => n23326);
   U23409 : NOR4_X1 port map( A1 => n23328, A2 => n23329, A3 => n23330, A4 => 
                           n23331, ZN => n23327);
   U23410 : OAI221_X1 port map( B1 => n20740, B2 => n24994, C1 => n8997, C2 => 
                           n24988, A => n23343, ZN => n23336);
   U23411 : NAND2_X1 port map( A1 => n23308, A2 => n23309, ZN => n5345);
   U23412 : NOR4_X1 port map( A1 => n23318, A2 => n23319, A3 => n23320, A4 => 
                           n23321, ZN => n23308);
   U23413 : NOR4_X1 port map( A1 => n23310, A2 => n23311, A3 => n23312, A4 => 
                           n23313, ZN => n23309);
   U23414 : OAI221_X1 port map( B1 => n20739, B2 => n24994, C1 => n8996, C2 => 
                           n24988, A => n23325, ZN => n23318);
   U23415 : NAND2_X1 port map( A1 => n23290, A2 => n23291, ZN => n5346);
   U23416 : NOR4_X1 port map( A1 => n23300, A2 => n23301, A3 => n23302, A4 => 
                           n23303, ZN => n23290);
   U23417 : NOR4_X1 port map( A1 => n23292, A2 => n23293, A3 => n23294, A4 => 
                           n23295, ZN => n23291);
   U23418 : OAI221_X1 port map( B1 => n20738, B2 => n24994, C1 => n8995, C2 => 
                           n24988, A => n23307, ZN => n23300);
   U23419 : NAND2_X1 port map( A1 => n23272, A2 => n23273, ZN => n5347);
   U23420 : NOR4_X1 port map( A1 => n23282, A2 => n23283, A3 => n23284, A4 => 
                           n23285, ZN => n23272);
   U23421 : NOR4_X1 port map( A1 => n23274, A2 => n23275, A3 => n23276, A4 => 
                           n23277, ZN => n23273);
   U23422 : OAI221_X1 port map( B1 => n20737, B2 => n24995, C1 => n8994, C2 => 
                           n24989, A => n23289, ZN => n23282);
   U23423 : NAND2_X1 port map( A1 => n23254, A2 => n23255, ZN => n5348);
   U23424 : NOR4_X1 port map( A1 => n23264, A2 => n23265, A3 => n23266, A4 => 
                           n23267, ZN => n23254);
   U23425 : NOR4_X1 port map( A1 => n23256, A2 => n23257, A3 => n23258, A4 => 
                           n23259, ZN => n23255);
   U23426 : OAI221_X1 port map( B1 => n20736, B2 => n24995, C1 => n8993, C2 => 
                           n24989, A => n23271, ZN => n23264);
   U23427 : NAND2_X1 port map( A1 => n23236, A2 => n23237, ZN => n5349);
   U23428 : NOR4_X1 port map( A1 => n23246, A2 => n23247, A3 => n23248, A4 => 
                           n23249, ZN => n23236);
   U23429 : NOR4_X1 port map( A1 => n23238, A2 => n23239, A3 => n23240, A4 => 
                           n23241, ZN => n23237);
   U23430 : OAI221_X1 port map( B1 => n20735, B2 => n24995, C1 => n8992, C2 => 
                           n24989, A => n23253, ZN => n23246);
   U23431 : NAND2_X1 port map( A1 => n23218, A2 => n23219, ZN => n5350);
   U23432 : NOR4_X1 port map( A1 => n23228, A2 => n23229, A3 => n23230, A4 => 
                           n23231, ZN => n23218);
   U23433 : NOR4_X1 port map( A1 => n23220, A2 => n23221, A3 => n23222, A4 => 
                           n23223, ZN => n23219);
   U23434 : OAI221_X1 port map( B1 => n20734, B2 => n24995, C1 => n8991, C2 => 
                           n24989, A => n23235, ZN => n23228);
   U23435 : NAND2_X1 port map( A1 => n23200, A2 => n23201, ZN => n5351);
   U23436 : NOR4_X1 port map( A1 => n23210, A2 => n23211, A3 => n23212, A4 => 
                           n23213, ZN => n23200);
   U23437 : NOR4_X1 port map( A1 => n23202, A2 => n23203, A3 => n23204, A4 => 
                           n23205, ZN => n23201);
   U23438 : OAI221_X1 port map( B1 => n20733, B2 => n24995, C1 => n8990, C2 => 
                           n24989, A => n23217, ZN => n23210);
   U23439 : NAND2_X1 port map( A1 => n23182, A2 => n23183, ZN => n5352);
   U23440 : NOR4_X1 port map( A1 => n23192, A2 => n23193, A3 => n23194, A4 => 
                           n23195, ZN => n23182);
   U23441 : NOR4_X1 port map( A1 => n23184, A2 => n23185, A3 => n23186, A4 => 
                           n23187, ZN => n23183);
   U23442 : OAI221_X1 port map( B1 => n20732, B2 => n24995, C1 => n8989, C2 => 
                           n24989, A => n23199, ZN => n23192);
   U23443 : NAND2_X1 port map( A1 => n23164, A2 => n23165, ZN => n5353);
   U23444 : NOR4_X1 port map( A1 => n23174, A2 => n23175, A3 => n23176, A4 => 
                           n23177, ZN => n23164);
   U23445 : NOR4_X1 port map( A1 => n23166, A2 => n23167, A3 => n23168, A4 => 
                           n23169, ZN => n23165);
   U23446 : OAI221_X1 port map( B1 => n20731, B2 => n24995, C1 => n8988, C2 => 
                           n24989, A => n23181, ZN => n23174);
   U23447 : NAND2_X1 port map( A1 => n23146, A2 => n23147, ZN => n5354);
   U23448 : NOR4_X1 port map( A1 => n23156, A2 => n23157, A3 => n23158, A4 => 
                           n23159, ZN => n23146);
   U23449 : NOR4_X1 port map( A1 => n23148, A2 => n23149, A3 => n23150, A4 => 
                           n23151, ZN => n23147);
   U23450 : OAI221_X1 port map( B1 => n20730, B2 => n24995, C1 => n8987, C2 => 
                           n24989, A => n23163, ZN => n23156);
   U23451 : NAND2_X1 port map( A1 => n23128, A2 => n23129, ZN => n5355);
   U23452 : NOR4_X1 port map( A1 => n23138, A2 => n23139, A3 => n23140, A4 => 
                           n23141, ZN => n23128);
   U23453 : NOR4_X1 port map( A1 => n23130, A2 => n23131, A3 => n23132, A4 => 
                           n23133, ZN => n23129);
   U23454 : OAI221_X1 port map( B1 => n20729, B2 => n24995, C1 => n8986, C2 => 
                           n24989, A => n23145, ZN => n23138);
   U23455 : NAND2_X1 port map( A1 => n23110, A2 => n23111, ZN => n5356);
   U23456 : NOR4_X1 port map( A1 => n23120, A2 => n23121, A3 => n23122, A4 => 
                           n23123, ZN => n23110);
   U23457 : NOR4_X1 port map( A1 => n23112, A2 => n23113, A3 => n23114, A4 => 
                           n23115, ZN => n23111);
   U23458 : OAI221_X1 port map( B1 => n20728, B2 => n24995, C1 => n8985, C2 => 
                           n24989, A => n23127, ZN => n23120);
   U23459 : NAND2_X1 port map( A1 => n23092, A2 => n23093, ZN => n5357);
   U23460 : NOR4_X1 port map( A1 => n23102, A2 => n23103, A3 => n23104, A4 => 
                           n23105, ZN => n23092);
   U23461 : NOR4_X1 port map( A1 => n23094, A2 => n23095, A3 => n23096, A4 => 
                           n23097, ZN => n23093);
   U23462 : OAI221_X1 port map( B1 => n20727, B2 => n24995, C1 => n8984, C2 => 
                           n24989, A => n23109, ZN => n23102);
   U23463 : NAND2_X1 port map( A1 => n23074, A2 => n23075, ZN => n5358);
   U23464 : NOR4_X1 port map( A1 => n23084, A2 => n23085, A3 => n23086, A4 => 
                           n23087, ZN => n23074);
   U23465 : NOR4_X1 port map( A1 => n23076, A2 => n23077, A3 => n23078, A4 => 
                           n23079, ZN => n23075);
   U23466 : OAI221_X1 port map( B1 => n20726, B2 => n24995, C1 => n8983, C2 => 
                           n24989, A => n23091, ZN => n23084);
   U23467 : NAND2_X1 port map( A1 => n23056, A2 => n23057, ZN => n5359);
   U23468 : NOR4_X1 port map( A1 => n23066, A2 => n23067, A3 => n23068, A4 => 
                           n23069, ZN => n23056);
   U23469 : NOR4_X1 port map( A1 => n23058, A2 => n23059, A3 => n23060, A4 => 
                           n23061, ZN => n23057);
   U23470 : OAI221_X1 port map( B1 => n20725, B2 => n24996, C1 => n8982, C2 => 
                           n24990, A => n23073, ZN => n23066);
   U23471 : NAND2_X1 port map( A1 => n23038, A2 => n23039, ZN => n5360);
   U23472 : NOR4_X1 port map( A1 => n23048, A2 => n23049, A3 => n23050, A4 => 
                           n23051, ZN => n23038);
   U23473 : NOR4_X1 port map( A1 => n23040, A2 => n23041, A3 => n23042, A4 => 
                           n23043, ZN => n23039);
   U23474 : OAI221_X1 port map( B1 => n20724, B2 => n24996, C1 => n8981, C2 => 
                           n24990, A => n23055, ZN => n23048);
   U23475 : NAND2_X1 port map( A1 => n23020, A2 => n23021, ZN => n5361);
   U23476 : NOR4_X1 port map( A1 => n23030, A2 => n23031, A3 => n23032, A4 => 
                           n23033, ZN => n23020);
   U23477 : NOR4_X1 port map( A1 => n23022, A2 => n23023, A3 => n23024, A4 => 
                           n23025, ZN => n23021);
   U23478 : OAI221_X1 port map( B1 => n20723, B2 => n24996, C1 => n8980, C2 => 
                           n24990, A => n23037, ZN => n23030);
   U23479 : NAND2_X1 port map( A1 => n23002, A2 => n23003, ZN => n5362);
   U23480 : NOR4_X1 port map( A1 => n23012, A2 => n23013, A3 => n23014, A4 => 
                           n23015, ZN => n23002);
   U23481 : NOR4_X1 port map( A1 => n23004, A2 => n23005, A3 => n23006, A4 => 
                           n23007, ZN => n23003);
   U23482 : OAI221_X1 port map( B1 => n20722, B2 => n24996, C1 => n8979, C2 => 
                           n24990, A => n23019, ZN => n23012);
   U23483 : NAND2_X1 port map( A1 => n22984, A2 => n22985, ZN => n5363);
   U23484 : NOR4_X1 port map( A1 => n22994, A2 => n22995, A3 => n22996, A4 => 
                           n22997, ZN => n22984);
   U23485 : NOR4_X1 port map( A1 => n22986, A2 => n22987, A3 => n22988, A4 => 
                           n22989, ZN => n22985);
   U23486 : OAI221_X1 port map( B1 => n20721, B2 => n24996, C1 => n8978, C2 => 
                           n24990, A => n23001, ZN => n22994);
   U23487 : NAND2_X1 port map( A1 => n22966, A2 => n22967, ZN => n5364);
   U23488 : NOR4_X1 port map( A1 => n22976, A2 => n22977, A3 => n22978, A4 => 
                           n22979, ZN => n22966);
   U23489 : NOR4_X1 port map( A1 => n22968, A2 => n22969, A3 => n22970, A4 => 
                           n22971, ZN => n22967);
   U23490 : OAI221_X1 port map( B1 => n20720, B2 => n24996, C1 => n8977, C2 => 
                           n24990, A => n22983, ZN => n22976);
   U23491 : NAND2_X1 port map( A1 => n22948, A2 => n22949, ZN => n5365);
   U23492 : NOR4_X1 port map( A1 => n22958, A2 => n22959, A3 => n22960, A4 => 
                           n22961, ZN => n22948);
   U23493 : NOR4_X1 port map( A1 => n22950, A2 => n22951, A3 => n22952, A4 => 
                           n22953, ZN => n22949);
   U23494 : OAI221_X1 port map( B1 => n20719, B2 => n24996, C1 => n8976, C2 => 
                           n24990, A => n22965, ZN => n22958);
   U23495 : NAND2_X1 port map( A1 => n22930, A2 => n22931, ZN => n5366);
   U23496 : NOR4_X1 port map( A1 => n22940, A2 => n22941, A3 => n22942, A4 => 
                           n22943, ZN => n22930);
   U23497 : NOR4_X1 port map( A1 => n22932, A2 => n22933, A3 => n22934, A4 => 
                           n22935, ZN => n22931);
   U23498 : OAI221_X1 port map( B1 => n20718, B2 => n24996, C1 => n8975, C2 => 
                           n24990, A => n22947, ZN => n22940);
   U23499 : NAND2_X1 port map( A1 => n22912, A2 => n22913, ZN => n5367);
   U23500 : NOR4_X1 port map( A1 => n22922, A2 => n22923, A3 => n22924, A4 => 
                           n22925, ZN => n22912);
   U23501 : NOR4_X1 port map( A1 => n22914, A2 => n22915, A3 => n22916, A4 => 
                           n22917, ZN => n22913);
   U23502 : OAI221_X1 port map( B1 => n20717, B2 => n24996, C1 => n8974, C2 => 
                           n24990, A => n22929, ZN => n22922);
   U23503 : NAND2_X1 port map( A1 => n22894, A2 => n22895, ZN => n5368);
   U23504 : NOR4_X1 port map( A1 => n22904, A2 => n22905, A3 => n22906, A4 => 
                           n22907, ZN => n22894);
   U23505 : NOR4_X1 port map( A1 => n22896, A2 => n22897, A3 => n22898, A4 => 
                           n22899, ZN => n22895);
   U23506 : OAI221_X1 port map( B1 => n20716, B2 => n24996, C1 => n8973, C2 => 
                           n24990, A => n22911, ZN => n22904);
   U23507 : NAND2_X1 port map( A1 => n22876, A2 => n22877, ZN => n5369);
   U23508 : NOR4_X1 port map( A1 => n22886, A2 => n22887, A3 => n22888, A4 => 
                           n22889, ZN => n22876);
   U23509 : NOR4_X1 port map( A1 => n22878, A2 => n22879, A3 => n22880, A4 => 
                           n22881, ZN => n22877);
   U23510 : OAI221_X1 port map( B1 => n20715, B2 => n24996, C1 => n8972, C2 => 
                           n24990, A => n22893, ZN => n22886);
   U23511 : NAND2_X1 port map( A1 => n22858, A2 => n22859, ZN => n5370);
   U23512 : NOR4_X1 port map( A1 => n22868, A2 => n22869, A3 => n22870, A4 => 
                           n22871, ZN => n22858);
   U23513 : NOR4_X1 port map( A1 => n22860, A2 => n22861, A3 => n22862, A4 => 
                           n22863, ZN => n22859);
   U23514 : OAI221_X1 port map( B1 => n20714, B2 => n24996, C1 => n8971, C2 => 
                           n24990, A => n22875, ZN => n22868);
   U23515 : NAND2_X1 port map( A1 => n22723, A2 => n22724, ZN => n5375);
   U23516 : NOR4_X1 port map( A1 => n22744, A2 => n22745, A3 => n22746, A4 => 
                           n22747, ZN => n22723);
   U23517 : NOR4_X1 port map( A1 => n22725, A2 => n22726, A3 => n22727, A4 => 
                           n22728, ZN => n22724);
   U23518 : OAI221_X1 port map( B1 => n20773, B2 => n25190, C1 => n9030, C2 => 
                           n25184, A => n22752, ZN => n22744);
   U23519 : NAND2_X1 port map( A1 => n22705, A2 => n22706, ZN => n5376);
   U23520 : NOR4_X1 port map( A1 => n22715, A2 => n22716, A3 => n22717, A4 => 
                           n22718, ZN => n22705);
   U23521 : NOR4_X1 port map( A1 => n22707, A2 => n22708, A3 => n22709, A4 => 
                           n22710, ZN => n22706);
   U23522 : OAI221_X1 port map( B1 => n20772, B2 => n25190, C1 => n9029, C2 => 
                           n25184, A => n22722, ZN => n22715);
   U23523 : NAND2_X1 port map( A1 => n22687, A2 => n22688, ZN => n5377);
   U23524 : NOR4_X1 port map( A1 => n22697, A2 => n22698, A3 => n22699, A4 => 
                           n22700, ZN => n22687);
   U23525 : NOR4_X1 port map( A1 => n22689, A2 => n22690, A3 => n22691, A4 => 
                           n22692, ZN => n22688);
   U23526 : OAI221_X1 port map( B1 => n20771, B2 => n25190, C1 => n9028, C2 => 
                           n25184, A => n22704, ZN => n22697);
   U23527 : NAND2_X1 port map( A1 => n22669, A2 => n22670, ZN => n5378);
   U23528 : NOR4_X1 port map( A1 => n22679, A2 => n22680, A3 => n22681, A4 => 
                           n22682, ZN => n22669);
   U23529 : NOR4_X1 port map( A1 => n22671, A2 => n22672, A3 => n22673, A4 => 
                           n22674, ZN => n22670);
   U23530 : OAI221_X1 port map( B1 => n20770, B2 => n25190, C1 => n9027, C2 => 
                           n25184, A => n22686, ZN => n22679);
   U23531 : NAND2_X1 port map( A1 => n22651, A2 => n22652, ZN => n5379);
   U23532 : NOR4_X1 port map( A1 => n22661, A2 => n22662, A3 => n22663, A4 => 
                           n22664, ZN => n22651);
   U23533 : NOR4_X1 port map( A1 => n22653, A2 => n22654, A3 => n22655, A4 => 
                           n22656, ZN => n22652);
   U23534 : OAI221_X1 port map( B1 => n20769, B2 => n25190, C1 => n9026, C2 => 
                           n25184, A => n22668, ZN => n22661);
   U23535 : NAND2_X1 port map( A1 => n22633, A2 => n22634, ZN => n5380);
   U23536 : NOR4_X1 port map( A1 => n22643, A2 => n22644, A3 => n22645, A4 => 
                           n22646, ZN => n22633);
   U23537 : NOR4_X1 port map( A1 => n22635, A2 => n22636, A3 => n22637, A4 => 
                           n22638, ZN => n22634);
   U23538 : OAI221_X1 port map( B1 => n20768, B2 => n25190, C1 => n9025, C2 => 
                           n25184, A => n22650, ZN => n22643);
   U23539 : NAND2_X1 port map( A1 => n22615, A2 => n22616, ZN => n5381);
   U23540 : NOR4_X1 port map( A1 => n22625, A2 => n22626, A3 => n22627, A4 => 
                           n22628, ZN => n22615);
   U23541 : NOR4_X1 port map( A1 => n22617, A2 => n22618, A3 => n22619, A4 => 
                           n22620, ZN => n22616);
   U23542 : OAI221_X1 port map( B1 => n20767, B2 => n25190, C1 => n9024, C2 => 
                           n25184, A => n22632, ZN => n22625);
   U23543 : NAND2_X1 port map( A1 => n22597, A2 => n22598, ZN => n5382);
   U23544 : NOR4_X1 port map( A1 => n22607, A2 => n22608, A3 => n22609, A4 => 
                           n22610, ZN => n22597);
   U23545 : NOR4_X1 port map( A1 => n22599, A2 => n22600, A3 => n22601, A4 => 
                           n22602, ZN => n22598);
   U23546 : OAI221_X1 port map( B1 => n20766, B2 => n25190, C1 => n9023, C2 => 
                           n25184, A => n22614, ZN => n22607);
   U23547 : NAND2_X1 port map( A1 => n22579, A2 => n22580, ZN => n5383);
   U23548 : NOR4_X1 port map( A1 => n22589, A2 => n22590, A3 => n22591, A4 => 
                           n22592, ZN => n22579);
   U23549 : NOR4_X1 port map( A1 => n22581, A2 => n22582, A3 => n22583, A4 => 
                           n22584, ZN => n22580);
   U23550 : OAI221_X1 port map( B1 => n20765, B2 => n25190, C1 => n9022, C2 => 
                           n25184, A => n22596, ZN => n22589);
   U23551 : NAND2_X1 port map( A1 => n22561, A2 => n22562, ZN => n5384);
   U23552 : NOR4_X1 port map( A1 => n22571, A2 => n22572, A3 => n22573, A4 => 
                           n22574, ZN => n22561);
   U23553 : NOR4_X1 port map( A1 => n22563, A2 => n22564, A3 => n22565, A4 => 
                           n22566, ZN => n22562);
   U23554 : OAI221_X1 port map( B1 => n20764, B2 => n25190, C1 => n9021, C2 => 
                           n25184, A => n22578, ZN => n22571);
   U23555 : NAND2_X1 port map( A1 => n22543, A2 => n22544, ZN => n5385);
   U23556 : NOR4_X1 port map( A1 => n22553, A2 => n22554, A3 => n22555, A4 => 
                           n22556, ZN => n22543);
   U23557 : NOR4_X1 port map( A1 => n22545, A2 => n22546, A3 => n22547, A4 => 
                           n22548, ZN => n22544);
   U23558 : OAI221_X1 port map( B1 => n20763, B2 => n25190, C1 => n9020, C2 => 
                           n25184, A => n22560, ZN => n22553);
   U23559 : NAND2_X1 port map( A1 => n22525, A2 => n22526, ZN => n5386);
   U23560 : NOR4_X1 port map( A1 => n22535, A2 => n22536, A3 => n22537, A4 => 
                           n22538, ZN => n22525);
   U23561 : NOR4_X1 port map( A1 => n22527, A2 => n22528, A3 => n22529, A4 => 
                           n22530, ZN => n22526);
   U23562 : OAI221_X1 port map( B1 => n20762, B2 => n25190, C1 => n9019, C2 => 
                           n25184, A => n22542, ZN => n22535);
   U23563 : NAND2_X1 port map( A1 => n22507, A2 => n22508, ZN => n5387);
   U23564 : NOR4_X1 port map( A1 => n22517, A2 => n22518, A3 => n22519, A4 => 
                           n22520, ZN => n22507);
   U23565 : NOR4_X1 port map( A1 => n22509, A2 => n22510, A3 => n22511, A4 => 
                           n22512, ZN => n22508);
   U23566 : OAI221_X1 port map( B1 => n20761, B2 => n25191, C1 => n9018, C2 => 
                           n25185, A => n22524, ZN => n22517);
   U23567 : NAND2_X1 port map( A1 => n22489, A2 => n22490, ZN => n5388);
   U23568 : NOR4_X1 port map( A1 => n22499, A2 => n22500, A3 => n22501, A4 => 
                           n22502, ZN => n22489);
   U23569 : NOR4_X1 port map( A1 => n22491, A2 => n22492, A3 => n22493, A4 => 
                           n22494, ZN => n22490);
   U23570 : OAI221_X1 port map( B1 => n20760, B2 => n25191, C1 => n9017, C2 => 
                           n25185, A => n22506, ZN => n22499);
   U23571 : NAND2_X1 port map( A1 => n22471, A2 => n22472, ZN => n5389);
   U23572 : NOR4_X1 port map( A1 => n22481, A2 => n22482, A3 => n22483, A4 => 
                           n22484, ZN => n22471);
   U23573 : NOR4_X1 port map( A1 => n22473, A2 => n22474, A3 => n22475, A4 => 
                           n22476, ZN => n22472);
   U23574 : OAI221_X1 port map( B1 => n20759, B2 => n25191, C1 => n9016, C2 => 
                           n25185, A => n22488, ZN => n22481);
   U23575 : NAND2_X1 port map( A1 => n22453, A2 => n22454, ZN => n5390);
   U23576 : NOR4_X1 port map( A1 => n22463, A2 => n22464, A3 => n22465, A4 => 
                           n22466, ZN => n22453);
   U23577 : NOR4_X1 port map( A1 => n22455, A2 => n22456, A3 => n22457, A4 => 
                           n22458, ZN => n22454);
   U23578 : OAI221_X1 port map( B1 => n20758, B2 => n25191, C1 => n9015, C2 => 
                           n25185, A => n22470, ZN => n22463);
   U23579 : NAND2_X1 port map( A1 => n22435, A2 => n22436, ZN => n5391);
   U23580 : NOR4_X1 port map( A1 => n22445, A2 => n22446, A3 => n22447, A4 => 
                           n22448, ZN => n22435);
   U23581 : NOR4_X1 port map( A1 => n22437, A2 => n22438, A3 => n22439, A4 => 
                           n22440, ZN => n22436);
   U23582 : OAI221_X1 port map( B1 => n20757, B2 => n25191, C1 => n9014, C2 => 
                           n25185, A => n22452, ZN => n22445);
   U23583 : NAND2_X1 port map( A1 => n22417, A2 => n22418, ZN => n5392);
   U23584 : NOR4_X1 port map( A1 => n22427, A2 => n22428, A3 => n22429, A4 => 
                           n22430, ZN => n22417);
   U23585 : NOR4_X1 port map( A1 => n22419, A2 => n22420, A3 => n22421, A4 => 
                           n22422, ZN => n22418);
   U23586 : OAI221_X1 port map( B1 => n20756, B2 => n25191, C1 => n9013, C2 => 
                           n25185, A => n22434, ZN => n22427);
   U23587 : NAND2_X1 port map( A1 => n22399, A2 => n22400, ZN => n5393);
   U23588 : NOR4_X1 port map( A1 => n22409, A2 => n22410, A3 => n22411, A4 => 
                           n22412, ZN => n22399);
   U23589 : NOR4_X1 port map( A1 => n22401, A2 => n22402, A3 => n22403, A4 => 
                           n22404, ZN => n22400);
   U23590 : OAI221_X1 port map( B1 => n20755, B2 => n25191, C1 => n9012, C2 => 
                           n25185, A => n22416, ZN => n22409);
   U23591 : NAND2_X1 port map( A1 => n22381, A2 => n22382, ZN => n5394);
   U23592 : NOR4_X1 port map( A1 => n22391, A2 => n22392, A3 => n22393, A4 => 
                           n22394, ZN => n22381);
   U23593 : NOR4_X1 port map( A1 => n22383, A2 => n22384, A3 => n22385, A4 => 
                           n22386, ZN => n22382);
   U23594 : OAI221_X1 port map( B1 => n20754, B2 => n25191, C1 => n9011, C2 => 
                           n25185, A => n22398, ZN => n22391);
   U23595 : NAND2_X1 port map( A1 => n22363, A2 => n22364, ZN => n5395);
   U23596 : NOR4_X1 port map( A1 => n22373, A2 => n22374, A3 => n22375, A4 => 
                           n22376, ZN => n22363);
   U23597 : NOR4_X1 port map( A1 => n22365, A2 => n22366, A3 => n22367, A4 => 
                           n22368, ZN => n22364);
   U23598 : OAI221_X1 port map( B1 => n20753, B2 => n25191, C1 => n9010, C2 => 
                           n25185, A => n22380, ZN => n22373);
   U23599 : NAND2_X1 port map( A1 => n22345, A2 => n22346, ZN => n5396);
   U23600 : NOR4_X1 port map( A1 => n22355, A2 => n22356, A3 => n22357, A4 => 
                           n22358, ZN => n22345);
   U23601 : NOR4_X1 port map( A1 => n22347, A2 => n22348, A3 => n22349, A4 => 
                           n22350, ZN => n22346);
   U23602 : OAI221_X1 port map( B1 => n20752, B2 => n25191, C1 => n9009, C2 => 
                           n25185, A => n22362, ZN => n22355);
   U23603 : NAND2_X1 port map( A1 => n22327, A2 => n22328, ZN => n5397);
   U23604 : NOR4_X1 port map( A1 => n22337, A2 => n22338, A3 => n22339, A4 => 
                           n22340, ZN => n22327);
   U23605 : NOR4_X1 port map( A1 => n22329, A2 => n22330, A3 => n22331, A4 => 
                           n22332, ZN => n22328);
   U23606 : OAI221_X1 port map( B1 => n20751, B2 => n25191, C1 => n9008, C2 => 
                           n25185, A => n22344, ZN => n22337);
   U23607 : NAND2_X1 port map( A1 => n22309, A2 => n22310, ZN => n5398);
   U23608 : NOR4_X1 port map( A1 => n22319, A2 => n22320, A3 => n22321, A4 => 
                           n22322, ZN => n22309);
   U23609 : NOR4_X1 port map( A1 => n22311, A2 => n22312, A3 => n22313, A4 => 
                           n22314, ZN => n22310);
   U23610 : OAI221_X1 port map( B1 => n20750, B2 => n25191, C1 => n9007, C2 => 
                           n25185, A => n22326, ZN => n22319);
   U23611 : NAND2_X1 port map( A1 => n22291, A2 => n22292, ZN => n5399);
   U23612 : NOR4_X1 port map( A1 => n22301, A2 => n22302, A3 => n22303, A4 => 
                           n22304, ZN => n22291);
   U23613 : NOR4_X1 port map( A1 => n22293, A2 => n22294, A3 => n22295, A4 => 
                           n22296, ZN => n22292);
   U23614 : OAI221_X1 port map( B1 => n20749, B2 => n25192, C1 => n9006, C2 => 
                           n25186, A => n22308, ZN => n22301);
   U23615 : NAND2_X1 port map( A1 => n22273, A2 => n22274, ZN => n5400);
   U23616 : NOR4_X1 port map( A1 => n22283, A2 => n22284, A3 => n22285, A4 => 
                           n22286, ZN => n22273);
   U23617 : NOR4_X1 port map( A1 => n22275, A2 => n22276, A3 => n22277, A4 => 
                           n22278, ZN => n22274);
   U23618 : OAI221_X1 port map( B1 => n20748, B2 => n25192, C1 => n9005, C2 => 
                           n25186, A => n22290, ZN => n22283);
   U23619 : NAND2_X1 port map( A1 => n22255, A2 => n22256, ZN => n5401);
   U23620 : NOR4_X1 port map( A1 => n22265, A2 => n22266, A3 => n22267, A4 => 
                           n22268, ZN => n22255);
   U23621 : NOR4_X1 port map( A1 => n22257, A2 => n22258, A3 => n22259, A4 => 
                           n22260, ZN => n22256);
   U23622 : OAI221_X1 port map( B1 => n20747, B2 => n25192, C1 => n9004, C2 => 
                           n25186, A => n22272, ZN => n22265);
   U23623 : NAND2_X1 port map( A1 => n22237, A2 => n22238, ZN => n5402);
   U23624 : NOR4_X1 port map( A1 => n22247, A2 => n22248, A3 => n22249, A4 => 
                           n22250, ZN => n22237);
   U23625 : NOR4_X1 port map( A1 => n22239, A2 => n22240, A3 => n22241, A4 => 
                           n22242, ZN => n22238);
   U23626 : OAI221_X1 port map( B1 => n20746, B2 => n25192, C1 => n9003, C2 => 
                           n25186, A => n22254, ZN => n22247);
   U23627 : NAND2_X1 port map( A1 => n22219, A2 => n22220, ZN => n5403);
   U23628 : NOR4_X1 port map( A1 => n22229, A2 => n22230, A3 => n22231, A4 => 
                           n22232, ZN => n22219);
   U23629 : NOR4_X1 port map( A1 => n22221, A2 => n22222, A3 => n22223, A4 => 
                           n22224, ZN => n22220);
   U23630 : OAI221_X1 port map( B1 => n20745, B2 => n25192, C1 => n9002, C2 => 
                           n25186, A => n22236, ZN => n22229);
   U23631 : NAND2_X1 port map( A1 => n22201, A2 => n22202, ZN => n5404);
   U23632 : NOR4_X1 port map( A1 => n22211, A2 => n22212, A3 => n22213, A4 => 
                           n22214, ZN => n22201);
   U23633 : NOR4_X1 port map( A1 => n22203, A2 => n22204, A3 => n22205, A4 => 
                           n22206, ZN => n22202);
   U23634 : OAI221_X1 port map( B1 => n20744, B2 => n25192, C1 => n9001, C2 => 
                           n25186, A => n22218, ZN => n22211);
   U23635 : NAND2_X1 port map( A1 => n22183, A2 => n22184, ZN => n5405);
   U23636 : NOR4_X1 port map( A1 => n22193, A2 => n22194, A3 => n22195, A4 => 
                           n22196, ZN => n22183);
   U23637 : NOR4_X1 port map( A1 => n22185, A2 => n22186, A3 => n22187, A4 => 
                           n22188, ZN => n22184);
   U23638 : OAI221_X1 port map( B1 => n20743, B2 => n25192, C1 => n9000, C2 => 
                           n25186, A => n22200, ZN => n22193);
   U23639 : NAND2_X1 port map( A1 => n22165, A2 => n22166, ZN => n5406);
   U23640 : NOR4_X1 port map( A1 => n22175, A2 => n22176, A3 => n22177, A4 => 
                           n22178, ZN => n22165);
   U23641 : NOR4_X1 port map( A1 => n22167, A2 => n22168, A3 => n22169, A4 => 
                           n22170, ZN => n22166);
   U23642 : OAI221_X1 port map( B1 => n20742, B2 => n25192, C1 => n8999, C2 => 
                           n25186, A => n22182, ZN => n22175);
   U23643 : NAND2_X1 port map( A1 => n22147, A2 => n22148, ZN => n5407);
   U23644 : NOR4_X1 port map( A1 => n22157, A2 => n22158, A3 => n22159, A4 => 
                           n22160, ZN => n22147);
   U23645 : NOR4_X1 port map( A1 => n22149, A2 => n22150, A3 => n22151, A4 => 
                           n22152, ZN => n22148);
   U23646 : OAI221_X1 port map( B1 => n20741, B2 => n25192, C1 => n8998, C2 => 
                           n25186, A => n22164, ZN => n22157);
   U23647 : NAND2_X1 port map( A1 => n22129, A2 => n22130, ZN => n5408);
   U23648 : NOR4_X1 port map( A1 => n22139, A2 => n22140, A3 => n22141, A4 => 
                           n22142, ZN => n22129);
   U23649 : NOR4_X1 port map( A1 => n22131, A2 => n22132, A3 => n22133, A4 => 
                           n22134, ZN => n22130);
   U23650 : OAI221_X1 port map( B1 => n20740, B2 => n25192, C1 => n8997, C2 => 
                           n25186, A => n22146, ZN => n22139);
   U23651 : NAND2_X1 port map( A1 => n22111, A2 => n22112, ZN => n5409);
   U23652 : NOR4_X1 port map( A1 => n22121, A2 => n22122, A3 => n22123, A4 => 
                           n22124, ZN => n22111);
   U23653 : NOR4_X1 port map( A1 => n22113, A2 => n22114, A3 => n22115, A4 => 
                           n22116, ZN => n22112);
   U23654 : OAI221_X1 port map( B1 => n20739, B2 => n25192, C1 => n8996, C2 => 
                           n25186, A => n22128, ZN => n22121);
   U23655 : NAND2_X1 port map( A1 => n22093, A2 => n22094, ZN => n5410);
   U23656 : NOR4_X1 port map( A1 => n22103, A2 => n22104, A3 => n22105, A4 => 
                           n22106, ZN => n22093);
   U23657 : NOR4_X1 port map( A1 => n22095, A2 => n22096, A3 => n22097, A4 => 
                           n22098, ZN => n22094);
   U23658 : OAI221_X1 port map( B1 => n20738, B2 => n25192, C1 => n8995, C2 => 
                           n25186, A => n22110, ZN => n22103);
   U23659 : NAND2_X1 port map( A1 => n22075, A2 => n22076, ZN => n5411);
   U23660 : NOR4_X1 port map( A1 => n22085, A2 => n22086, A3 => n22087, A4 => 
                           n22088, ZN => n22075);
   U23661 : NOR4_X1 port map( A1 => n22077, A2 => n22078, A3 => n22079, A4 => 
                           n22080, ZN => n22076);
   U23662 : OAI221_X1 port map( B1 => n20737, B2 => n25193, C1 => n8994, C2 => 
                           n25187, A => n22092, ZN => n22085);
   U23663 : NAND2_X1 port map( A1 => n22057, A2 => n22058, ZN => n5412);
   U23664 : NOR4_X1 port map( A1 => n22067, A2 => n22068, A3 => n22069, A4 => 
                           n22070, ZN => n22057);
   U23665 : NOR4_X1 port map( A1 => n22059, A2 => n22060, A3 => n22061, A4 => 
                           n22062, ZN => n22058);
   U23666 : OAI221_X1 port map( B1 => n20736, B2 => n25193, C1 => n8993, C2 => 
                           n25187, A => n22074, ZN => n22067);
   U23667 : NAND2_X1 port map( A1 => n22039, A2 => n22040, ZN => n5413);
   U23668 : NOR4_X1 port map( A1 => n22049, A2 => n22050, A3 => n22051, A4 => 
                           n22052, ZN => n22039);
   U23669 : NOR4_X1 port map( A1 => n22041, A2 => n22042, A3 => n22043, A4 => 
                           n22044, ZN => n22040);
   U23670 : OAI221_X1 port map( B1 => n20735, B2 => n25193, C1 => n8992, C2 => 
                           n25187, A => n22056, ZN => n22049);
   U23671 : NAND2_X1 port map( A1 => n22021, A2 => n22022, ZN => n5414);
   U23672 : NOR4_X1 port map( A1 => n22031, A2 => n22032, A3 => n22033, A4 => 
                           n22034, ZN => n22021);
   U23673 : NOR4_X1 port map( A1 => n22023, A2 => n22024, A3 => n22025, A4 => 
                           n22026, ZN => n22022);
   U23674 : OAI221_X1 port map( B1 => n20734, B2 => n25193, C1 => n8991, C2 => 
                           n25187, A => n22038, ZN => n22031);
   U23675 : NAND2_X1 port map( A1 => n22003, A2 => n22004, ZN => n5415);
   U23676 : NOR4_X1 port map( A1 => n22013, A2 => n22014, A3 => n22015, A4 => 
                           n22016, ZN => n22003);
   U23677 : NOR4_X1 port map( A1 => n22005, A2 => n22006, A3 => n22007, A4 => 
                           n22008, ZN => n22004);
   U23678 : OAI221_X1 port map( B1 => n20733, B2 => n25193, C1 => n8990, C2 => 
                           n25187, A => n22020, ZN => n22013);
   U23679 : NAND2_X1 port map( A1 => n21985, A2 => n21986, ZN => n5416);
   U23680 : NOR4_X1 port map( A1 => n21995, A2 => n21996, A3 => n21997, A4 => 
                           n21998, ZN => n21985);
   U23681 : NOR4_X1 port map( A1 => n21987, A2 => n21988, A3 => n21989, A4 => 
                           n21990, ZN => n21986);
   U23682 : OAI221_X1 port map( B1 => n20732, B2 => n25193, C1 => n8989, C2 => 
                           n25187, A => n22002, ZN => n21995);
   U23683 : NAND2_X1 port map( A1 => n21967, A2 => n21968, ZN => n5417);
   U23684 : NOR4_X1 port map( A1 => n21977, A2 => n21978, A3 => n21979, A4 => 
                           n21980, ZN => n21967);
   U23685 : NOR4_X1 port map( A1 => n21969, A2 => n21970, A3 => n21971, A4 => 
                           n21972, ZN => n21968);
   U23686 : OAI221_X1 port map( B1 => n20731, B2 => n25193, C1 => n8988, C2 => 
                           n25187, A => n21984, ZN => n21977);
   U23687 : NAND2_X1 port map( A1 => n21949, A2 => n21950, ZN => n5418);
   U23688 : NOR4_X1 port map( A1 => n21959, A2 => n21960, A3 => n21961, A4 => 
                           n21962, ZN => n21949);
   U23689 : NOR4_X1 port map( A1 => n21951, A2 => n21952, A3 => n21953, A4 => 
                           n21954, ZN => n21950);
   U23690 : OAI221_X1 port map( B1 => n20730, B2 => n25193, C1 => n8987, C2 => 
                           n25187, A => n21966, ZN => n21959);
   U23691 : NAND2_X1 port map( A1 => n21931, A2 => n21932, ZN => n5419);
   U23692 : NOR4_X1 port map( A1 => n21941, A2 => n21942, A3 => n21943, A4 => 
                           n21944, ZN => n21931);
   U23693 : NOR4_X1 port map( A1 => n21933, A2 => n21934, A3 => n21935, A4 => 
                           n21936, ZN => n21932);
   U23694 : OAI221_X1 port map( B1 => n20729, B2 => n25193, C1 => n8986, C2 => 
                           n25187, A => n21948, ZN => n21941);
   U23695 : NAND2_X1 port map( A1 => n21913, A2 => n21914, ZN => n5420);
   U23696 : NOR4_X1 port map( A1 => n21923, A2 => n21924, A3 => n21925, A4 => 
                           n21926, ZN => n21913);
   U23697 : NOR4_X1 port map( A1 => n21915, A2 => n21916, A3 => n21917, A4 => 
                           n21918, ZN => n21914);
   U23698 : OAI221_X1 port map( B1 => n20728, B2 => n25193, C1 => n8985, C2 => 
                           n25187, A => n21930, ZN => n21923);
   U23699 : NAND2_X1 port map( A1 => n21895, A2 => n21896, ZN => n5421);
   U23700 : NOR4_X1 port map( A1 => n21905, A2 => n21906, A3 => n21907, A4 => 
                           n21908, ZN => n21895);
   U23701 : NOR4_X1 port map( A1 => n21897, A2 => n21898, A3 => n21899, A4 => 
                           n21900, ZN => n21896);
   U23702 : OAI221_X1 port map( B1 => n20727, B2 => n25193, C1 => n8984, C2 => 
                           n25187, A => n21912, ZN => n21905);
   U23703 : NAND2_X1 port map( A1 => n21877, A2 => n21878, ZN => n5422);
   U23704 : NOR4_X1 port map( A1 => n21887, A2 => n21888, A3 => n21889, A4 => 
                           n21890, ZN => n21877);
   U23705 : NOR4_X1 port map( A1 => n21879, A2 => n21880, A3 => n21881, A4 => 
                           n21882, ZN => n21878);
   U23706 : OAI221_X1 port map( B1 => n20726, B2 => n25193, C1 => n8983, C2 => 
                           n25187, A => n21894, ZN => n21887);
   U23707 : NAND2_X1 port map( A1 => n21859, A2 => n21860, ZN => n5423);
   U23708 : NOR4_X1 port map( A1 => n21869, A2 => n21870, A3 => n21871, A4 => 
                           n21872, ZN => n21859);
   U23709 : NOR4_X1 port map( A1 => n21861, A2 => n21862, A3 => n21863, A4 => 
                           n21864, ZN => n21860);
   U23710 : OAI221_X1 port map( B1 => n20725, B2 => n25194, C1 => n8982, C2 => 
                           n25188, A => n21876, ZN => n21869);
   U23711 : NAND2_X1 port map( A1 => n21841, A2 => n21842, ZN => n5424);
   U23712 : NOR4_X1 port map( A1 => n21851, A2 => n21852, A3 => n21853, A4 => 
                           n21854, ZN => n21841);
   U23713 : NOR4_X1 port map( A1 => n21843, A2 => n21844, A3 => n21845, A4 => 
                           n21846, ZN => n21842);
   U23714 : OAI221_X1 port map( B1 => n20724, B2 => n25194, C1 => n8981, C2 => 
                           n25188, A => n21858, ZN => n21851);
   U23715 : NAND2_X1 port map( A1 => n21823, A2 => n21824, ZN => n5425);
   U23716 : NOR4_X1 port map( A1 => n21833, A2 => n21834, A3 => n21835, A4 => 
                           n21836, ZN => n21823);
   U23717 : NOR4_X1 port map( A1 => n21825, A2 => n21826, A3 => n21827, A4 => 
                           n21828, ZN => n21824);
   U23718 : OAI221_X1 port map( B1 => n20723, B2 => n25194, C1 => n8980, C2 => 
                           n25188, A => n21840, ZN => n21833);
   U23719 : NAND2_X1 port map( A1 => n21805, A2 => n21806, ZN => n5426);
   U23720 : NOR4_X1 port map( A1 => n21815, A2 => n21816, A3 => n21817, A4 => 
                           n21818, ZN => n21805);
   U23721 : NOR4_X1 port map( A1 => n21807, A2 => n21808, A3 => n21809, A4 => 
                           n21810, ZN => n21806);
   U23722 : OAI221_X1 port map( B1 => n20722, B2 => n25194, C1 => n8979, C2 => 
                           n25188, A => n21822, ZN => n21815);
   U23723 : NAND2_X1 port map( A1 => n21787, A2 => n21788, ZN => n5427);
   U23724 : NOR4_X1 port map( A1 => n21797, A2 => n21798, A3 => n21799, A4 => 
                           n21800, ZN => n21787);
   U23725 : NOR4_X1 port map( A1 => n21789, A2 => n21790, A3 => n21791, A4 => 
                           n21792, ZN => n21788);
   U23726 : OAI221_X1 port map( B1 => n20721, B2 => n25194, C1 => n8978, C2 => 
                           n25188, A => n21804, ZN => n21797);
   U23727 : NAND2_X1 port map( A1 => n21769, A2 => n21770, ZN => n5428);
   U23728 : NOR4_X1 port map( A1 => n21779, A2 => n21780, A3 => n21781, A4 => 
                           n21782, ZN => n21769);
   U23729 : NOR4_X1 port map( A1 => n21771, A2 => n21772, A3 => n21773, A4 => 
                           n21774, ZN => n21770);
   U23730 : OAI221_X1 port map( B1 => n20720, B2 => n25194, C1 => n8977, C2 => 
                           n25188, A => n21786, ZN => n21779);
   U23731 : NAND2_X1 port map( A1 => n21751, A2 => n21752, ZN => n5429);
   U23732 : NOR4_X1 port map( A1 => n21761, A2 => n21762, A3 => n21763, A4 => 
                           n21764, ZN => n21751);
   U23733 : NOR4_X1 port map( A1 => n21753, A2 => n21754, A3 => n21755, A4 => 
                           n21756, ZN => n21752);
   U23734 : OAI221_X1 port map( B1 => n20719, B2 => n25194, C1 => n8976, C2 => 
                           n25188, A => n21768, ZN => n21761);
   U23735 : NAND2_X1 port map( A1 => n21733, A2 => n21734, ZN => n5430);
   U23736 : NOR4_X1 port map( A1 => n21743, A2 => n21744, A3 => n21745, A4 => 
                           n21746, ZN => n21733);
   U23737 : NOR4_X1 port map( A1 => n21735, A2 => n21736, A3 => n21737, A4 => 
                           n21738, ZN => n21734);
   U23738 : OAI221_X1 port map( B1 => n20718, B2 => n25194, C1 => n8975, C2 => 
                           n25188, A => n21750, ZN => n21743);
   U23739 : NAND2_X1 port map( A1 => n21715, A2 => n21716, ZN => n5431);
   U23740 : NOR4_X1 port map( A1 => n21725, A2 => n21726, A3 => n21727, A4 => 
                           n21728, ZN => n21715);
   U23741 : NOR4_X1 port map( A1 => n21717, A2 => n21718, A3 => n21719, A4 => 
                           n21720, ZN => n21716);
   U23742 : OAI221_X1 port map( B1 => n20717, B2 => n25194, C1 => n8974, C2 => 
                           n25188, A => n21732, ZN => n21725);
   U23743 : NAND2_X1 port map( A1 => n21697, A2 => n21698, ZN => n5432);
   U23744 : NOR4_X1 port map( A1 => n21707, A2 => n21708, A3 => n21709, A4 => 
                           n21710, ZN => n21697);
   U23745 : NOR4_X1 port map( A1 => n21699, A2 => n21700, A3 => n21701, A4 => 
                           n21702, ZN => n21698);
   U23746 : OAI221_X1 port map( B1 => n20716, B2 => n25194, C1 => n8973, C2 => 
                           n25188, A => n21714, ZN => n21707);
   U23747 : NAND2_X1 port map( A1 => n21679, A2 => n21680, ZN => n5433);
   U23748 : NOR4_X1 port map( A1 => n21689, A2 => n21690, A3 => n21691, A4 => 
                           n21692, ZN => n21679);
   U23749 : NOR4_X1 port map( A1 => n21681, A2 => n21682, A3 => n21683, A4 => 
                           n21684, ZN => n21680);
   U23750 : OAI221_X1 port map( B1 => n20715, B2 => n25194, C1 => n8972, C2 => 
                           n25188, A => n21696, ZN => n21689);
   U23751 : NAND2_X1 port map( A1 => n21661, A2 => n21662, ZN => n5434);
   U23752 : NOR4_X1 port map( A1 => n21671, A2 => n21672, A3 => n21673, A4 => 
                           n21674, ZN => n21661);
   U23753 : NOR4_X1 port map( A1 => n21663, A2 => n21664, A3 => n21665, A4 => 
                           n21666, ZN => n21662);
   U23754 : OAI221_X1 port map( B1 => n20714, B2 => n25194, C1 => n8971, C2 => 
                           n25188, A => n21678, ZN => n21671);
   U23755 : OAI22_X1 port map( A1 => n25597, A2 => n21477, B1 => n25782, B2 => 
                           n25589, ZN => n6527);
   U23756 : OAI22_X1 port map( A1 => n25597, A2 => n21476, B1 => n25785, B2 => 
                           n25589, ZN => n6528);
   U23757 : OAI22_X1 port map( A1 => n25597, A2 => n21475, B1 => n25788, B2 => 
                           n25589, ZN => n6529);
   U23758 : OAI22_X1 port map( A1 => n25597, A2 => n21474, B1 => n25791, B2 => 
                           n25589, ZN => n6530);
   U23759 : OAI22_X1 port map( A1 => n25597, A2 => n21473, B1 => n25794, B2 => 
                           n25589, ZN => n6531);
   U23760 : OAI22_X1 port map( A1 => n25597, A2 => n21472, B1 => n25797, B2 => 
                           n25589, ZN => n6532);
   U23761 : OAI22_X1 port map( A1 => n25597, A2 => n21471, B1 => n25800, B2 => 
                           n25589, ZN => n6533);
   U23762 : OAI22_X1 port map( A1 => n25597, A2 => n21470, B1 => n25803, B2 => 
                           n25589, ZN => n6534);
   U23763 : OAI22_X1 port map( A1 => n25597, A2 => n21469, B1 => n25806, B2 => 
                           n25589, ZN => n6535);
   U23764 : OAI22_X1 port map( A1 => n25597, A2 => n21468, B1 => n25809, B2 => 
                           n25589, ZN => n6536);
   U23765 : OAI22_X1 port map( A1 => n25597, A2 => n21467, B1 => n25812, B2 => 
                           n25589, ZN => n6537);
   U23766 : OAI22_X1 port map( A1 => n25597, A2 => n21466, B1 => n25815, B2 => 
                           n25589, ZN => n6538);
   U23767 : OAI22_X1 port map( A1 => n25598, A2 => n21465, B1 => n25818, B2 => 
                           n25590, ZN => n6539);
   U23768 : OAI22_X1 port map( A1 => n25598, A2 => n21464, B1 => n25821, B2 => 
                           n25590, ZN => n6540);
   U23769 : OAI22_X1 port map( A1 => n25598, A2 => n21463, B1 => n25824, B2 => 
                           n25590, ZN => n6541);
   U23770 : OAI22_X1 port map( A1 => n25598, A2 => n21462, B1 => n25827, B2 => 
                           n25590, ZN => n6542);
   U23771 : OAI22_X1 port map( A1 => n25598, A2 => n21461, B1 => n25830, B2 => 
                           n25590, ZN => n6543);
   U23772 : OAI22_X1 port map( A1 => n25598, A2 => n21460, B1 => n25833, B2 => 
                           n25590, ZN => n6544);
   U23773 : OAI22_X1 port map( A1 => n25598, A2 => n21459, B1 => n25836, B2 => 
                           n25590, ZN => n6545);
   U23774 : OAI22_X1 port map( A1 => n25598, A2 => n21458, B1 => n25839, B2 => 
                           n25590, ZN => n6546);
   U23775 : OAI22_X1 port map( A1 => n25598, A2 => n21457, B1 => n25842, B2 => 
                           n25590, ZN => n6547);
   U23776 : OAI22_X1 port map( A1 => n25598, A2 => n21456, B1 => n25845, B2 => 
                           n25590, ZN => n6548);
   U23777 : OAI22_X1 port map( A1 => n25598, A2 => n21455, B1 => n25848, B2 => 
                           n25590, ZN => n6549);
   U23778 : OAI22_X1 port map( A1 => n25598, A2 => n21454, B1 => n25851, B2 => 
                           n25590, ZN => n6550);
   U23779 : OAI22_X1 port map( A1 => n25598, A2 => n21453, B1 => n25854, B2 => 
                           n25591, ZN => n6551);
   U23780 : OAI22_X1 port map( A1 => n25599, A2 => n21452, B1 => n25857, B2 => 
                           n25591, ZN => n6552);
   U23781 : OAI22_X1 port map( A1 => n25599, A2 => n21451, B1 => n25860, B2 => 
                           n25591, ZN => n6553);
   U23782 : OAI22_X1 port map( A1 => n25599, A2 => n21450, B1 => n25863, B2 => 
                           n25591, ZN => n6554);
   U23783 : OAI22_X1 port map( A1 => n25599, A2 => n21449, B1 => n25866, B2 => 
                           n25591, ZN => n6555);
   U23784 : OAI22_X1 port map( A1 => n25599, A2 => n21448, B1 => n25869, B2 => 
                           n25591, ZN => n6556);
   U23785 : OAI22_X1 port map( A1 => n25599, A2 => n21447, B1 => n25872, B2 => 
                           n25591, ZN => n6557);
   U23786 : OAI22_X1 port map( A1 => n25599, A2 => n21446, B1 => n25875, B2 => 
                           n25591, ZN => n6558);
   U23787 : OAI22_X1 port map( A1 => n25599, A2 => n21445, B1 => n25878, B2 => 
                           n25591, ZN => n6559);
   U23788 : OAI22_X1 port map( A1 => n25599, A2 => n21444, B1 => n25881, B2 => 
                           n25591, ZN => n6560);
   U23789 : OAI22_X1 port map( A1 => n25599, A2 => n21443, B1 => n25884, B2 => 
                           n25591, ZN => n6561);
   U23790 : OAI22_X1 port map( A1 => n25599, A2 => n21442, B1 => n25887, B2 => 
                           n25591, ZN => n6562);
   U23791 : OAI22_X1 port map( A1 => n25599, A2 => n21441, B1 => n25890, B2 => 
                           n25592, ZN => n6563);
   U23792 : OAI22_X1 port map( A1 => n25599, A2 => n21440, B1 => n25893, B2 => 
                           n25592, ZN => n6564);
   U23793 : OAI22_X1 port map( A1 => n25600, A2 => n21439, B1 => n25896, B2 => 
                           n25592, ZN => n6565);
   U23794 : OAI22_X1 port map( A1 => n25600, A2 => n21438, B1 => n25899, B2 => 
                           n25592, ZN => n6566);
   U23795 : OAI22_X1 port map( A1 => n25600, A2 => n21437, B1 => n25902, B2 => 
                           n25592, ZN => n6567);
   U23796 : OAI22_X1 port map( A1 => n25600, A2 => n21436, B1 => n25905, B2 => 
                           n25592, ZN => n6568);
   U23797 : OAI22_X1 port map( A1 => n25600, A2 => n21435, B1 => n25908, B2 => 
                           n25592, ZN => n6569);
   U23798 : OAI22_X1 port map( A1 => n25600, A2 => n21434, B1 => n25911, B2 => 
                           n25592, ZN => n6570);
   U23799 : OAI22_X1 port map( A1 => n25600, A2 => n21433, B1 => n25914, B2 => 
                           n25592, ZN => n6571);
   U23800 : OAI22_X1 port map( A1 => n25600, A2 => n21432, B1 => n25917, B2 => 
                           n25592, ZN => n6572);
   U23801 : OAI22_X1 port map( A1 => n25600, A2 => n21431, B1 => n25920, B2 => 
                           n25592, ZN => n6573);
   U23802 : OAI22_X1 port map( A1 => n25600, A2 => n21430, B1 => n25923, B2 => 
                           n25592, ZN => n6574);
   U23803 : OAI22_X1 port map( A1 => n25600, A2 => n21429, B1 => n25926, B2 => 
                           n25593, ZN => n6575);
   U23804 : OAI22_X1 port map( A1 => n25600, A2 => n21428, B1 => n25929, B2 => 
                           n25593, ZN => n6576);
   U23805 : OAI22_X1 port map( A1 => n25600, A2 => n21427, B1 => n25932, B2 => 
                           n25593, ZN => n6577);
   U23806 : OAI22_X1 port map( A1 => n25601, A2 => n21426, B1 => n25935, B2 => 
                           n25593, ZN => n6578);
   U23807 : OAI22_X1 port map( A1 => n25601, A2 => n21425, B1 => n25938, B2 => 
                           n25593, ZN => n6579);
   U23808 : OAI22_X1 port map( A1 => n25601, A2 => n21424, B1 => n25941, B2 => 
                           n25593, ZN => n6580);
   U23809 : OAI22_X1 port map( A1 => n25601, A2 => n21423, B1 => n25944, B2 => 
                           n25593, ZN => n6581);
   U23810 : OAI22_X1 port map( A1 => n25601, A2 => n21422, B1 => n25947, B2 => 
                           n25593, ZN => n6582);
   U23811 : OAI22_X1 port map( A1 => n25601, A2 => n21421, B1 => n25950, B2 => 
                           n25593, ZN => n6583);
   U23812 : OAI22_X1 port map( A1 => n25601, A2 => n21420, B1 => n25953, B2 => 
                           n25593, ZN => n6584);
   U23813 : OAI22_X1 port map( A1 => n25601, A2 => n21419, B1 => n25956, B2 => 
                           n25593, ZN => n6585);
   U23814 : OAI22_X1 port map( A1 => n25601, A2 => n21418, B1 => n25959, B2 => 
                           n25593, ZN => n6586);
   U23815 : OAI22_X1 port map( A1 => n25572, A2 => n20965, B1 => n25782, B2 => 
                           n25564, ZN => n6399);
   U23816 : OAI22_X1 port map( A1 => n25572, A2 => n20964, B1 => n25785, B2 => 
                           n25564, ZN => n6400);
   U23817 : OAI22_X1 port map( A1 => n25572, A2 => n20963, B1 => n25788, B2 => 
                           n25564, ZN => n6401);
   U23818 : OAI22_X1 port map( A1 => n25572, A2 => n20962, B1 => n25791, B2 => 
                           n25564, ZN => n6402);
   U23819 : OAI22_X1 port map( A1 => n25572, A2 => n20961, B1 => n25794, B2 => 
                           n25564, ZN => n6403);
   U23820 : OAI22_X1 port map( A1 => n25572, A2 => n20960, B1 => n25797, B2 => 
                           n25564, ZN => n6404);
   U23821 : OAI22_X1 port map( A1 => n25572, A2 => n20959, B1 => n25800, B2 => 
                           n25564, ZN => n6405);
   U23822 : OAI22_X1 port map( A1 => n25572, A2 => n20958, B1 => n25803, B2 => 
                           n25564, ZN => n6406);
   U23823 : OAI22_X1 port map( A1 => n25572, A2 => n20957, B1 => n25806, B2 => 
                           n25564, ZN => n6407);
   U23824 : OAI22_X1 port map( A1 => n25572, A2 => n20956, B1 => n25809, B2 => 
                           n25564, ZN => n6408);
   U23825 : OAI22_X1 port map( A1 => n25572, A2 => n20955, B1 => n25812, B2 => 
                           n25564, ZN => n6409);
   U23826 : OAI22_X1 port map( A1 => n25572, A2 => n20954, B1 => n25815, B2 => 
                           n25564, ZN => n6410);
   U23827 : OAI22_X1 port map( A1 => n25573, A2 => n20953, B1 => n25818, B2 => 
                           n25565, ZN => n6411);
   U23828 : OAI22_X1 port map( A1 => n25573, A2 => n20952, B1 => n25821, B2 => 
                           n25565, ZN => n6412);
   U23829 : OAI22_X1 port map( A1 => n25573, A2 => n20951, B1 => n25824, B2 => 
                           n25565, ZN => n6413);
   U23830 : OAI22_X1 port map( A1 => n25573, A2 => n20950, B1 => n25827, B2 => 
                           n25565, ZN => n6414);
   U23831 : OAI22_X1 port map( A1 => n25573, A2 => n20949, B1 => n25830, B2 => 
                           n25565, ZN => n6415);
   U23832 : OAI22_X1 port map( A1 => n25573, A2 => n20948, B1 => n25833, B2 => 
                           n25565, ZN => n6416);
   U23833 : OAI22_X1 port map( A1 => n25573, A2 => n20947, B1 => n25836, B2 => 
                           n25565, ZN => n6417);
   U23834 : OAI22_X1 port map( A1 => n25573, A2 => n20946, B1 => n25839, B2 => 
                           n25565, ZN => n6418);
   U23835 : OAI22_X1 port map( A1 => n25573, A2 => n20945, B1 => n25842, B2 => 
                           n25565, ZN => n6419);
   U23836 : OAI22_X1 port map( A1 => n25573, A2 => n20944, B1 => n25845, B2 => 
                           n25565, ZN => n6420);
   U23837 : OAI22_X1 port map( A1 => n25573, A2 => n20943, B1 => n25848, B2 => 
                           n25565, ZN => n6421);
   U23838 : OAI22_X1 port map( A1 => n25573, A2 => n20942, B1 => n25851, B2 => 
                           n25565, ZN => n6422);
   U23839 : OAI22_X1 port map( A1 => n25573, A2 => n20941, B1 => n25854, B2 => 
                           n25566, ZN => n6423);
   U23840 : OAI22_X1 port map( A1 => n25574, A2 => n20940, B1 => n25857, B2 => 
                           n25566, ZN => n6424);
   U23841 : OAI22_X1 port map( A1 => n25574, A2 => n20939, B1 => n25860, B2 => 
                           n25566, ZN => n6425);
   U23842 : OAI22_X1 port map( A1 => n25574, A2 => n20938, B1 => n25863, B2 => 
                           n25566, ZN => n6426);
   U23843 : OAI22_X1 port map( A1 => n25574, A2 => n20937, B1 => n25866, B2 => 
                           n25566, ZN => n6427);
   U23844 : OAI22_X1 port map( A1 => n25574, A2 => n20936, B1 => n25869, B2 => 
                           n25566, ZN => n6428);
   U23845 : OAI22_X1 port map( A1 => n25574, A2 => n20935, B1 => n25872, B2 => 
                           n25566, ZN => n6429);
   U23846 : OAI22_X1 port map( A1 => n25574, A2 => n20934, B1 => n25875, B2 => 
                           n25566, ZN => n6430);
   U23847 : OAI22_X1 port map( A1 => n25574, A2 => n20933, B1 => n25878, B2 => 
                           n25566, ZN => n6431);
   U23848 : OAI22_X1 port map( A1 => n25574, A2 => n20932, B1 => n25881, B2 => 
                           n25566, ZN => n6432);
   U23849 : OAI22_X1 port map( A1 => n25574, A2 => n20931, B1 => n25884, B2 => 
                           n25566, ZN => n6433);
   U23850 : OAI22_X1 port map( A1 => n25574, A2 => n20930, B1 => n25887, B2 => 
                           n25566, ZN => n6434);
   U23851 : OAI22_X1 port map( A1 => n25574, A2 => n20929, B1 => n25890, B2 => 
                           n25567, ZN => n6435);
   U23852 : OAI22_X1 port map( A1 => n25574, A2 => n20928, B1 => n25893, B2 => 
                           n25567, ZN => n6436);
   U23853 : OAI22_X1 port map( A1 => n25575, A2 => n20927, B1 => n25896, B2 => 
                           n25567, ZN => n6437);
   U23854 : OAI22_X1 port map( A1 => n25575, A2 => n20926, B1 => n25899, B2 => 
                           n25567, ZN => n6438);
   U23855 : OAI22_X1 port map( A1 => n25575, A2 => n20925, B1 => n25902, B2 => 
                           n25567, ZN => n6439);
   U23856 : OAI22_X1 port map( A1 => n25575, A2 => n20924, B1 => n25905, B2 => 
                           n25567, ZN => n6440);
   U23857 : OAI22_X1 port map( A1 => n25575, A2 => n20923, B1 => n25908, B2 => 
                           n25567, ZN => n6441);
   U23858 : OAI22_X1 port map( A1 => n25575, A2 => n20922, B1 => n25911, B2 => 
                           n25567, ZN => n6442);
   U23859 : OAI22_X1 port map( A1 => n25575, A2 => n20921, B1 => n25914, B2 => 
                           n25567, ZN => n6443);
   U23860 : OAI22_X1 port map( A1 => n25575, A2 => n20920, B1 => n25917, B2 => 
                           n25567, ZN => n6444);
   U23861 : OAI22_X1 port map( A1 => n25575, A2 => n20919, B1 => n25920, B2 => 
                           n25567, ZN => n6445);
   U23862 : OAI22_X1 port map( A1 => n25575, A2 => n20918, B1 => n25923, B2 => 
                           n25567, ZN => n6446);
   U23863 : OAI22_X1 port map( A1 => n25575, A2 => n20917, B1 => n25926, B2 => 
                           n25568, ZN => n6447);
   U23864 : OAI22_X1 port map( A1 => n25575, A2 => n20916, B1 => n25929, B2 => 
                           n25568, ZN => n6448);
   U23865 : OAI22_X1 port map( A1 => n25575, A2 => n20915, B1 => n25932, B2 => 
                           n25568, ZN => n6449);
   U23866 : OAI22_X1 port map( A1 => n25576, A2 => n20914, B1 => n25935, B2 => 
                           n25568, ZN => n6450);
   U23867 : OAI22_X1 port map( A1 => n25576, A2 => n20913, B1 => n25938, B2 => 
                           n25568, ZN => n6451);
   U23868 : OAI22_X1 port map( A1 => n25576, A2 => n20912, B1 => n25941, B2 => 
                           n25568, ZN => n6452);
   U23869 : OAI22_X1 port map( A1 => n25576, A2 => n20911, B1 => n25944, B2 => 
                           n25568, ZN => n6453);
   U23870 : OAI22_X1 port map( A1 => n25576, A2 => n20910, B1 => n25947, B2 => 
                           n25568, ZN => n6454);
   U23871 : OAI22_X1 port map( A1 => n25576, A2 => n20909, B1 => n25950, B2 => 
                           n25568, ZN => n6455);
   U23872 : OAI22_X1 port map( A1 => n25576, A2 => n20908, B1 => n25953, B2 => 
                           n25568, ZN => n6456);
   U23873 : OAI22_X1 port map( A1 => n25576, A2 => n20907, B1 => n25956, B2 => 
                           n25568, ZN => n6457);
   U23874 : OAI22_X1 port map( A1 => n25576, A2 => n20906, B1 => n25959, B2 => 
                           n25568, ZN => n6458);
   U23875 : OAI22_X1 port map( A1 => n25382, A2 => n20777, B1 => n25963, B2 => 
                           n25375, ZN => n5499);
   U23876 : OAI22_X1 port map( A1 => n25382, A2 => n20776, B1 => n25966, B2 => 
                           n25375, ZN => n5500);
   U23877 : OAI22_X1 port map( A1 => n25382, A2 => n20775, B1 => n25969, B2 => 
                           n25375, ZN => n5501);
   U23878 : OAI22_X1 port map( A1 => n25382, A2 => n20774, B1 => n25972, B2 => 
                           n25375, ZN => n5502);
   U23879 : OAI22_X1 port map( A1 => n25675, A2 => n19749, B1 => n25781, B2 => 
                           n25667, ZN => n6911);
   U23880 : OAI22_X1 port map( A1 => n25675, A2 => n19748, B1 => n25784, B2 => 
                           n25667, ZN => n6912);
   U23881 : OAI22_X1 port map( A1 => n25675, A2 => n19747, B1 => n25787, B2 => 
                           n25667, ZN => n6913);
   U23882 : OAI22_X1 port map( A1 => n25675, A2 => n19746, B1 => n25790, B2 => 
                           n25667, ZN => n6914);
   U23883 : OAI22_X1 port map( A1 => n25675, A2 => n19745, B1 => n25793, B2 => 
                           n25667, ZN => n6915);
   U23884 : OAI22_X1 port map( A1 => n25675, A2 => n19744, B1 => n25796, B2 => 
                           n25667, ZN => n6916);
   U23885 : OAI22_X1 port map( A1 => n25675, A2 => n19743, B1 => n25799, B2 => 
                           n25667, ZN => n6917);
   U23886 : OAI22_X1 port map( A1 => n25675, A2 => n19742, B1 => n25802, B2 => 
                           n25667, ZN => n6918);
   U23887 : OAI22_X1 port map( A1 => n25675, A2 => n19741, B1 => n25805, B2 => 
                           n25667, ZN => n6919);
   U23888 : OAI22_X1 port map( A1 => n25675, A2 => n19740, B1 => n25808, B2 => 
                           n25667, ZN => n6920);
   U23889 : OAI22_X1 port map( A1 => n25675, A2 => n19739, B1 => n25811, B2 => 
                           n25667, ZN => n6921);
   U23890 : OAI22_X1 port map( A1 => n25675, A2 => n19738, B1 => n25814, B2 => 
                           n25667, ZN => n6922);
   U23891 : OAI22_X1 port map( A1 => n25676, A2 => n19737, B1 => n25817, B2 => 
                           n25668, ZN => n6923);
   U23892 : OAI22_X1 port map( A1 => n25676, A2 => n19736, B1 => n25820, B2 => 
                           n25668, ZN => n6924);
   U23893 : OAI22_X1 port map( A1 => n25676, A2 => n19735, B1 => n25823, B2 => 
                           n25668, ZN => n6925);
   U23894 : OAI22_X1 port map( A1 => n25676, A2 => n19734, B1 => n25826, B2 => 
                           n25668, ZN => n6926);
   U23895 : OAI22_X1 port map( A1 => n25676, A2 => n19733, B1 => n25829, B2 => 
                           n25668, ZN => n6927);
   U23896 : OAI22_X1 port map( A1 => n25676, A2 => n19732, B1 => n25832, B2 => 
                           n25668, ZN => n6928);
   U23897 : OAI22_X1 port map( A1 => n25676, A2 => n19731, B1 => n25835, B2 => 
                           n25668, ZN => n6929);
   U23898 : OAI22_X1 port map( A1 => n25676, A2 => n19730, B1 => n25838, B2 => 
                           n25668, ZN => n6930);
   U23899 : OAI22_X1 port map( A1 => n25676, A2 => n19729, B1 => n25841, B2 => 
                           n25668, ZN => n6931);
   U23900 : OAI22_X1 port map( A1 => n25676, A2 => n19728, B1 => n25844, B2 => 
                           n25668, ZN => n6932);
   U23901 : OAI22_X1 port map( A1 => n25676, A2 => n19727, B1 => n25847, B2 => 
                           n25668, ZN => n6933);
   U23902 : OAI22_X1 port map( A1 => n25676, A2 => n19726, B1 => n25850, B2 => 
                           n25668, ZN => n6934);
   U23903 : OAI22_X1 port map( A1 => n25676, A2 => n19725, B1 => n25853, B2 => 
                           n25669, ZN => n6935);
   U23904 : OAI22_X1 port map( A1 => n25677, A2 => n19724, B1 => n25856, B2 => 
                           n25669, ZN => n6936);
   U23905 : OAI22_X1 port map( A1 => n25677, A2 => n19723, B1 => n25859, B2 => 
                           n25669, ZN => n6937);
   U23906 : OAI22_X1 port map( A1 => n25677, A2 => n19722, B1 => n25862, B2 => 
                           n25669, ZN => n6938);
   U23907 : OAI22_X1 port map( A1 => n25677, A2 => n19721, B1 => n25865, B2 => 
                           n25669, ZN => n6939);
   U23908 : OAI22_X1 port map( A1 => n25677, A2 => n19720, B1 => n25868, B2 => 
                           n25669, ZN => n6940);
   U23909 : OAI22_X1 port map( A1 => n25677, A2 => n19719, B1 => n25871, B2 => 
                           n25669, ZN => n6941);
   U23910 : OAI22_X1 port map( A1 => n25677, A2 => n19718, B1 => n25874, B2 => 
                           n25669, ZN => n6942);
   U23911 : OAI22_X1 port map( A1 => n25677, A2 => n19717, B1 => n25877, B2 => 
                           n25669, ZN => n6943);
   U23912 : OAI22_X1 port map( A1 => n25677, A2 => n19716, B1 => n25880, B2 => 
                           n25669, ZN => n6944);
   U23913 : OAI22_X1 port map( A1 => n25677, A2 => n19715, B1 => n25883, B2 => 
                           n25669, ZN => n6945);
   U23914 : OAI22_X1 port map( A1 => n25677, A2 => n19714, B1 => n25886, B2 => 
                           n25669, ZN => n6946);
   U23915 : OAI22_X1 port map( A1 => n25677, A2 => n19713, B1 => n25889, B2 => 
                           n25670, ZN => n6947);
   U23916 : OAI22_X1 port map( A1 => n25677, A2 => n19712, B1 => n25892, B2 => 
                           n25670, ZN => n6948);
   U23917 : OAI22_X1 port map( A1 => n25678, A2 => n19711, B1 => n25895, B2 => 
                           n25670, ZN => n6949);
   U23918 : OAI22_X1 port map( A1 => n25678, A2 => n19710, B1 => n25898, B2 => 
                           n25670, ZN => n6950);
   U23919 : OAI22_X1 port map( A1 => n25678, A2 => n19709, B1 => n25901, B2 => 
                           n25670, ZN => n6951);
   U23920 : OAI22_X1 port map( A1 => n25678, A2 => n19708, B1 => n25904, B2 => 
                           n25670, ZN => n6952);
   U23921 : OAI22_X1 port map( A1 => n25678, A2 => n19707, B1 => n25907, B2 => 
                           n25670, ZN => n6953);
   U23922 : OAI22_X1 port map( A1 => n25678, A2 => n19706, B1 => n25910, B2 => 
                           n25670, ZN => n6954);
   U23923 : OAI22_X1 port map( A1 => n25678, A2 => n19705, B1 => n25913, B2 => 
                           n25670, ZN => n6955);
   U23924 : OAI22_X1 port map( A1 => n25678, A2 => n19704, B1 => n25916, B2 => 
                           n25670, ZN => n6956);
   U23925 : OAI22_X1 port map( A1 => n25678, A2 => n19703, B1 => n25919, B2 => 
                           n25670, ZN => n6957);
   U23926 : OAI22_X1 port map( A1 => n25678, A2 => n19702, B1 => n25922, B2 => 
                           n25670, ZN => n6958);
   U23927 : OAI22_X1 port map( A1 => n25678, A2 => n19701, B1 => n25925, B2 => 
                           n25671, ZN => n6959);
   U23928 : OAI22_X1 port map( A1 => n25678, A2 => n19700, B1 => n25928, B2 => 
                           n25671, ZN => n6960);
   U23929 : OAI22_X1 port map( A1 => n25678, A2 => n19699, B1 => n25931, B2 => 
                           n25671, ZN => n6961);
   U23930 : OAI22_X1 port map( A1 => n25679, A2 => n19698, B1 => n25934, B2 => 
                           n25671, ZN => n6962);
   U23931 : OAI22_X1 port map( A1 => n25679, A2 => n19697, B1 => n25937, B2 => 
                           n25671, ZN => n6963);
   U23932 : OAI22_X1 port map( A1 => n25679, A2 => n19696, B1 => n25940, B2 => 
                           n25671, ZN => n6964);
   U23933 : OAI22_X1 port map( A1 => n25679, A2 => n19695, B1 => n25943, B2 => 
                           n25671, ZN => n6965);
   U23934 : OAI22_X1 port map( A1 => n25679, A2 => n19694, B1 => n25946, B2 => 
                           n25671, ZN => n6966);
   U23935 : OAI22_X1 port map( A1 => n25679, A2 => n19693, B1 => n25949, B2 => 
                           n25671, ZN => n6967);
   U23936 : OAI22_X1 port map( A1 => n25679, A2 => n19692, B1 => n25952, B2 => 
                           n25671, ZN => n6968);
   U23937 : OAI22_X1 port map( A1 => n25679, A2 => n19691, B1 => n25955, B2 => 
                           n25671, ZN => n6969);
   U23938 : OAI22_X1 port map( A1 => n25679, A2 => n19690, B1 => n25958, B2 => 
                           n25671, ZN => n6970);
   U23939 : OAI22_X1 port map( A1 => n25482, A2 => n21093, B1 => n25782, B2 => 
                           n25474, ZN => n5951);
   U23940 : OAI22_X1 port map( A1 => n25482, A2 => n21092, B1 => n25785, B2 => 
                           n25474, ZN => n5952);
   U23941 : OAI22_X1 port map( A1 => n25482, A2 => n21091, B1 => n25788, B2 => 
                           n25474, ZN => n5953);
   U23942 : OAI22_X1 port map( A1 => n25482, A2 => n21090, B1 => n25791, B2 => 
                           n25474, ZN => n5954);
   U23943 : OAI22_X1 port map( A1 => n25482, A2 => n21089, B1 => n25794, B2 => 
                           n25474, ZN => n5955);
   U23944 : OAI22_X1 port map( A1 => n25482, A2 => n21088, B1 => n25797, B2 => 
                           n25474, ZN => n5956);
   U23945 : OAI22_X1 port map( A1 => n25482, A2 => n21087, B1 => n25800, B2 => 
                           n25474, ZN => n5957);
   U23946 : OAI22_X1 port map( A1 => n25482, A2 => n21086, B1 => n25803, B2 => 
                           n25474, ZN => n5958);
   U23947 : OAI22_X1 port map( A1 => n25482, A2 => n21085, B1 => n25806, B2 => 
                           n25474, ZN => n5959);
   U23948 : OAI22_X1 port map( A1 => n25482, A2 => n21084, B1 => n25809, B2 => 
                           n25474, ZN => n5960);
   U23949 : OAI22_X1 port map( A1 => n25482, A2 => n21083, B1 => n25812, B2 => 
                           n25474, ZN => n5961);
   U23950 : OAI22_X1 port map( A1 => n25482, A2 => n21082, B1 => n25815, B2 => 
                           n25474, ZN => n5962);
   U23951 : OAI22_X1 port map( A1 => n25483, A2 => n21081, B1 => n25818, B2 => 
                           n25475, ZN => n5963);
   U23952 : OAI22_X1 port map( A1 => n25483, A2 => n21080, B1 => n25821, B2 => 
                           n25475, ZN => n5964);
   U23953 : OAI22_X1 port map( A1 => n25483, A2 => n21079, B1 => n25824, B2 => 
                           n25475, ZN => n5965);
   U23954 : OAI22_X1 port map( A1 => n25483, A2 => n21078, B1 => n25827, B2 => 
                           n25475, ZN => n5966);
   U23955 : OAI22_X1 port map( A1 => n25483, A2 => n21077, B1 => n25830, B2 => 
                           n25475, ZN => n5967);
   U23956 : OAI22_X1 port map( A1 => n25483, A2 => n21076, B1 => n25833, B2 => 
                           n25475, ZN => n5968);
   U23957 : OAI22_X1 port map( A1 => n25483, A2 => n21075, B1 => n25836, B2 => 
                           n25475, ZN => n5969);
   U23958 : OAI22_X1 port map( A1 => n25483, A2 => n21074, B1 => n25839, B2 => 
                           n25475, ZN => n5970);
   U23959 : OAI22_X1 port map( A1 => n25483, A2 => n21073, B1 => n25842, B2 => 
                           n25475, ZN => n5971);
   U23960 : OAI22_X1 port map( A1 => n25483, A2 => n21072, B1 => n25845, B2 => 
                           n25475, ZN => n5972);
   U23961 : OAI22_X1 port map( A1 => n25483, A2 => n21071, B1 => n25848, B2 => 
                           n25475, ZN => n5973);
   U23962 : OAI22_X1 port map( A1 => n25483, A2 => n21070, B1 => n25851, B2 => 
                           n25475, ZN => n5974);
   U23963 : OAI22_X1 port map( A1 => n25483, A2 => n21069, B1 => n25854, B2 => 
                           n25476, ZN => n5975);
   U23964 : OAI22_X1 port map( A1 => n25484, A2 => n21068, B1 => n25857, B2 => 
                           n25476, ZN => n5976);
   U23965 : OAI22_X1 port map( A1 => n25484, A2 => n21067, B1 => n25860, B2 => 
                           n25476, ZN => n5977);
   U23966 : OAI22_X1 port map( A1 => n25484, A2 => n21066, B1 => n25863, B2 => 
                           n25476, ZN => n5978);
   U23967 : OAI22_X1 port map( A1 => n25484, A2 => n21065, B1 => n25866, B2 => 
                           n25476, ZN => n5979);
   U23968 : OAI22_X1 port map( A1 => n25484, A2 => n21064, B1 => n25869, B2 => 
                           n25476, ZN => n5980);
   U23969 : OAI22_X1 port map( A1 => n25484, A2 => n21063, B1 => n25872, B2 => 
                           n25476, ZN => n5981);
   U23970 : OAI22_X1 port map( A1 => n25484, A2 => n21062, B1 => n25875, B2 => 
                           n25476, ZN => n5982);
   U23971 : OAI22_X1 port map( A1 => n25484, A2 => n21061, B1 => n25878, B2 => 
                           n25476, ZN => n5983);
   U23972 : OAI22_X1 port map( A1 => n25484, A2 => n21060, B1 => n25881, B2 => 
                           n25476, ZN => n5984);
   U23973 : OAI22_X1 port map( A1 => n25484, A2 => n21059, B1 => n25884, B2 => 
                           n25476, ZN => n5985);
   U23974 : OAI22_X1 port map( A1 => n25484, A2 => n21058, B1 => n25887, B2 => 
                           n25476, ZN => n5986);
   U23975 : OAI22_X1 port map( A1 => n25484, A2 => n21057, B1 => n25890, B2 => 
                           n25477, ZN => n5987);
   U23976 : OAI22_X1 port map( A1 => n25484, A2 => n21056, B1 => n25893, B2 => 
                           n25477, ZN => n5988);
   U23977 : OAI22_X1 port map( A1 => n25485, A2 => n21055, B1 => n25896, B2 => 
                           n25477, ZN => n5989);
   U23978 : OAI22_X1 port map( A1 => n25485, A2 => n21054, B1 => n25899, B2 => 
                           n25477, ZN => n5990);
   U23979 : OAI22_X1 port map( A1 => n25485, A2 => n21053, B1 => n25902, B2 => 
                           n25477, ZN => n5991);
   U23980 : OAI22_X1 port map( A1 => n25485, A2 => n21052, B1 => n25905, B2 => 
                           n25477, ZN => n5992);
   U23981 : OAI22_X1 port map( A1 => n25485, A2 => n21051, B1 => n25908, B2 => 
                           n25477, ZN => n5993);
   U23982 : OAI22_X1 port map( A1 => n25485, A2 => n21050, B1 => n25911, B2 => 
                           n25477, ZN => n5994);
   U23983 : OAI22_X1 port map( A1 => n25485, A2 => n21049, B1 => n25914, B2 => 
                           n25477, ZN => n5995);
   U23984 : OAI22_X1 port map( A1 => n25485, A2 => n21048, B1 => n25917, B2 => 
                           n25477, ZN => n5996);
   U23985 : OAI22_X1 port map( A1 => n25485, A2 => n21047, B1 => n25920, B2 => 
                           n25477, ZN => n5997);
   U23986 : OAI22_X1 port map( A1 => n25485, A2 => n21046, B1 => n25923, B2 => 
                           n25477, ZN => n5998);
   U23987 : OAI22_X1 port map( A1 => n25485, A2 => n21045, B1 => n25926, B2 => 
                           n25478, ZN => n5999);
   U23988 : OAI22_X1 port map( A1 => n25485, A2 => n21044, B1 => n25929, B2 => 
                           n25478, ZN => n6000);
   U23989 : OAI22_X1 port map( A1 => n25485, A2 => n21043, B1 => n25932, B2 => 
                           n25478, ZN => n6001);
   U23990 : OAI22_X1 port map( A1 => n25486, A2 => n21042, B1 => n25935, B2 => 
                           n25478, ZN => n6002);
   U23991 : OAI22_X1 port map( A1 => n25486, A2 => n21041, B1 => n25938, B2 => 
                           n25478, ZN => n6003);
   U23992 : OAI22_X1 port map( A1 => n25486, A2 => n21040, B1 => n25941, B2 => 
                           n25478, ZN => n6004);
   U23993 : OAI22_X1 port map( A1 => n25486, A2 => n21039, B1 => n25944, B2 => 
                           n25478, ZN => n6005);
   U23994 : OAI22_X1 port map( A1 => n25486, A2 => n21038, B1 => n25947, B2 => 
                           n25478, ZN => n6006);
   U23995 : OAI22_X1 port map( A1 => n25486, A2 => n21037, B1 => n25950, B2 => 
                           n25478, ZN => n6007);
   U23996 : OAI22_X1 port map( A1 => n25486, A2 => n21036, B1 => n25953, B2 => 
                           n25478, ZN => n6008);
   U23997 : OAI22_X1 port map( A1 => n25486, A2 => n21035, B1 => n25956, B2 => 
                           n25478, ZN => n6009);
   U23998 : OAI22_X1 port map( A1 => n25486, A2 => n21034, B1 => n25959, B2 => 
                           n25478, ZN => n6010);
   U23999 : NOR3_X1 port map( A1 => n19493, A2 => ADD_RD2(3), A3 => n19489, ZN 
                           => n23940);
   U24000 : NOR3_X1 port map( A1 => n19488, A2 => ADD_RD1(3), A3 => n19484, ZN 
                           => n22743);
   U24001 : NOR3_X1 port map( A1 => n19493, A2 => ADD_RD2(4), A3 => n19490, ZN 
                           => n23929);
   U24002 : NOR3_X1 port map( A1 => n19488, A2 => ADD_RD1(4), A3 => n19485, ZN 
                           => n22732);
   U24003 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n19493,
                           ZN => n23937);
   U24004 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n19488,
                           ZN => n22740);
   U24005 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n23935);
   U24006 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n22738);
   U24007 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n19489,
                           ZN => n23933);
   U24008 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(3), A3 => n19484,
                           ZN => n22736);
   U24009 : NOR3_X1 port map( A1 => n19489, A2 => ADD_RD2(0), A3 => n19490, ZN 
                           => n23939);
   U24010 : NOR3_X1 port map( A1 => n19484, A2 => ADD_RD1(0), A3 => n19485, ZN 
                           => n22742);
   U24011 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n19490,
                           ZN => n23927);
   U24012 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n19485,
                           ZN => n22730);
   U24013 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), ZN => n21490);
   U24014 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n19483, ZN => n21487);
   U24015 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => n19482, ZN => n21484);
   U24016 : INV_X1 port map( A => ADD_RD2(3), ZN => n19490);
   U24017 : INV_X1 port map( A => ADD_RD1(3), ZN => n19485);
   U24018 : INV_X1 port map( A => ADD_RD2(4), ZN => n19489);
   U24019 : INV_X1 port map( A => ADD_RD1(4), ZN => n19484);
   U24020 : INV_X1 port map( A => ADD_RD2(0), ZN => n19493);
   U24021 : INV_X1 port map( A => ADD_RD1(0), ZN => n19488);
   U24022 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => ADD_WR(4), ZN => 
                           n21528);
   U24023 : AND3_X1 port map( A1 => ENABLE, A2 => n19479, A3 => WR, ZN => 
                           n21491);
   U24024 : INV_X1 port map( A => ADD_WR(4), ZN => n19479);
   U24025 : INV_X1 port map( A => RESET, ZN => n19478);
   U24026 : INV_X1 port map( A => DATAIN(0), ZN => n19557);
   U24027 : INV_X1 port map( A => DATAIN(1), ZN => n19556);
   U24028 : INV_X1 port map( A => DATAIN(2), ZN => n19555);
   U24029 : INV_X1 port map( A => DATAIN(3), ZN => n19554);
   U24030 : INV_X1 port map( A => DATAIN(4), ZN => n19553);
   U24031 : INV_X1 port map( A => DATAIN(5), ZN => n19552);
   U24032 : INV_X1 port map( A => DATAIN(6), ZN => n19551);
   U24033 : INV_X1 port map( A => DATAIN(7), ZN => n19550);
   U24034 : INV_X1 port map( A => DATAIN(8), ZN => n19549);
   U24035 : INV_X1 port map( A => DATAIN(9), ZN => n19548);
   U24036 : INV_X1 port map( A => DATAIN(10), ZN => n19547);
   U24037 : INV_X1 port map( A => DATAIN(11), ZN => n19546);
   U24038 : INV_X1 port map( A => DATAIN(12), ZN => n19545);
   U24039 : INV_X1 port map( A => DATAIN(13), ZN => n19544);
   U24040 : INV_X1 port map( A => DATAIN(14), ZN => n19543);
   U24041 : INV_X1 port map( A => DATAIN(15), ZN => n19542);
   U24042 : INV_X1 port map( A => DATAIN(16), ZN => n19541);
   U24043 : INV_X1 port map( A => DATAIN(17), ZN => n19540);
   U24044 : INV_X1 port map( A => DATAIN(18), ZN => n19539);
   U24045 : INV_X1 port map( A => DATAIN(19), ZN => n19538);
   U24046 : INV_X1 port map( A => DATAIN(20), ZN => n19537);
   U24047 : INV_X1 port map( A => DATAIN(21), ZN => n19536);
   U24048 : INV_X1 port map( A => DATAIN(22), ZN => n19535);
   U24049 : INV_X1 port map( A => DATAIN(23), ZN => n19534);
   U24050 : INV_X1 port map( A => DATAIN(24), ZN => n19533);
   U24051 : INV_X1 port map( A => DATAIN(25), ZN => n19532);
   U24052 : INV_X1 port map( A => DATAIN(26), ZN => n19531);
   U24053 : INV_X1 port map( A => DATAIN(27), ZN => n19530);
   U24054 : INV_X1 port map( A => DATAIN(28), ZN => n19529);
   U24055 : INV_X1 port map( A => DATAIN(29), ZN => n19528);
   U24056 : INV_X1 port map( A => DATAIN(30), ZN => n19527);
   U24057 : INV_X1 port map( A => DATAIN(31), ZN => n19526);
   U24058 : INV_X1 port map( A => DATAIN(32), ZN => n19525);
   U24059 : INV_X1 port map( A => DATAIN(33), ZN => n19524);
   U24060 : INV_X1 port map( A => DATAIN(34), ZN => n19523);
   U24061 : INV_X1 port map( A => DATAIN(35), ZN => n19522);
   U24062 : INV_X1 port map( A => DATAIN(36), ZN => n19521);
   U24063 : INV_X1 port map( A => DATAIN(37), ZN => n19520);
   U24064 : INV_X1 port map( A => DATAIN(38), ZN => n19519);
   U24065 : INV_X1 port map( A => DATAIN(39), ZN => n19518);
   U24066 : INV_X1 port map( A => DATAIN(40), ZN => n19517);
   U24067 : INV_X1 port map( A => DATAIN(41), ZN => n19516);
   U24068 : INV_X1 port map( A => DATAIN(42), ZN => n19515);
   U24069 : INV_X1 port map( A => DATAIN(43), ZN => n19514);
   U24070 : INV_X1 port map( A => DATAIN(44), ZN => n19513);
   U24071 : INV_X1 port map( A => DATAIN(45), ZN => n19512);
   U24072 : INV_X1 port map( A => DATAIN(46), ZN => n19511);
   U24073 : INV_X1 port map( A => DATAIN(47), ZN => n19510);
   U24074 : INV_X1 port map( A => DATAIN(48), ZN => n19509);
   U24075 : INV_X1 port map( A => DATAIN(49), ZN => n19508);
   U24076 : INV_X1 port map( A => DATAIN(50), ZN => n19507);
   U24077 : INV_X1 port map( A => DATAIN(51), ZN => n19506);
   U24078 : INV_X1 port map( A => DATAIN(52), ZN => n19505);
   U24079 : INV_X1 port map( A => DATAIN(53), ZN => n19504);
   U24080 : INV_X1 port map( A => DATAIN(54), ZN => n19503);
   U24081 : INV_X1 port map( A => DATAIN(55), ZN => n19502);
   U24082 : INV_X1 port map( A => DATAIN(56), ZN => n19501);
   U24083 : INV_X1 port map( A => DATAIN(57), ZN => n19500);
   U24084 : INV_X1 port map( A => DATAIN(58), ZN => n19499);
   U24085 : INV_X1 port map( A => DATAIN(59), ZN => n19498);
   U24086 : INV_X1 port map( A => DATAIN(60), ZN => n19497);
   U24087 : INV_X1 port map( A => DATAIN(61), ZN => n19496);
   U24088 : INV_X1 port map( A => DATAIN(62), ZN => n19495);
   U24089 : INV_X1 port map( A => DATAIN(63), ZN => n19494);
   U24090 : INV_X1 port map( A => ADD_WR(3), ZN => n19480);
   U24091 : INV_X1 port map( A => ADD_WR(2), ZN => n19481);
   U24092 : INV_X1 port map( A => ADD_WR(0), ZN => n19483);
   U24093 : INV_X1 port map( A => ADD_RD2(2), ZN => n19491);
   U24094 : INV_X1 port map( A => ADD_RD1(2), ZN => n19486);
   U24095 : INV_X1 port map( A => ADD_RD2(1), ZN => n19492);
   U24096 : INV_X1 port map( A => ADD_RD1(1), ZN => n19487);
   U24097 : INV_X1 port map( A => ADD_WR(1), ZN => n19482);
   U24098 : CLKBUF_X1 port map( A => n22803, Z => n24979);
   U24099 : CLKBUF_X1 port map( A => n22802, Z => n24985);
   U24100 : CLKBUF_X1 port map( A => n22800, Z => n24991);
   U24101 : CLKBUF_X1 port map( A => n22799, Z => n24997);
   U24102 : CLKBUF_X1 port map( A => n22798, Z => n25003);
   U24103 : CLKBUF_X1 port map( A => n22797, Z => n25009);
   U24104 : CLKBUF_X1 port map( A => n22795, Z => n25015);
   U24105 : CLKBUF_X1 port map( A => n22794, Z => n25021);
   U24106 : CLKBUF_X1 port map( A => n22793, Z => n25027);
   U24107 : CLKBUF_X1 port map( A => n22792, Z => n25033);
   U24108 : CLKBUF_X1 port map( A => n22790, Z => n25039);
   U24109 : CLKBUF_X1 port map( A => n22789, Z => n25045);
   U24110 : CLKBUF_X1 port map( A => n22788, Z => n25051);
   U24111 : CLKBUF_X1 port map( A => n22787, Z => n25057);
   U24112 : CLKBUF_X1 port map( A => n22785, Z => n25063);
   U24113 : CLKBUF_X1 port map( A => n22784, Z => n25069);
   U24114 : CLKBUF_X1 port map( A => n22779, Z => n25075);
   U24115 : CLKBUF_X1 port map( A => n22778, Z => n25081);
   U24116 : CLKBUF_X1 port map( A => n22777, Z => n25087);
   U24117 : CLKBUF_X1 port map( A => n22775, Z => n25093);
   U24118 : CLKBUF_X1 port map( A => n22774, Z => n25099);
   U24119 : CLKBUF_X1 port map( A => n22773, Z => n25105);
   U24120 : CLKBUF_X1 port map( A => n22772, Z => n25111);
   U24121 : CLKBUF_X1 port map( A => n22770, Z => n25117);
   U24122 : CLKBUF_X1 port map( A => n22769, Z => n25123);
   U24123 : CLKBUF_X1 port map( A => n22768, Z => n25129);
   U24124 : CLKBUF_X1 port map( A => n22767, Z => n25135);
   U24125 : CLKBUF_X1 port map( A => n22765, Z => n25141);
   U24126 : CLKBUF_X1 port map( A => n22764, Z => n25147);
   U24127 : CLKBUF_X1 port map( A => n22763, Z => n25153);
   U24128 : CLKBUF_X1 port map( A => n22762, Z => n25159);
   U24129 : CLKBUF_X1 port map( A => n22760, Z => n25165);
   U24130 : CLKBUF_X1 port map( A => n22759, Z => n25171);
   U24131 : CLKBUF_X1 port map( A => n21606, Z => n25177);
   U24132 : CLKBUF_X1 port map( A => n21605, Z => n25183);
   U24133 : CLKBUF_X1 port map( A => n21603, Z => n25189);
   U24134 : CLKBUF_X1 port map( A => n21602, Z => n25195);
   U24135 : CLKBUF_X1 port map( A => n21601, Z => n25201);
   U24136 : CLKBUF_X1 port map( A => n21600, Z => n25207);
   U24137 : CLKBUF_X1 port map( A => n21598, Z => n25213);
   U24138 : CLKBUF_X1 port map( A => n21597, Z => n25219);
   U24139 : CLKBUF_X1 port map( A => n21596, Z => n25225);
   U24140 : CLKBUF_X1 port map( A => n21595, Z => n25231);
   U24141 : CLKBUF_X1 port map( A => n21593, Z => n25237);
   U24142 : CLKBUF_X1 port map( A => n21592, Z => n25243);
   U24143 : CLKBUF_X1 port map( A => n21591, Z => n25249);
   U24144 : CLKBUF_X1 port map( A => n21590, Z => n25255);
   U24145 : CLKBUF_X1 port map( A => n21588, Z => n25261);
   U24146 : CLKBUF_X1 port map( A => n21587, Z => n25267);
   U24147 : CLKBUF_X1 port map( A => n21582, Z => n25273);
   U24148 : CLKBUF_X1 port map( A => n21581, Z => n25279);
   U24149 : CLKBUF_X1 port map( A => n21580, Z => n25285);
   U24150 : CLKBUF_X1 port map( A => n21578, Z => n25291);
   U24151 : CLKBUF_X1 port map( A => n21577, Z => n25297);
   U24152 : CLKBUF_X1 port map( A => n21576, Z => n25303);
   U24153 : CLKBUF_X1 port map( A => n21575, Z => n25309);
   U24154 : CLKBUF_X1 port map( A => n21573, Z => n25315);
   U24155 : CLKBUF_X1 port map( A => n21572, Z => n25321);
   U24156 : CLKBUF_X1 port map( A => n21571, Z => n25327);
   U24157 : CLKBUF_X1 port map( A => n21570, Z => n25333);
   U24158 : CLKBUF_X1 port map( A => n21568, Z => n25339);
   U24159 : CLKBUF_X1 port map( A => n21567, Z => n25345);
   U24160 : CLKBUF_X1 port map( A => n21566, Z => n25351);
   U24161 : CLKBUF_X1 port map( A => n21565, Z => n25357);
   U24162 : CLKBUF_X1 port map( A => n21563, Z => n25363);
   U24163 : CLKBUF_X1 port map( A => n21562, Z => n25369);
   U24164 : CLKBUF_X1 port map( A => n21555, Z => n25375);
   U24165 : CLKBUF_X1 port map( A => n21553, Z => n25388);
   U24166 : CLKBUF_X1 port map( A => n21551, Z => n25401);
   U24167 : CLKBUF_X1 port map( A => n21548, Z => n25414);
   U24168 : CLKBUF_X1 port map( A => n21546, Z => n25427);
   U24169 : CLKBUF_X1 port map( A => n21544, Z => n25440);
   U24170 : CLKBUF_X1 port map( A => n21542, Z => n25453);
   U24171 : CLKBUF_X1 port map( A => n21539, Z => n25466);
   U24172 : CLKBUF_X1 port map( A => n21537, Z => n25479);
   U24173 : CLKBUF_X1 port map( A => n21535, Z => n25492);
   U24174 : CLKBUF_X1 port map( A => n21533, Z => n25505);
   U24175 : CLKBUF_X1 port map( A => n21532, Z => n25511);
   U24176 : CLKBUF_X1 port map( A => n21530, Z => n25517);
   U24177 : CLKBUF_X1 port map( A => n21527, Z => n25530);
   U24178 : CLKBUF_X1 port map( A => n21525, Z => n25543);
   U24179 : CLKBUF_X1 port map( A => n21523, Z => n25556);
   U24180 : CLKBUF_X1 port map( A => n21520, Z => n25569);
   U24181 : CLKBUF_X1 port map( A => n21518, Z => n25582);
   U24182 : CLKBUF_X1 port map( A => n21517, Z => n25588);
   U24183 : CLKBUF_X1 port map( A => n21516, Z => n25594);
   U24184 : CLKBUF_X1 port map( A => n21514, Z => n25607);
   U24185 : CLKBUF_X1 port map( A => n21511, Z => n25620);
   U24186 : CLKBUF_X1 port map( A => n21509, Z => n25633);
   U24187 : CLKBUF_X1 port map( A => n21507, Z => n25646);
   U24188 : CLKBUF_X1 port map( A => n21505, Z => n25659);
   U24189 : CLKBUF_X1 port map( A => n21502, Z => n25672);
   U24190 : CLKBUF_X1 port map( A => n21500, Z => n25685);
   U24191 : CLKBUF_X1 port map( A => n21499, Z => n25691);
   U24192 : CLKBUF_X1 port map( A => n21498, Z => n25697);
   U24193 : CLKBUF_X1 port map( A => n21496, Z => n25710);
   U24194 : CLKBUF_X1 port map( A => n21493, Z => n25723);
   U24195 : CLKBUF_X1 port map( A => n21489, Z => n25736);
   U24196 : CLKBUF_X1 port map( A => n21486, Z => n25749);
   U24197 : CLKBUF_X1 port map( A => n21485, Z => n25755);
   U24198 : CLKBUF_X1 port map( A => n21483, Z => n25761);
   U24199 : CLKBUF_X1 port map( A => n21479, Z => n25774);
   U24200 : CLKBUF_X1 port map( A => n21478, Z => n25780);
   U24201 : CLKBUF_X1 port map( A => n19478, Z => n25978);

end SYN_A;
