
module register_file_NBIT64_NREG32 ( CLK, RESET, ENABLE, RD1, RD2, WR, ADD_WR, 
        ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [63:0] DATAIN;
  output [63:0] OUT1;
  output [63:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7149, n7150, n7151, n7152, n7153, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7490, n7491, n7492, n7493, n7494,
         n7495, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7653, n7654, n7655, n7656, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4642,
         n4643, n4646, n4647, n4648, n4649, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4682, n4683, n4684, n4685, n7080, n7081, n7084,
         n7085, n7088, n7089, n7092, n7093, n7096, n7097, n7100, n7101, n7104,
         n7105, n7130, n7131, n7154, n7155, n7158, n7159, n7162, n7163, n7166,
         n7167, n7170, n7171, n7174, n7175, n7178, n7179, n7182, n7183, n7186,
         n7187, n7190, n7191, n7194, n7195, n7198, n7199, n7202, n7205, n7208,
         n7211, n7214, n7217, n7220, n7223, n7226, n7229, n7232, n7245, n7278,
         n7279, n7282, n7283, n7286, n7287, n7290, n7291, n7294, n7295, n7298,
         n7299, n7302, n7303, n7306, n7307, n7310, n7311, n7314, n7315, n7318,
         n7319, n7322, n7323, n8599, n8600, n8603, n8604, n8605, n8606, n8611,
         n8612, n8613, n8614, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466;

  DFF_X1 \REGISTERS_reg[0][63]  ( .D(n7037), .CK(CLK), .QN(n13392) );
  DFF_X1 \REGISTERS_reg[0][54]  ( .D(n7028), .CK(CLK), .QN(n13393) );
  DFF_X1 \REGISTERS_reg[0][53]  ( .D(n7027), .CK(CLK), .QN(n13394) );
  DFF_X1 \REGISTERS_reg[0][52]  ( .D(n7026), .CK(CLK), .QN(n13395) );
  DFF_X1 \REGISTERS_reg[0][51]  ( .D(n7025), .CK(CLK), .QN(n13396) );
  DFF_X1 \REGISTERS_reg[0][50]  ( .D(n7024), .CK(CLK), .QN(n13397) );
  DFF_X1 \REGISTERS_reg[0][49]  ( .D(n7023), .CK(CLK), .QN(n13398) );
  DFF_X1 \REGISTERS_reg[0][48]  ( .D(n7022), .CK(CLK), .QN(n13399) );
  DFF_X1 \REGISTERS_reg[0][47]  ( .D(n7021), .CK(CLK), .QN(n13400) );
  DFF_X1 \REGISTERS_reg[0][46]  ( .D(n7020), .CK(CLK), .QN(n13401) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n6938), .CK(CLK), .QN(n13402) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n6937), .CK(CLK), .QN(n13403) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n6936), .CK(CLK), .QN(n13404) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n6935), .CK(CLK), .QN(n13405) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n6934), .CK(CLK), .QN(n13406) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n6933), .CK(CLK), .QN(n13407) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n6932), .CK(CLK), .QN(n13408) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n6931), .CK(CLK), .QN(n13409) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n6930), .CK(CLK), .QN(n13410) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n6929), .CK(CLK), .QN(n13411) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n6928), .CK(CLK), .QN(n13412) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n6927), .CK(CLK), .QN(n13413) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n6926), .CK(CLK), .QN(n13414) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n6925), .CK(CLK), .QN(n13415) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n6924), .CK(CLK), .QN(n13416) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n6923), .CK(CLK), .QN(n13417) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n6922), .CK(CLK), .QN(n13418) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n6921), .CK(CLK), .QN(n13419) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n6920), .CK(CLK), .QN(n13420) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n6919), .CK(CLK), .QN(n13421) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n6918), .CK(CLK), .QN(n13422) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n6917), .CK(CLK), .QN(n13423) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n6916), .CK(CLK), .QN(n13424) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n6915), .CK(CLK), .QN(n13425) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n6914), .CK(CLK), .QN(n13426) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n6913), .CK(CLK), .QN(n13427) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n6912), .CK(CLK), .QN(n13428) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n6911), .CK(CLK), .QN(n13429) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n6910), .CK(CLK), .QN(n13430) );
  DFF_X1 \REGISTERS_reg[10][59]  ( .D(n6393), .CK(CLK), .QN(n13435) );
  DFF_X1 \REGISTERS_reg[10][58]  ( .D(n6392), .CK(CLK), .QN(n13436) );
  DFF_X1 \REGISTERS_reg[10][57]  ( .D(n6391), .CK(CLK), .QN(n13437) );
  DFF_X1 \REGISTERS_reg[10][56]  ( .D(n6390), .CK(CLK), .QN(n13438) );
  DFF_X1 \REGISTERS_reg[10][55]  ( .D(n6389), .CK(CLK), .QN(n13439) );
  DFF_X1 \REGISTERS_reg[10][54]  ( .D(n6388), .CK(CLK), .QN(n13440) );
  DFF_X1 \REGISTERS_reg[10][53]  ( .D(n6387), .CK(CLK), .QN(n13441) );
  DFF_X1 \REGISTERS_reg[10][52]  ( .D(n6386), .CK(CLK), .QN(n13442) );
  DFF_X1 \REGISTERS_reg[10][51]  ( .D(n6385), .CK(CLK), .QN(n13443) );
  DFF_X1 \REGISTERS_reg[10][50]  ( .D(n6384), .CK(CLK), .QN(n13444) );
  DFF_X1 \REGISTERS_reg[10][49]  ( .D(n6383), .CK(CLK), .QN(n13445) );
  DFF_X1 \REGISTERS_reg[10][48]  ( .D(n6382), .CK(CLK), .QN(n13446) );
  DFF_X1 \REGISTERS_reg[10][47]  ( .D(n6381), .CK(CLK), .QN(n13447) );
  DFF_X1 \REGISTERS_reg[10][46]  ( .D(n6380), .CK(CLK), .QN(n13448) );
  DFF_X1 \REGISTERS_reg[10][45]  ( .D(n6379), .CK(CLK), .QN(n13449) );
  DFF_X1 \REGISTERS_reg[10][44]  ( .D(n6378), .CK(CLK), .QN(n13450) );
  DFF_X1 \REGISTERS_reg[10][43]  ( .D(n6377), .CK(CLK), .QN(n13451) );
  DFF_X1 \REGISTERS_reg[10][42]  ( .D(n6376), .CK(CLK), .QN(n13452) );
  DFF_X1 \REGISTERS_reg[10][41]  ( .D(n6375), .CK(CLK), .QN(n13453) );
  DFF_X1 \REGISTERS_reg[10][40]  ( .D(n6374), .CK(CLK), .QN(n13454) );
  DFF_X1 \REGISTERS_reg[10][39]  ( .D(n6373), .CK(CLK), .QN(n13455) );
  DFF_X1 \REGISTERS_reg[10][38]  ( .D(n6372), .CK(CLK), .QN(n13456) );
  DFF_X1 \REGISTERS_reg[10][37]  ( .D(n6371), .CK(CLK), .QN(n13457) );
  DFF_X1 \REGISTERS_reg[10][36]  ( .D(n6370), .CK(CLK), .QN(n13458) );
  DFF_X1 \REGISTERS_reg[10][35]  ( .D(n6369), .CK(CLK), .QN(n13459) );
  DFF_X1 \REGISTERS_reg[10][34]  ( .D(n6368), .CK(CLK), .QN(n13460) );
  DFF_X1 \REGISTERS_reg[10][33]  ( .D(n6367), .CK(CLK), .QN(n13461) );
  DFF_X1 \REGISTERS_reg[10][32]  ( .D(n6366), .CK(CLK), .QN(n13462) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n6365), .CK(CLK), .QN(n13463) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n6364), .CK(CLK), .QN(n13464) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n6363), .CK(CLK), .QN(n13465) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n6362), .CK(CLK), .QN(n13466) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n6361), .CK(CLK), .QN(n13467) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n6360), .CK(CLK), .QN(n13468) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n6359), .CK(CLK), .QN(n13469) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n6358), .CK(CLK), .QN(n13470) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n6357), .CK(CLK), .QN(n13471) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n6356), .CK(CLK), .QN(n13472) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n6355), .CK(CLK), .QN(n13473) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n6354), .CK(CLK), .QN(n13474) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n6353), .CK(CLK), .QN(n13475) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n6352), .CK(CLK), .QN(n13476) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n6351), .CK(CLK), .QN(n13477) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n6350), .CK(CLK), .QN(n13478) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n6349), .CK(CLK), .QN(n13479) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n6348), .CK(CLK), .QN(n13480) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n6347), .CK(CLK), .QN(n13481) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n6346), .CK(CLK), .QN(n13482) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n6345), .CK(CLK), .QN(n13483) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n6344), .CK(CLK), .QN(n13484) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n6343), .CK(CLK), .QN(n13485) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n6342), .CK(CLK), .QN(n13486) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n6341), .CK(CLK), .QN(n13487) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n6340), .CK(CLK), .QN(n13488) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n6339), .CK(CLK), .QN(n13489) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n6338), .CK(CLK), .QN(n13490) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n6337), .CK(CLK), .QN(n13491) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n6336), .CK(CLK), .QN(n13492) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n6335), .CK(CLK), .QN(n13493) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n6334), .CK(CLK), .QN(n13494) );
  DFF_X1 \REGISTERS_reg[11][59]  ( .D(n6329), .CK(CLK), .QN(n13499) );
  DFF_X1 \REGISTERS_reg[11][58]  ( .D(n6328), .CK(CLK), .QN(n13500) );
  DFF_X1 \REGISTERS_reg[11][57]  ( .D(n6327), .CK(CLK), .QN(n13501) );
  DFF_X1 \REGISTERS_reg[11][56]  ( .D(n6326), .CK(CLK), .QN(n13502) );
  DFF_X1 \REGISTERS_reg[11][55]  ( .D(n6325), .CK(CLK), .QN(n13503) );
  DFF_X1 \REGISTERS_reg[11][54]  ( .D(n6324), .CK(CLK), .QN(n13504) );
  DFF_X1 \REGISTERS_reg[11][53]  ( .D(n6323), .CK(CLK), .QN(n13505) );
  DFF_X1 \REGISTERS_reg[11][52]  ( .D(n6322), .CK(CLK), .QN(n13506) );
  DFF_X1 \REGISTERS_reg[11][51]  ( .D(n6321), .CK(CLK), .QN(n13507) );
  DFF_X1 \REGISTERS_reg[11][50]  ( .D(n6320), .CK(CLK), .QN(n13508) );
  DFF_X1 \REGISTERS_reg[11][49]  ( .D(n6319), .CK(CLK), .QN(n13509) );
  DFF_X1 \REGISTERS_reg[11][48]  ( .D(n6318), .CK(CLK), .QN(n13510) );
  DFF_X1 \REGISTERS_reg[11][47]  ( .D(n6317), .CK(CLK), .QN(n13511) );
  DFF_X1 \REGISTERS_reg[11][46]  ( .D(n6316), .CK(CLK), .QN(n13512) );
  DFF_X1 \REGISTERS_reg[11][45]  ( .D(n6315), .CK(CLK), .QN(n13513) );
  DFF_X1 \REGISTERS_reg[11][44]  ( .D(n6314), .CK(CLK), .QN(n13514) );
  DFF_X1 \REGISTERS_reg[11][43]  ( .D(n6313), .CK(CLK), .QN(n13515) );
  DFF_X1 \REGISTERS_reg[11][38]  ( .D(n6308), .CK(CLK), .QN(n13516) );
  DFF_X1 \REGISTERS_reg[11][37]  ( .D(n6307), .CK(CLK), .QN(n13517) );
  DFF_X1 \REGISTERS_reg[11][36]  ( .D(n6306), .CK(CLK), .QN(n13518) );
  DFF_X1 \REGISTERS_reg[11][35]  ( .D(n6305), .CK(CLK), .QN(n13519) );
  DFF_X1 \REGISTERS_reg[11][34]  ( .D(n6304), .CK(CLK), .QN(n13520) );
  DFF_X1 \REGISTERS_reg[11][33]  ( .D(n6303), .CK(CLK), .QN(n13521) );
  DFF_X1 \REGISTERS_reg[11][32]  ( .D(n6302), .CK(CLK), .QN(n13522) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n6301), .CK(CLK), .QN(n13523) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n6300), .CK(CLK), .QN(n13524) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n6299), .CK(CLK), .QN(n13525) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n6298), .CK(CLK), .QN(n13526) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n6297), .CK(CLK), .QN(n13527) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n6296), .CK(CLK), .QN(n13528) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n6295), .CK(CLK), .QN(n13529) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n6294), .CK(CLK), .QN(n13530) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n6293), .CK(CLK), .QN(n13531) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n6292), .CK(CLK), .QN(n13532) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n6291), .CK(CLK), .QN(n13533) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n6290), .CK(CLK), .QN(n13534) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n6286), .CK(CLK), .QN(n13535) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n6273), .CK(CLK), .QN(n13536) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n6272), .CK(CLK), .QN(n13537) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n6271), .CK(CLK), .QN(n13538) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n6270), .CK(CLK), .QN(n13539) );
  DFF_X1 \REGISTERS_reg[14][59]  ( .D(n6137), .CK(CLK), .QN(n13544) );
  DFF_X1 \REGISTERS_reg[14][58]  ( .D(n6136), .CK(CLK), .QN(n13545) );
  DFF_X1 \REGISTERS_reg[14][57]  ( .D(n6135), .CK(CLK), .QN(n13546) );
  DFF_X1 \REGISTERS_reg[14][56]  ( .D(n6134), .CK(CLK), .QN(n13547) );
  DFF_X1 \REGISTERS_reg[14][55]  ( .D(n6133), .CK(CLK), .QN(n13548) );
  DFF_X1 \REGISTERS_reg[14][54]  ( .D(n6132), .CK(CLK), .QN(n13549) );
  DFF_X1 \REGISTERS_reg[14][53]  ( .D(n6131), .CK(CLK), .QN(n13550) );
  DFF_X1 \REGISTERS_reg[14][52]  ( .D(n6130), .CK(CLK), .QN(n13551) );
  DFF_X1 \REGISTERS_reg[14][51]  ( .D(n6129), .CK(CLK), .QN(n13552) );
  DFF_X1 \REGISTERS_reg[14][50]  ( .D(n6128), .CK(CLK), .QN(n13553) );
  DFF_X1 \REGISTERS_reg[14][49]  ( .D(n6127), .CK(CLK), .QN(n13554) );
  DFF_X1 \REGISTERS_reg[14][48]  ( .D(n6126), .CK(CLK), .QN(n13555) );
  DFF_X1 \REGISTERS_reg[14][47]  ( .D(n6125), .CK(CLK), .QN(n13556) );
  DFF_X1 \REGISTERS_reg[14][46]  ( .D(n6124), .CK(CLK), .QN(n13557) );
  DFF_X1 \REGISTERS_reg[14][45]  ( .D(n6123), .CK(CLK), .QN(n13558) );
  DFF_X1 \REGISTERS_reg[14][44]  ( .D(n6122), .CK(CLK), .QN(n13559) );
  DFF_X1 \REGISTERS_reg[14][43]  ( .D(n6121), .CK(CLK), .QN(n13560) );
  DFF_X1 \REGISTERS_reg[14][42]  ( .D(n6120), .CK(CLK), .QN(n13561) );
  DFF_X1 \REGISTERS_reg[14][41]  ( .D(n6119), .CK(CLK), .QN(n13562) );
  DFF_X1 \REGISTERS_reg[14][40]  ( .D(n6118), .CK(CLK), .QN(n13563) );
  DFF_X1 \REGISTERS_reg[14][39]  ( .D(n6117), .CK(CLK), .QN(n13564) );
  DFF_X1 \REGISTERS_reg[14][38]  ( .D(n6116), .CK(CLK), .QN(n13565) );
  DFF_X1 \REGISTERS_reg[14][37]  ( .D(n6115), .CK(CLK), .QN(n13566) );
  DFF_X1 \REGISTERS_reg[14][36]  ( .D(n6114), .CK(CLK), .QN(n13567) );
  DFF_X1 \REGISTERS_reg[14][35]  ( .D(n6113), .CK(CLK), .QN(n13568) );
  DFF_X1 \REGISTERS_reg[14][34]  ( .D(n6112), .CK(CLK), .QN(n13569) );
  DFF_X1 \REGISTERS_reg[14][33]  ( .D(n6111), .CK(CLK), .QN(n13570) );
  DFF_X1 \REGISTERS_reg[14][32]  ( .D(n6110), .CK(CLK), .QN(n13571) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n6109), .CK(CLK), .QN(n13572) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n6108), .CK(CLK), .QN(n13573) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n6107), .CK(CLK), .QN(n13574) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n6106), .CK(CLK), .QN(n13575) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n6105), .CK(CLK), .QN(n13576) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n6104), .CK(CLK), .QN(n13577) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n6103), .CK(CLK), .QN(n13578) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n6102), .CK(CLK), .QN(n13579) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n6101), .CK(CLK), .QN(n13580) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n6100), .CK(CLK), .QN(n13581) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n6099), .CK(CLK), .QN(n13582) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n6098), .CK(CLK), .QN(n13583) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n6097), .CK(CLK), .QN(n13584) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n6096), .CK(CLK), .QN(n13585) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n6095), .CK(CLK), .QN(n13586) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n6094), .CK(CLK), .QN(n13587) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n6093), .CK(CLK), .QN(n13588) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n6092), .CK(CLK), .QN(n13589) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n6091), .CK(CLK), .QN(n13590) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n6090), .CK(CLK), .QN(n13591) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n6089), .CK(CLK), .QN(n13592) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n6088), .CK(CLK), .QN(n13593) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n6087), .CK(CLK), .QN(n13594) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n6086), .CK(CLK), .QN(n13595) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n6085), .CK(CLK), .QN(n13596) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n6084), .CK(CLK), .QN(n13597) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n6083), .CK(CLK), .QN(n13598) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n6082), .CK(CLK), .QN(n13599) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n6081), .CK(CLK), .QN(n13600) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n6080), .CK(CLK), .QN(n13601) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n6079), .CK(CLK), .QN(n13602) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n6078), .CK(CLK), .QN(n13603) );
  DFF_X1 \REGISTERS_reg[15][59]  ( .D(n6073), .CK(CLK), .QN(n13608) );
  DFF_X1 \REGISTERS_reg[15][58]  ( .D(n6072), .CK(CLK), .QN(n13609) );
  DFF_X1 \REGISTERS_reg[15][57]  ( .D(n6071), .CK(CLK), .QN(n13610) );
  DFF_X1 \REGISTERS_reg[15][56]  ( .D(n6070), .CK(CLK), .QN(n13611) );
  DFF_X1 \REGISTERS_reg[15][55]  ( .D(n6069), .CK(CLK), .QN(n13612) );
  DFF_X1 \REGISTERS_reg[15][54]  ( .D(n6068), .CK(CLK), .QN(n13613) );
  DFF_X1 \REGISTERS_reg[15][53]  ( .D(n6067), .CK(CLK), .QN(n13614) );
  DFF_X1 \REGISTERS_reg[15][52]  ( .D(n6066), .CK(CLK), .QN(n13615) );
  DFF_X1 \REGISTERS_reg[15][51]  ( .D(n6065), .CK(CLK), .QN(n13616) );
  DFF_X1 \REGISTERS_reg[15][50]  ( .D(n6064), .CK(CLK), .QN(n13617) );
  DFF_X1 \REGISTERS_reg[15][49]  ( .D(n6063), .CK(CLK), .QN(n13618) );
  DFF_X1 \REGISTERS_reg[15][48]  ( .D(n6062), .CK(CLK), .QN(n13619) );
  DFF_X1 \REGISTERS_reg[15][47]  ( .D(n6061), .CK(CLK), .QN(n13620) );
  DFF_X1 \REGISTERS_reg[15][46]  ( .D(n6060), .CK(CLK), .QN(n13621) );
  DFF_X1 \REGISTERS_reg[15][45]  ( .D(n6059), .CK(CLK), .QN(n13622) );
  DFF_X1 \REGISTERS_reg[15][44]  ( .D(n6058), .CK(CLK), .QN(n13623) );
  DFF_X1 \REGISTERS_reg[15][43]  ( .D(n6057), .CK(CLK), .QN(n13624) );
  DFF_X1 \REGISTERS_reg[15][42]  ( .D(n6056), .CK(CLK), .QN(n13625) );
  DFF_X1 \REGISTERS_reg[15][41]  ( .D(n6055), .CK(CLK), .QN(n13626) );
  DFF_X1 \REGISTERS_reg[15][40]  ( .D(n6054), .CK(CLK), .QN(n13627) );
  DFF_X1 \REGISTERS_reg[15][39]  ( .D(n6053), .CK(CLK), .QN(n13628) );
  DFF_X1 \REGISTERS_reg[15][38]  ( .D(n6052), .CK(CLK), .QN(n13629) );
  DFF_X1 \REGISTERS_reg[15][37]  ( .D(n6051), .CK(CLK), .QN(n13630) );
  DFF_X1 \REGISTERS_reg[15][36]  ( .D(n6050), .CK(CLK), .QN(n13631) );
  DFF_X1 \REGISTERS_reg[15][35]  ( .D(n6049), .CK(CLK), .QN(n13632) );
  DFF_X1 \REGISTERS_reg[15][34]  ( .D(n6048), .CK(CLK), .QN(n13633) );
  DFF_X1 \REGISTERS_reg[15][33]  ( .D(n6047), .CK(CLK), .QN(n13634) );
  DFF_X1 \REGISTERS_reg[15][32]  ( .D(n6046), .CK(CLK), .QN(n13635) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n6045), .CK(CLK), .QN(n13636) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n6044), .CK(CLK), .QN(n13637) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n6043), .CK(CLK), .QN(n13638) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n6042), .CK(CLK), .QN(n13639) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n6041), .CK(CLK), .QN(n13640) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n6040), .CK(CLK), .QN(n13641) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n6039), .CK(CLK), .QN(n13642) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n6038), .CK(CLK), .QN(n13643) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n6037), .CK(CLK), .QN(n13644) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n6036), .CK(CLK), .QN(n13645) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n6030), .CK(CLK), .QN(n13646) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n6017), .CK(CLK), .QN(n13647) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n6016), .CK(CLK), .QN(n13648) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n6015), .CK(CLK), .QN(n13649) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n6014), .CK(CLK), .QN(n13650) );
  DFF_X1 \REGISTERS_reg[18][59]  ( .D(n5881), .CK(CLK), .Q(n4682), .QN(n12128)
         );
  DFF_X1 \REGISTERS_reg[18][58]  ( .D(n5880), .CK(CLK), .Q(n4678), .QN(n12127)
         );
  DFF_X1 \REGISTERS_reg[18][57]  ( .D(n5879), .CK(CLK), .Q(n4676), .QN(n12126)
         );
  DFF_X1 \REGISTERS_reg[18][56]  ( .D(n5878), .CK(CLK), .Q(n4674), .QN(n12125)
         );
  DFF_X1 \REGISTERS_reg[18][55]  ( .D(n5877), .CK(CLK), .Q(n4672), .QN(n12124)
         );
  DFF_X1 \REGISTERS_reg[18][54]  ( .D(n5876), .CK(CLK), .Q(n4670), .QN(n12123)
         );
  DFF_X1 \REGISTERS_reg[18][53]  ( .D(n5875), .CK(CLK), .Q(n4668), .QN(n12122)
         );
  DFF_X1 \REGISTERS_reg[18][52]  ( .D(n5874), .CK(CLK), .Q(n4666), .QN(n12121)
         );
  DFF_X1 \REGISTERS_reg[18][51]  ( .D(n5873), .CK(CLK), .Q(n4664), .QN(n12120)
         );
  DFF_X1 \REGISTERS_reg[18][50]  ( .D(n5872), .CK(CLK), .Q(n4662), .QN(n12119)
         );
  DFF_X1 \REGISTERS_reg[18][49]  ( .D(n5871), .CK(CLK), .Q(n4660), .QN(n12118)
         );
  DFF_X1 \REGISTERS_reg[18][48]  ( .D(n5870), .CK(CLK), .Q(n4658), .QN(n12117)
         );
  DFF_X1 \REGISTERS_reg[18][47]  ( .D(n5869), .CK(CLK), .Q(n4656), .QN(n12116)
         );
  DFF_X1 \REGISTERS_reg[18][46]  ( .D(n5868), .CK(CLK), .Q(n8695), .QN(n12115)
         );
  DFF_X1 \REGISTERS_reg[18][45]  ( .D(n5867), .CK(CLK), .Q(n8693), .QN(n12114)
         );
  DFF_X1 \REGISTERS_reg[18][44]  ( .D(n5866), .CK(CLK), .Q(n8691), .QN(n12113)
         );
  DFF_X1 \REGISTERS_reg[18][43]  ( .D(n5865), .CK(CLK), .Q(n8689), .QN(n12112)
         );
  DFF_X1 \REGISTERS_reg[18][42]  ( .D(n5864), .CK(CLK), .Q(n8687), .QN(n12111)
         );
  DFF_X1 \REGISTERS_reg[18][41]  ( .D(n5863), .CK(CLK), .Q(n8685), .QN(n12110)
         );
  DFF_X1 \REGISTERS_reg[18][40]  ( .D(n5862), .CK(CLK), .Q(n8683), .QN(n12109)
         );
  DFF_X1 \REGISTERS_reg[18][39]  ( .D(n5861), .CK(CLK), .Q(n8681), .QN(n12108)
         );
  DFF_X1 \REGISTERS_reg[18][38]  ( .D(n5860), .CK(CLK), .Q(n8679), .QN(n12107)
         );
  DFF_X1 \REGISTERS_reg[18][37]  ( .D(n5859), .CK(CLK), .Q(n8677), .QN(n12106)
         );
  DFF_X1 \REGISTERS_reg[18][36]  ( .D(n5858), .CK(CLK), .Q(n8675), .QN(n12105)
         );
  DFF_X1 \REGISTERS_reg[18][35]  ( .D(n5857), .CK(CLK), .Q(n8673), .QN(n12104)
         );
  DFF_X1 \REGISTERS_reg[18][34]  ( .D(n5856), .CK(CLK), .Q(n8671), .QN(n12103)
         );
  DFF_X1 \REGISTERS_reg[18][33]  ( .D(n5855), .CK(CLK), .Q(n8669), .QN(n12102)
         );
  DFF_X1 \REGISTERS_reg[18][32]  ( .D(n5854), .CK(CLK), .Q(n8667), .QN(n12101)
         );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n5853), .CK(CLK), .Q(n8665), .QN(n12100)
         );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n5852), .CK(CLK), .Q(n8663), .QN(n12099)
         );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n5851), .CK(CLK), .Q(n8661), .QN(n12098)
         );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n5850), .CK(CLK), .Q(n8659), .QN(n12097)
         );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n5849), .CK(CLK), .Q(n8657), .QN(n12096)
         );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n5848), .CK(CLK), .Q(n8655), .QN(n12095)
         );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n5847), .CK(CLK), .Q(n8653), .QN(n12094)
         );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n5846), .CK(CLK), .Q(n8651), .QN(n12093)
         );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n5845), .CK(CLK), .Q(n8649), .QN(n12045)
         );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n5844), .CK(CLK), .Q(n8647), .QN(n12044)
         );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n5843), .CK(CLK), .Q(n8645), .QN(n12043)
         );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n5842), .CK(CLK), .Q(n8643), .QN(n12042)
         );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n5841), .CK(CLK), .Q(n8641), .QN(n12041)
         );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n5840), .CK(CLK), .Q(n8639), .QN(n12040)
         );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n5839), .CK(CLK), .Q(n8637), .QN(n12039)
         );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n5838), .CK(CLK), .Q(n8635), .QN(n12038)
         );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n5837), .CK(CLK), .Q(n8633), .QN(n12037)
         );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n5836), .CK(CLK), .Q(n8631), .QN(n12036)
         );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n5835), .CK(CLK), .Q(n8629), .QN(n12035)
         );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n5834), .CK(CLK), .Q(n8627), .QN(n12034)
         );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n5833), .CK(CLK), .Q(n8625), .QN(n12033)
         );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n5832), .CK(CLK), .Q(n8623), .QN(n12032)
         );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n5831), .CK(CLK), .Q(n8621), .QN(n12031)
         );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n5830), .CK(CLK), .Q(n8619), .QN(n12030)
         );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n5829), .CK(CLK), .Q(n8617), .QN(n12029)
         );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n5828), .CK(CLK), .Q(n8611), .QN(n12028)
         );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n5827), .CK(CLK), .Q(n8603), .QN(n12027)
         );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n5826), .CK(CLK), .Q(n8599), .QN(n12026)
         );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n5825), .CK(CLK), .Q(n4654), .QN(n12025)
         );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n5824), .CK(CLK), .Q(n4652), .QN(n12024)
         );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n5823), .CK(CLK), .Q(n4646), .QN(n12023)
         );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n5822), .CK(CLK), .Q(n4642), .QN(n12022)
         );
  DFF_X1 \REGISTERS_reg[19][59]  ( .D(n5817), .CK(CLK), .Q(n4683), .QN(n11958)
         );
  DFF_X1 \REGISTERS_reg[19][58]  ( .D(n5816), .CK(CLK), .Q(n4679), .QN(n11957)
         );
  DFF_X1 \REGISTERS_reg[19][57]  ( .D(n5815), .CK(CLK), .Q(n4677), .QN(n11956)
         );
  DFF_X1 \REGISTERS_reg[19][56]  ( .D(n5814), .CK(CLK), .Q(n4675), .QN(n11955)
         );
  DFF_X1 \REGISTERS_reg[19][55]  ( .D(n5813), .CK(CLK), .Q(n4673), .QN(n11954)
         );
  DFF_X1 \REGISTERS_reg[19][54]  ( .D(n5812), .CK(CLK), .Q(n4671), .QN(n11953)
         );
  DFF_X1 \REGISTERS_reg[19][53]  ( .D(n5811), .CK(CLK), .Q(n4669), .QN(n11952)
         );
  DFF_X1 \REGISTERS_reg[19][52]  ( .D(n5810), .CK(CLK), .Q(n4667), .QN(n11951)
         );
  DFF_X1 \REGISTERS_reg[19][51]  ( .D(n5809), .CK(CLK), .Q(n4665), .QN(n11950)
         );
  DFF_X1 \REGISTERS_reg[19][50]  ( .D(n5808), .CK(CLK), .Q(n4663), .QN(n11949)
         );
  DFF_X1 \REGISTERS_reg[19][49]  ( .D(n5807), .CK(CLK), .Q(n4661), .QN(n11948)
         );
  DFF_X1 \REGISTERS_reg[19][48]  ( .D(n5806), .CK(CLK), .Q(n4659), .QN(n11947)
         );
  DFF_X1 \REGISTERS_reg[19][47]  ( .D(n5805), .CK(CLK), .Q(n4657), .QN(n11946)
         );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n5761), .CK(CLK), .Q(n4655), .QN(n11850)
         );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n5760), .CK(CLK), .Q(n4653), .QN(n11849)
         );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n5759), .CK(CLK), .Q(n4647), .QN(n11848)
         );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n5758), .CK(CLK), .Q(n4643), .QN(n11847)
         );
  DFF_X1 \REGISTERS_reg[22][59]  ( .D(n5625), .CK(CLK), .Q(n4684), .QN(n12092)
         );
  DFF_X1 \REGISTERS_reg[22][58]  ( .D(n5624), .CK(CLK), .Q(n4502), .QN(n12091)
         );
  DFF_X1 \REGISTERS_reg[22][57]  ( .D(n5623), .CK(CLK), .Q(n4500), .QN(n12090)
         );
  DFF_X1 \REGISTERS_reg[22][56]  ( .D(n5622), .CK(CLK), .Q(n4498), .QN(n12089)
         );
  DFF_X1 \REGISTERS_reg[22][55]  ( .D(n5621), .CK(CLK), .Q(n4496), .QN(n12088)
         );
  DFF_X1 \REGISTERS_reg[22][54]  ( .D(n5620), .CK(CLK), .Q(n4494), .QN(n12087)
         );
  DFF_X1 \REGISTERS_reg[22][53]  ( .D(n5619), .CK(CLK), .Q(n4492), .QN(n12086)
         );
  DFF_X1 \REGISTERS_reg[22][52]  ( .D(n5618), .CK(CLK), .Q(n4490), .QN(n12085)
         );
  DFF_X1 \REGISTERS_reg[22][51]  ( .D(n5617), .CK(CLK), .Q(n4488), .QN(n12084)
         );
  DFF_X1 \REGISTERS_reg[22][50]  ( .D(n5616), .CK(CLK), .Q(n4486), .QN(n12083)
         );
  DFF_X1 \REGISTERS_reg[22][49]  ( .D(n5615), .CK(CLK), .Q(n7322), .QN(n12082)
         );
  DFF_X1 \REGISTERS_reg[22][48]  ( .D(n5614), .CK(CLK), .Q(n7318), .QN(n12081)
         );
  DFF_X1 \REGISTERS_reg[22][47]  ( .D(n5613), .CK(CLK), .Q(n7314), .QN(n12080)
         );
  DFF_X1 \REGISTERS_reg[22][46]  ( .D(n5612), .CK(CLK), .Q(n7310), .QN(n12079)
         );
  DFF_X1 \REGISTERS_reg[22][45]  ( .D(n5611), .CK(CLK), .Q(n7306), .QN(n12078)
         );
  DFF_X1 \REGISTERS_reg[22][44]  ( .D(n5610), .CK(CLK), .Q(n7302), .QN(n12077)
         );
  DFF_X1 \REGISTERS_reg[22][43]  ( .D(n5609), .CK(CLK), .Q(n7298), .QN(n12076)
         );
  DFF_X1 \REGISTERS_reg[22][42]  ( .D(n5608), .CK(CLK), .Q(n7294), .QN(n12075)
         );
  DFF_X1 \REGISTERS_reg[22][41]  ( .D(n5607), .CK(CLK), .Q(n7290), .QN(n12074)
         );
  DFF_X1 \REGISTERS_reg[22][40]  ( .D(n5606), .CK(CLK), .Q(n7286), .QN(n12073)
         );
  DFF_X1 \REGISTERS_reg[22][39]  ( .D(n5605), .CK(CLK), .Q(n7282), .QN(n12072)
         );
  DFF_X1 \REGISTERS_reg[22][38]  ( .D(n5604), .CK(CLK), .Q(n7278), .QN(n12071)
         );
  DFF_X1 \REGISTERS_reg[22][37]  ( .D(n5603), .CK(CLK), .Q(n7245), .QN(n12070)
         );
  DFF_X1 \REGISTERS_reg[22][36]  ( .D(n5602), .CK(CLK), .Q(n7232), .QN(n12069)
         );
  DFF_X1 \REGISTERS_reg[22][35]  ( .D(n5601), .CK(CLK), .Q(n7229), .QN(n12068)
         );
  DFF_X1 \REGISTERS_reg[22][34]  ( .D(n5600), .CK(CLK), .Q(n7226), .QN(n12067)
         );
  DFF_X1 \REGISTERS_reg[22][33]  ( .D(n5599), .CK(CLK), .Q(n7223), .QN(n12066)
         );
  DFF_X1 \REGISTERS_reg[22][32]  ( .D(n5598), .CK(CLK), .Q(n7220), .QN(n12065)
         );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n5597), .CK(CLK), .Q(n7217), .QN(n12064)
         );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n5596), .CK(CLK), .Q(n7214), .QN(n12063)
         );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n5595), .CK(CLK), .Q(n7211), .QN(n12062)
         );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n5594), .CK(CLK), .Q(n7208), .QN(n12061)
         );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n5593), .CK(CLK), .Q(n7205), .QN(n12060)
         );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n5592), .CK(CLK), .Q(n7202), .QN(n12059)
         );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n5591), .CK(CLK), .Q(n7198), .QN(n12058)
         );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n5590), .CK(CLK), .Q(n7194), .QN(n12057)
         );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n5589), .CK(CLK), .Q(n7190), .QN(n12021)
         );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n5588), .CK(CLK), .Q(n7186), .QN(n12020)
         );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n5587), .CK(CLK), .Q(n7182), .QN(n12019)
         );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n5586), .CK(CLK), .Q(n7178), .QN(n12018)
         );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n5585), .CK(CLK), .Q(n7174), .QN(n12017)
         );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n5584), .CK(CLK), .Q(n7170), .QN(n12016)
         );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n5583), .CK(CLK), .Q(n7166), .QN(n12015)
         );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n5582), .CK(CLK), .Q(n7162), .QN(n12014)
         );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n5581), .CK(CLK), .Q(n7158), .QN(n12013)
         );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n5580), .CK(CLK), .Q(n7154), .QN(n12012)
         );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n5579), .CK(CLK), .Q(n7130), .QN(n12011)
         );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n5578), .CK(CLK), .Q(n7104), .QN(n12010)
         );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n5577), .CK(CLK), .Q(n7100), .QN(n12009)
         );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n5576), .CK(CLK), .Q(n7096), .QN(n12008)
         );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n5575), .CK(CLK), .Q(n7092), .QN(n12007)
         );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n5574), .CK(CLK), .Q(n7088), .QN(n12006)
         );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n5573), .CK(CLK), .Q(n7084), .QN(n12005)
         );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n5572), .CK(CLK), .Q(n8613), .QN(n12004)
         );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n5571), .CK(CLK), .Q(n8605), .QN(n12003)
         );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n5570), .CK(CLK), .Q(n7080), .QN(n12002)
         );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n5569), .CK(CLK), .Q(n4484), .QN(n12001)
         );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n5568), .CK(CLK), .Q(n4482), .QN(n12000)
         );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n5567), .CK(CLK), .Q(n4648), .QN(n11999)
         );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n5566), .CK(CLK), .Q(n4480), .QN(n11998)
         );
  DFF_X1 \REGISTERS_reg[23][59]  ( .D(n5561), .CK(CLK), .Q(n4685), .QN(n11945)
         );
  DFF_X1 \REGISTERS_reg[23][58]  ( .D(n5560), .CK(CLK), .Q(n4503), .QN(n11944)
         );
  DFF_X1 \REGISTERS_reg[23][57]  ( .D(n5559), .CK(CLK), .Q(n4501), .QN(n11943)
         );
  DFF_X1 \REGISTERS_reg[23][56]  ( .D(n5558), .CK(CLK), .Q(n4499), .QN(n11942)
         );
  DFF_X1 \REGISTERS_reg[23][55]  ( .D(n5557), .CK(CLK), .Q(n4497), .QN(n11941)
         );
  DFF_X1 \REGISTERS_reg[23][54]  ( .D(n5556), .CK(CLK), .Q(n4495), .QN(n11940)
         );
  DFF_X1 \REGISTERS_reg[23][53]  ( .D(n5555), .CK(CLK), .Q(n4493), .QN(n11939)
         );
  DFF_X1 \REGISTERS_reg[23][52]  ( .D(n5554), .CK(CLK), .Q(n4491), .QN(n11938)
         );
  DFF_X1 \REGISTERS_reg[23][51]  ( .D(n5553), .CK(CLK), .Q(n4489), .QN(n11937)
         );
  DFF_X1 \REGISTERS_reg[23][50]  ( .D(n5552), .CK(CLK), .Q(n4487), .QN(n11936)
         );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n5505), .CK(CLK), .Q(n4485), .QN(n11846)
         );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n5504), .CK(CLK), .Q(n4483), .QN(n11845)
         );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n5503), .CK(CLK), .Q(n4649), .QN(n11844)
         );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n5502), .CK(CLK), .Q(n4481), .QN(n11843)
         );
  DFF_X1 \REGISTERS_reg[24][59]  ( .D(n5497), .CK(CLK), .QN(n13671) );
  DFF_X1 \REGISTERS_reg[24][58]  ( .D(n5496), .CK(CLK), .QN(n13672) );
  DFF_X1 \REGISTERS_reg[24][57]  ( .D(n5495), .CK(CLK), .QN(n13673) );
  DFF_X1 \REGISTERS_reg[24][56]  ( .D(n5494), .CK(CLK), .QN(n13674) );
  DFF_X1 \REGISTERS_reg[24][55]  ( .D(n5493), .CK(CLK), .QN(n13675) );
  DFF_X1 \REGISTERS_reg[24][54]  ( .D(n5492), .CK(CLK), .QN(n13676) );
  DFF_X1 \REGISTERS_reg[24][53]  ( .D(n5491), .CK(CLK), .QN(n13677) );
  DFF_X1 \REGISTERS_reg[24][52]  ( .D(n5490), .CK(CLK), .QN(n13678) );
  DFF_X1 \REGISTERS_reg[24][51]  ( .D(n5489), .CK(CLK), .QN(n13679) );
  DFF_X1 \REGISTERS_reg[24][50]  ( .D(n5488), .CK(CLK), .QN(n13680) );
  DFF_X1 \REGISTERS_reg[24][49]  ( .D(n5487), .CK(CLK), .QN(n13681) );
  DFF_X1 \REGISTERS_reg[24][48]  ( .D(n5486), .CK(CLK), .QN(n13682) );
  DFF_X1 \REGISTERS_reg[24][47]  ( .D(n5485), .CK(CLK), .QN(n13683) );
  DFF_X1 \REGISTERS_reg[24][46]  ( .D(n5484), .CK(CLK), .QN(n13684) );
  DFF_X1 \REGISTERS_reg[24][45]  ( .D(n5483), .CK(CLK), .QN(n13685) );
  DFF_X1 \REGISTERS_reg[24][44]  ( .D(n5482), .CK(CLK), .QN(n13686) );
  DFF_X1 \REGISTERS_reg[24][43]  ( .D(n5481), .CK(CLK), .QN(n13687) );
  DFF_X1 \REGISTERS_reg[24][42]  ( .D(n5480), .CK(CLK), .QN(n13688) );
  DFF_X1 \REGISTERS_reg[24][41]  ( .D(n5479), .CK(CLK), .QN(n13689) );
  DFF_X1 \REGISTERS_reg[24][40]  ( .D(n5478), .CK(CLK), .QN(n13690) );
  DFF_X1 \REGISTERS_reg[24][39]  ( .D(n5477), .CK(CLK), .QN(n13691) );
  DFF_X1 \REGISTERS_reg[24][38]  ( .D(n5476), .CK(CLK), .QN(n13692) );
  DFF_X1 \REGISTERS_reg[24][37]  ( .D(n5475), .CK(CLK), .QN(n13693) );
  DFF_X1 \REGISTERS_reg[24][36]  ( .D(n5474), .CK(CLK), .QN(n13694) );
  DFF_X1 \REGISTERS_reg[24][35]  ( .D(n5473), .CK(CLK), .QN(n13695) );
  DFF_X1 \REGISTERS_reg[24][34]  ( .D(n5472), .CK(CLK), .QN(n13696) );
  DFF_X1 \REGISTERS_reg[24][33]  ( .D(n5471), .CK(CLK), .QN(n13697) );
  DFF_X1 \REGISTERS_reg[24][32]  ( .D(n5470), .CK(CLK), .QN(n13698) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n5469), .CK(CLK), .QN(n13699) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n5468), .CK(CLK), .QN(n13700) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n5467), .CK(CLK), .QN(n13701) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n5466), .CK(CLK), .QN(n13702) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n5465), .CK(CLK), .QN(n13703) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n5464), .CK(CLK), .QN(n13704) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n5463), .CK(CLK), .QN(n13705) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n5462), .CK(CLK), .QN(n13706) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n5461), .CK(CLK), .QN(n13707) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n5460), .CK(CLK), .QN(n13708) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n5459), .CK(CLK), .QN(n13709) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n5458), .CK(CLK), .QN(n13710) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n5457), .CK(CLK), .QN(n13711) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n5456), .CK(CLK), .QN(n13712) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n5455), .CK(CLK), .QN(n13713) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n5454), .CK(CLK), .QN(n13714) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n5453), .CK(CLK), .QN(n13715) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n5452), .CK(CLK), .QN(n13716) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n5451), .CK(CLK), .QN(n13717) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n5450), .CK(CLK), .QN(n13718) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n5449), .CK(CLK), .QN(n13719) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n5448), .CK(CLK), .QN(n13720) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n5447), .CK(CLK), .QN(n13721) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n5446), .CK(CLK), .QN(n13722) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n5445), .CK(CLK), .QN(n13723) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n5444), .CK(CLK), .QN(n13724) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n5443), .CK(CLK), .QN(n13725) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n5442), .CK(CLK), .QN(n13726) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n5441), .CK(CLK), .QN(n13727) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n5440), .CK(CLK), .QN(n13728) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n5439), .CK(CLK), .QN(n13729) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n5438), .CK(CLK), .QN(n13730) );
  DFF_X1 \REGISTERS_reg[25][59]  ( .D(n5433), .CK(CLK), .QN(n13735) );
  DFF_X1 \REGISTERS_reg[25][58]  ( .D(n5432), .CK(CLK), .QN(n13736) );
  DFF_X1 \REGISTERS_reg[25][57]  ( .D(n5431), .CK(CLK), .QN(n13737) );
  DFF_X1 \REGISTERS_reg[25][56]  ( .D(n5430), .CK(CLK), .QN(n13738) );
  DFF_X1 \REGISTERS_reg[25][55]  ( .D(n5429), .CK(CLK), .QN(n13739) );
  DFF_X1 \REGISTERS_reg[25][54]  ( .D(n5428), .CK(CLK), .QN(n13740) );
  DFF_X1 \REGISTERS_reg[25][53]  ( .D(n5427), .CK(CLK), .QN(n13741) );
  DFF_X1 \REGISTERS_reg[25][52]  ( .D(n5426), .CK(CLK), .QN(n13742) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n5377), .CK(CLK), .QN(n13743) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n5376), .CK(CLK), .QN(n13744) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n5375), .CK(CLK), .QN(n13745) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n5374), .CK(CLK), .QN(n13746) );
  DFF_X1 \REGISTERS_reg[28][59]  ( .D(n5241), .CK(CLK), .QN(n13751) );
  DFF_X1 \REGISTERS_reg[28][58]  ( .D(n5240), .CK(CLK), .QN(n13752) );
  DFF_X1 \REGISTERS_reg[28][57]  ( .D(n5239), .CK(CLK), .QN(n13753) );
  DFF_X1 \REGISTERS_reg[28][56]  ( .D(n5238), .CK(CLK), .QN(n13754) );
  DFF_X1 \REGISTERS_reg[28][55]  ( .D(n5237), .CK(CLK), .QN(n13755) );
  DFF_X1 \REGISTERS_reg[28][54]  ( .D(n5236), .CK(CLK), .QN(n13756) );
  DFF_X1 \REGISTERS_reg[28][53]  ( .D(n5235), .CK(CLK), .QN(n13757) );
  DFF_X1 \REGISTERS_reg[28][52]  ( .D(n5234), .CK(CLK), .QN(n13758) );
  DFF_X1 \REGISTERS_reg[28][51]  ( .D(n5233), .CK(CLK), .QN(n13759) );
  DFF_X1 \REGISTERS_reg[28][50]  ( .D(n5232), .CK(CLK), .QN(n13760) );
  DFF_X1 \REGISTERS_reg[28][49]  ( .D(n5231), .CK(CLK), .QN(n13761) );
  DFF_X1 \REGISTERS_reg[28][48]  ( .D(n5230), .CK(CLK), .QN(n13762) );
  DFF_X1 \REGISTERS_reg[28][47]  ( .D(n5229), .CK(CLK), .QN(n13763) );
  DFF_X1 \REGISTERS_reg[28][46]  ( .D(n5228), .CK(CLK), .QN(n13764) );
  DFF_X1 \REGISTERS_reg[28][45]  ( .D(n5227), .CK(CLK), .QN(n13765) );
  DFF_X1 \REGISTERS_reg[28][44]  ( .D(n5226), .CK(CLK), .QN(n13766) );
  DFF_X1 \REGISTERS_reg[28][43]  ( .D(n5225), .CK(CLK), .QN(n13767) );
  DFF_X1 \REGISTERS_reg[28][42]  ( .D(n5224), .CK(CLK), .QN(n13768) );
  DFF_X1 \REGISTERS_reg[28][41]  ( .D(n5223), .CK(CLK), .QN(n13769) );
  DFF_X1 \REGISTERS_reg[28][40]  ( .D(n5222), .CK(CLK), .QN(n13770) );
  DFF_X1 \REGISTERS_reg[28][39]  ( .D(n5221), .CK(CLK), .QN(n13771) );
  DFF_X1 \REGISTERS_reg[28][38]  ( .D(n5220), .CK(CLK), .QN(n13772) );
  DFF_X1 \REGISTERS_reg[28][37]  ( .D(n5219), .CK(CLK), .QN(n13773) );
  DFF_X1 \REGISTERS_reg[28][36]  ( .D(n5218), .CK(CLK), .QN(n13774) );
  DFF_X1 \REGISTERS_reg[28][35]  ( .D(n5217), .CK(CLK), .QN(n13775) );
  DFF_X1 \REGISTERS_reg[28][34]  ( .D(n5216), .CK(CLK), .QN(n13776) );
  DFF_X1 \REGISTERS_reg[28][33]  ( .D(n5215), .CK(CLK), .QN(n13777) );
  DFF_X1 \REGISTERS_reg[28][32]  ( .D(n5214), .CK(CLK), .QN(n13778) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n5213), .CK(CLK), .QN(n13779) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n5212), .CK(CLK), .QN(n13780) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n5211), .CK(CLK), .QN(n13781) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n5210), .CK(CLK), .QN(n13782) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n5209), .CK(CLK), .QN(n13783) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n5208), .CK(CLK), .QN(n13784) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n5207), .CK(CLK), .QN(n13785) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n5206), .CK(CLK), .QN(n13786) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n5205), .CK(CLK), .QN(n13787) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n5204), .CK(CLK), .QN(n13788) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n5203), .CK(CLK), .QN(n13789) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n5202), .CK(CLK), .QN(n13790) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n5201), .CK(CLK), .QN(n13791) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n5200), .CK(CLK), .QN(n13792) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n5199), .CK(CLK), .QN(n13793) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n5198), .CK(CLK), .QN(n13794) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n5197), .CK(CLK), .QN(n13795) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n5196), .CK(CLK), .QN(n13796) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n5195), .CK(CLK), .QN(n13797) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n5194), .CK(CLK), .QN(n13798) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n5193), .CK(CLK), .QN(n13799) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n5192), .CK(CLK), .QN(n13800) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n5191), .CK(CLK), .QN(n13801) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n5190), .CK(CLK), .QN(n13802) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n5189), .CK(CLK), .QN(n13803) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n5188), .CK(CLK), .QN(n13804) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n5187), .CK(CLK), .QN(n13805) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n5186), .CK(CLK), .QN(n13806) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n5185), .CK(CLK), .QN(n13807) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n5184), .CK(CLK), .QN(n13808) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n5183), .CK(CLK), .QN(n13809) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n5182), .CK(CLK), .QN(n13810) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n5122), .CK(CLK), .QN(n13811) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n5121), .CK(CLK), .QN(n13812) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n5120), .CK(CLK), .QN(n13813) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n5119), .CK(CLK), .QN(n13814) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n5118), .CK(CLK), .QN(n13815) );
  DFF_X1 \OUT1_reg[63]  ( .D(n4989), .CK(CLK), .Q(OUT1[63]), .QN(n4765) );
  DFF_X1 \OUT1_reg[62]  ( .D(n4988), .CK(CLK), .Q(OUT1[62]), .QN(n4766) );
  DFF_X1 \OUT1_reg[61]  ( .D(n4987), .CK(CLK), .Q(OUT1[61]), .QN(n4767) );
  DFF_X1 \OUT1_reg[60]  ( .D(n4986), .CK(CLK), .Q(OUT1[60]), .QN(n4768) );
  DFF_X1 \OUT1_reg[59]  ( .D(n4985), .CK(CLK), .Q(OUT1[59]), .QN(n4769) );
  DFF_X1 \OUT1_reg[58]  ( .D(n4984), .CK(CLK), .Q(OUT1[58]), .QN(n4770) );
  DFF_X1 \OUT1_reg[57]  ( .D(n4983), .CK(CLK), .Q(OUT1[57]), .QN(n4771) );
  DFF_X1 \OUT1_reg[56]  ( .D(n4982), .CK(CLK), .Q(OUT1[56]), .QN(n4772) );
  DFF_X1 \OUT1_reg[55]  ( .D(n4981), .CK(CLK), .Q(OUT1[55]), .QN(n4773) );
  DFF_X1 \OUT1_reg[54]  ( .D(n4980), .CK(CLK), .Q(OUT1[54]), .QN(n4774) );
  DFF_X1 \OUT1_reg[53]  ( .D(n4979), .CK(CLK), .Q(OUT1[53]), .QN(n4775) );
  DFF_X1 \OUT1_reg[52]  ( .D(n4978), .CK(CLK), .Q(OUT1[52]), .QN(n4776) );
  DFF_X1 \OUT1_reg[51]  ( .D(n4977), .CK(CLK), .Q(OUT1[51]), .QN(n4777) );
  DFF_X1 \OUT1_reg[50]  ( .D(n4976), .CK(CLK), .Q(OUT1[50]), .QN(n4778) );
  DFF_X1 \OUT1_reg[49]  ( .D(n4975), .CK(CLK), .Q(OUT1[49]), .QN(n4779) );
  DFF_X1 \OUT1_reg[48]  ( .D(n4974), .CK(CLK), .Q(OUT1[48]), .QN(n4780) );
  DFF_X1 \OUT1_reg[47]  ( .D(n4973), .CK(CLK), .Q(OUT1[47]), .QN(n4781) );
  DFF_X1 \OUT1_reg[46]  ( .D(n4972), .CK(CLK), .Q(OUT1[46]), .QN(n4782) );
  DFF_X1 \OUT1_reg[45]  ( .D(n4971), .CK(CLK), .Q(OUT1[45]), .QN(n4783) );
  DFF_X1 \OUT1_reg[44]  ( .D(n4970), .CK(CLK), .Q(OUT1[44]), .QN(n4784) );
  DFF_X1 \OUT1_reg[43]  ( .D(n4969), .CK(CLK), .Q(OUT1[43]), .QN(n4785) );
  DFF_X1 \OUT1_reg[42]  ( .D(n4968), .CK(CLK), .Q(OUT1[42]), .QN(n4786) );
  DFF_X1 \OUT1_reg[41]  ( .D(n4967), .CK(CLK), .Q(OUT1[41]), .QN(n4787) );
  DFF_X1 \OUT1_reg[40]  ( .D(n4966), .CK(CLK), .Q(OUT1[40]), .QN(n4788) );
  DFF_X1 \OUT1_reg[39]  ( .D(n4965), .CK(CLK), .Q(OUT1[39]), .QN(n4789) );
  DFF_X1 \OUT1_reg[38]  ( .D(n4964), .CK(CLK), .Q(OUT1[38]), .QN(n4790) );
  DFF_X1 \OUT1_reg[37]  ( .D(n4963), .CK(CLK), .Q(OUT1[37]), .QN(n4791) );
  DFF_X1 \OUT1_reg[36]  ( .D(n4962), .CK(CLK), .Q(OUT1[36]), .QN(n4792) );
  DFF_X1 \OUT1_reg[35]  ( .D(n4961), .CK(CLK), .Q(OUT1[35]), .QN(n4793) );
  DFF_X1 \OUT1_reg[34]  ( .D(n4960), .CK(CLK), .Q(OUT1[34]), .QN(n4794) );
  DFF_X1 \OUT1_reg[33]  ( .D(n4959), .CK(CLK), .Q(OUT1[33]), .QN(n4795) );
  DFF_X1 \OUT1_reg[32]  ( .D(n4958), .CK(CLK), .Q(OUT1[32]), .QN(n4796) );
  DFF_X1 \OUT1_reg[31]  ( .D(n4957), .CK(CLK), .Q(OUT1[31]), .QN(n4797) );
  DFF_X1 \OUT1_reg[30]  ( .D(n4956), .CK(CLK), .Q(OUT1[30]), .QN(n4803) );
  DFF_X1 \OUT1_reg[29]  ( .D(n4955), .CK(CLK), .Q(OUT1[29]), .QN(n4804) );
  DFF_X1 \OUT1_reg[28]  ( .D(n4954), .CK(CLK), .Q(OUT1[28]), .QN(n4805) );
  DFF_X1 \OUT1_reg[27]  ( .D(n4953), .CK(CLK), .Q(OUT1[27]), .QN(n4806) );
  DFF_X1 \OUT1_reg[26]  ( .D(n4952), .CK(CLK), .Q(OUT1[26]), .QN(n4807) );
  DFF_X1 \OUT1_reg[25]  ( .D(n4951), .CK(CLK), .Q(OUT1[25]), .QN(n4808) );
  DFF_X1 \OUT1_reg[24]  ( .D(n4950), .CK(CLK), .Q(OUT1[24]), .QN(n4809) );
  DFF_X1 \OUT1_reg[23]  ( .D(n4949), .CK(CLK), .Q(OUT1[23]), .QN(n4810) );
  DFF_X1 \OUT1_reg[22]  ( .D(n4948), .CK(CLK), .Q(OUT1[22]), .QN(n4811) );
  DFF_X1 \OUT1_reg[21]  ( .D(n4947), .CK(CLK), .Q(OUT1[21]), .QN(n4812) );
  DFF_X1 \OUT1_reg[20]  ( .D(n4946), .CK(CLK), .Q(OUT1[20]), .QN(n4813) );
  DFF_X1 \OUT1_reg[19]  ( .D(n4945), .CK(CLK), .Q(OUT1[19]), .QN(n4814) );
  DFF_X1 \OUT1_reg[18]  ( .D(n4944), .CK(CLK), .Q(OUT1[18]), .QN(n4815) );
  DFF_X1 \OUT1_reg[17]  ( .D(n4943), .CK(CLK), .Q(OUT1[17]), .QN(n4816) );
  DFF_X1 \OUT1_reg[16]  ( .D(n4942), .CK(CLK), .Q(OUT1[16]), .QN(n4817) );
  DFF_X1 \OUT1_reg[15]  ( .D(n4941), .CK(CLK), .Q(OUT1[15]), .QN(n4818) );
  DFF_X1 \OUT1_reg[14]  ( .D(n4940), .CK(CLK), .Q(OUT1[14]), .QN(n4819) );
  DFF_X1 \OUT1_reg[13]  ( .D(n4939), .CK(CLK), .Q(OUT1[13]), .QN(n4820) );
  DFF_X1 \OUT1_reg[12]  ( .D(n4938), .CK(CLK), .Q(OUT1[12]), .QN(n4821) );
  DFF_X1 \OUT1_reg[11]  ( .D(n4937), .CK(CLK), .Q(OUT1[11]), .QN(n4822) );
  DFF_X1 \OUT1_reg[10]  ( .D(n4936), .CK(CLK), .Q(OUT1[10]), .QN(n4823) );
  DFF_X1 \OUT1_reg[9]  ( .D(n4935), .CK(CLK), .Q(OUT1[9]), .QN(n4824) );
  DFF_X1 \OUT1_reg[8]  ( .D(n4934), .CK(CLK), .Q(OUT1[8]), .QN(n4825) );
  DFF_X1 \OUT1_reg[7]  ( .D(n4933), .CK(CLK), .Q(OUT1[7]), .QN(n4826) );
  DFF_X1 \OUT1_reg[6]  ( .D(n4932), .CK(CLK), .Q(OUT1[6]), .QN(n4827) );
  DFF_X1 \OUT1_reg[5]  ( .D(n4931), .CK(CLK), .Q(OUT1[5]), .QN(n4828) );
  DFF_X1 \OUT1_reg[4]  ( .D(n4930), .CK(CLK), .Q(OUT1[4]), .QN(n4829) );
  DFF_X1 \OUT1_reg[3]  ( .D(n4929), .CK(CLK), .Q(OUT1[3]), .QN(n4830) );
  DFF_X1 \OUT1_reg[2]  ( .D(n4928), .CK(CLK), .Q(OUT1[2]), .QN(n4831) );
  DFF_X1 \OUT1_reg[1]  ( .D(n4927), .CK(CLK), .Q(OUT1[1]), .QN(n4832) );
  DFF_X1 \OUT1_reg[0]  ( .D(n4926), .CK(CLK), .Q(OUT1[0]), .QN(n4833) );
  DFF_X1 \OUT2_reg[63]  ( .D(n4925), .CK(CLK), .Q(OUT2[63]), .QN(n4834) );
  DFF_X1 \OUT2_reg[62]  ( .D(n4924), .CK(CLK), .Q(OUT2[62]), .QN(n4851) );
  DFF_X1 \OUT2_reg[61]  ( .D(n4923), .CK(CLK), .Q(OUT2[61]), .QN(n7112) );
  DFF_X1 \OUT2_reg[60]  ( .D(n4922), .CK(CLK), .Q(OUT2[60]), .QN(n7129) );
  DFF_X1 \OUT2_reg[59]  ( .D(n4921), .CK(CLK), .Q(OUT2[59]), .QN(n7146) );
  DFF_X1 \OUT2_reg[58]  ( .D(n4920), .CK(CLK), .Q(OUT2[58]), .QN(n7243) );
  DFF_X1 \OUT2_reg[57]  ( .D(n4919), .CK(CLK), .Q(OUT2[57]), .QN(n7260) );
  DFF_X1 \OUT2_reg[56]  ( .D(n4918), .CK(CLK), .Q(OUT2[56]), .QN(n7277) );
  DFF_X1 \OUT2_reg[55]  ( .D(n4917), .CK(CLK), .Q(OUT2[55]), .QN(n7376) );
  DFF_X1 \OUT2_reg[54]  ( .D(n4916), .CK(CLK), .Q(OUT2[54]), .QN(n7393) );
  DFF_X1 \OUT2_reg[53]  ( .D(n4915), .CK(CLK), .Q(OUT2[53]), .QN(n7495) );
  DFF_X1 \OUT2_reg[52]  ( .D(n4914), .CK(CLK), .Q(OUT2[52]), .QN(n7512) );
  DFF_X1 \OUT2_reg[51]  ( .D(n4913), .CK(CLK), .Q(OUT2[51]), .QN(n7529) );
  DFF_X1 \OUT2_reg[50]  ( .D(n4912), .CK(CLK), .Q(OUT2[50]), .QN(n7633) );
  DFF_X1 \OUT2_reg[49]  ( .D(n4911), .CK(CLK), .Q(OUT2[49]), .QN(n7650) );
  DFF_X1 \OUT2_reg[48]  ( .D(n4910), .CK(CLK), .Q(OUT2[48]), .QN(n7752) );
  DFF_X1 \OUT2_reg[47]  ( .D(n4909), .CK(CLK), .Q(OUT2[47]), .QN(n7769) );
  DFF_X1 \OUT2_reg[46]  ( .D(n4908), .CK(CLK), .Q(OUT2[46]), .QN(n7786) );
  DFF_X1 \OUT2_reg[45]  ( .D(n4907), .CK(CLK), .Q(OUT2[45]), .QN(n7803) );
  DFF_X1 \OUT2_reg[44]  ( .D(n4906), .CK(CLK), .Q(OUT2[44]), .QN(n7820) );
  DFF_X1 \OUT2_reg[43]  ( .D(n4905), .CK(CLK), .Q(OUT2[43]), .QN(n7837) );
  DFF_X1 \OUT2_reg[42]  ( .D(n4904), .CK(CLK), .Q(OUT2[42]), .QN(n7854) );
  DFF_X1 \OUT2_reg[41]  ( .D(n4903), .CK(CLK), .Q(OUT2[41]), .QN(n7871) );
  DFF_X1 \OUT2_reg[40]  ( .D(n4902), .CK(CLK), .Q(OUT2[40]), .QN(n7888) );
  DFF_X1 \OUT2_reg[39]  ( .D(n4901), .CK(CLK), .Q(OUT2[39]), .QN(n7905) );
  DFF_X1 \OUT2_reg[38]  ( .D(n4900), .CK(CLK), .Q(OUT2[38]), .QN(n7922) );
  DFF_X1 \OUT2_reg[37]  ( .D(n4899), .CK(CLK), .Q(OUT2[37]), .QN(n7939) );
  DFF_X1 \OUT2_reg[36]  ( .D(n4898), .CK(CLK), .Q(OUT2[36]), .QN(n7956) );
  DFF_X1 \OUT2_reg[35]  ( .D(n4897), .CK(CLK), .Q(OUT2[35]), .QN(n7973) );
  DFF_X1 \OUT2_reg[34]  ( .D(n4896), .CK(CLK), .Q(OUT2[34]), .QN(n7990) );
  DFF_X1 \OUT2_reg[33]  ( .D(n4895), .CK(CLK), .Q(OUT2[33]), .QN(n8007) );
  DFF_X1 \OUT2_reg[32]  ( .D(n4894), .CK(CLK), .Q(OUT2[32]), .QN(n8024) );
  DFF_X1 \OUT2_reg[31]  ( .D(n4893), .CK(CLK), .Q(OUT2[31]), .QN(n8041) );
  DFF_X1 \OUT2_reg[30]  ( .D(n4892), .CK(CLK), .Q(OUT2[30]), .QN(n8058) );
  DFF_X1 \OUT2_reg[29]  ( .D(n4891), .CK(CLK), .Q(OUT2[29]), .QN(n8075) );
  DFF_X1 \OUT2_reg[28]  ( .D(n4890), .CK(CLK), .Q(OUT2[28]), .QN(n8092) );
  DFF_X1 \OUT2_reg[27]  ( .D(n4889), .CK(CLK), .Q(OUT2[27]), .QN(n8109) );
  DFF_X1 \OUT2_reg[26]  ( .D(n4888), .CK(CLK), .Q(OUT2[26]), .QN(n8126) );
  DFF_X1 \OUT2_reg[25]  ( .D(n4887), .CK(CLK), .Q(OUT2[25]), .QN(n8143) );
  DFF_X1 \OUT2_reg[24]  ( .D(n4886), .CK(CLK), .Q(OUT2[24]), .QN(n8160) );
  DFF_X1 \OUT2_reg[23]  ( .D(n4885), .CK(CLK), .Q(OUT2[23]), .QN(n8177) );
  DFF_X1 \OUT2_reg[22]  ( .D(n4884), .CK(CLK), .Q(OUT2[22]), .QN(n8194) );
  DFF_X1 \OUT2_reg[21]  ( .D(n4883), .CK(CLK), .Q(OUT2[21]), .QN(n8211) );
  DFF_X1 \OUT2_reg[20]  ( .D(n4882), .CK(CLK), .Q(OUT2[20]), .QN(n8228) );
  DFF_X1 \OUT2_reg[19]  ( .D(n4881), .CK(CLK), .Q(OUT2[19]), .QN(n8245) );
  DFF_X1 \OUT2_reg[18]  ( .D(n4880), .CK(CLK), .Q(OUT2[18]), .QN(n8262) );
  DFF_X1 \OUT2_reg[17]  ( .D(n4879), .CK(CLK), .Q(OUT2[17]), .QN(n8279) );
  DFF_X1 \OUT2_reg[16]  ( .D(n4878), .CK(CLK), .Q(OUT2[16]), .QN(n8296) );
  DFF_X1 \OUT2_reg[15]  ( .D(n4877), .CK(CLK), .Q(OUT2[15]), .QN(n8313) );
  DFF_X1 \OUT2_reg[14]  ( .D(n4876), .CK(CLK), .Q(OUT2[14]), .QN(n8330) );
  DFF_X1 \OUT2_reg[13]  ( .D(n4875), .CK(CLK), .Q(OUT2[13]), .QN(n8347) );
  DFF_X1 \OUT2_reg[12]  ( .D(n4874), .CK(CLK), .Q(OUT2[12]), .QN(n8364) );
  DFF_X1 \OUT2_reg[11]  ( .D(n4873), .CK(CLK), .Q(OUT2[11]), .QN(n8381) );
  DFF_X1 \OUT2_reg[10]  ( .D(n4872), .CK(CLK), .Q(OUT2[10]), .QN(n8398) );
  DFF_X1 \OUT2_reg[9]  ( .D(n4871), .CK(CLK), .Q(OUT2[9]), .QN(n8415) );
  DFF_X1 \OUT2_reg[8]  ( .D(n4870), .CK(CLK), .Q(OUT2[8]), .QN(n8432) );
  DFF_X1 \OUT2_reg[7]  ( .D(n4869), .CK(CLK), .Q(OUT2[7]), .QN(n8449) );
  DFF_X1 \OUT2_reg[6]  ( .D(n4868), .CK(CLK), .Q(OUT2[6]), .QN(n8466) );
  DFF_X1 \OUT2_reg[5]  ( .D(n4867), .CK(CLK), .Q(OUT2[5]), .QN(n8483) );
  DFF_X1 \OUT2_reg[4]  ( .D(n4866), .CK(CLK), .Q(OUT2[4]), .QN(n8500) );
  DFF_X1 \OUT2_reg[3]  ( .D(n4865), .CK(CLK), .Q(OUT2[3]), .QN(n8517) );
  DFF_X1 \OUT2_reg[2]  ( .D(n4864), .CK(CLK), .Q(OUT2[2]), .QN(n8534) );
  DFF_X1 \OUT2_reg[1]  ( .D(n4863), .CK(CLK), .Q(OUT2[1]), .QN(n8551) );
  DFF_X1 \OUT2_reg[0]  ( .D(n4862), .CK(CLK), .Q(OUT2[0]), .QN(n8568) );
  DFF_X1 \REGISTERS_reg[3][62]  ( .D(n6844), .CK(CLK), .Q(n9950), .QN(n11997)
         );
  DFF_X1 \REGISTERS_reg[3][61]  ( .D(n6843), .CK(CLK), .Q(n9951), .QN(n11996)
         );
  DFF_X1 \REGISTERS_reg[3][60]  ( .D(n6842), .CK(CLK), .Q(n9952), .QN(n11995)
         );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n5401), .CK(CLK), .QN(n13869) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n5400), .CK(CLK), .QN(n13870) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n5399), .CK(CLK), .QN(n13871) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n5398), .CK(CLK), .QN(n13872) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n5397), .CK(CLK), .QN(n13873) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n5396), .CK(CLK), .QN(n13874) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n5395), .CK(CLK), .QN(n13875) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n5394), .CK(CLK), .QN(n13876) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n5393), .CK(CLK), .QN(n13877) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n5392), .CK(CLK), .QN(n13878) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n5391), .CK(CLK), .QN(n13879) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n5390), .CK(CLK), .QN(n13880) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n5389), .CK(CLK), .QN(n13881) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n5388), .CK(CLK), .QN(n13882) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n5387), .CK(CLK), .QN(n13883) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n5386), .CK(CLK), .QN(n13884) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n5385), .CK(CLK), .QN(n13885) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n5384), .CK(CLK), .QN(n13886) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n5383), .CK(CLK), .QN(n13887) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n5382), .CK(CLK), .QN(n13888) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n5381), .CK(CLK), .QN(n13889) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n5380), .CK(CLK), .QN(n13890) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n5379), .CK(CLK), .QN(n13891) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n5378), .CK(CLK), .QN(n13892) );
  DFF_X1 \REGISTERS_reg[29][39]  ( .D(n5157), .CK(CLK), .QN(n13929) );
  DFF_X1 \REGISTERS_reg[29][38]  ( .D(n5156), .CK(CLK), .QN(n13930) );
  DFF_X1 \REGISTERS_reg[29][37]  ( .D(n5155), .CK(CLK), .QN(n13931) );
  DFF_X1 \REGISTERS_reg[29][36]  ( .D(n5154), .CK(CLK), .QN(n13932) );
  DFF_X1 \REGISTERS_reg[29][35]  ( .D(n5153), .CK(CLK), .QN(n13933) );
  DFF_X1 \REGISTERS_reg[29][34]  ( .D(n5152), .CK(CLK), .QN(n13934) );
  DFF_X1 \REGISTERS_reg[29][33]  ( .D(n5151), .CK(CLK), .QN(n13935) );
  DFF_X1 \REGISTERS_reg[29][32]  ( .D(n5150), .CK(CLK), .QN(n13936) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n5149), .CK(CLK), .QN(n13937) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n5148), .CK(CLK), .QN(n13938) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n5147), .CK(CLK), .QN(n13939) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n5146), .CK(CLK), .QN(n13940) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n5145), .CK(CLK), .QN(n13941) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n5144), .CK(CLK), .QN(n13942) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n5143), .CK(CLK), .QN(n13943) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n5142), .CK(CLK), .QN(n13944) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n5141), .CK(CLK), .QN(n13945) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n5140), .CK(CLK), .QN(n13946) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n5139), .CK(CLK), .QN(n13947) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n5138), .CK(CLK), .QN(n13948) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n5137), .CK(CLK), .QN(n13949) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n5136), .CK(CLK), .QN(n13950) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n5135), .CK(CLK), .QN(n13951) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n5134), .CK(CLK), .QN(n13952) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n5133), .CK(CLK), .QN(n14025) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n5132), .CK(CLK), .QN(n14026) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n5131), .CK(CLK), .QN(n14027) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n5130), .CK(CLK), .QN(n14028) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n5129), .CK(CLK), .QN(n14029) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n5128), .CK(CLK), .QN(n14030) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n5127), .CK(CLK), .QN(n14031) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n5126), .CK(CLK), .QN(n14032) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n5125), .CK(CLK), .QN(n14033) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n5124), .CK(CLK), .QN(n14034) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n5123), .CK(CLK), .QN(n14035) );
  DFF_X1 \REGISTERS_reg[25][51]  ( .D(n5425), .CK(CLK), .QN(n14036) );
  DFF_X1 \REGISTERS_reg[25][50]  ( .D(n5424), .CK(CLK), .QN(n14037) );
  DFF_X1 \REGISTERS_reg[25][49]  ( .D(n5423), .CK(CLK), .QN(n14038) );
  DFF_X1 \REGISTERS_reg[25][48]  ( .D(n5422), .CK(CLK), .QN(n14039) );
  DFF_X1 \REGISTERS_reg[25][47]  ( .D(n5421), .CK(CLK), .QN(n14040) );
  DFF_X1 \REGISTERS_reg[25][46]  ( .D(n5420), .CK(CLK), .QN(n14041) );
  DFF_X1 \REGISTERS_reg[25][45]  ( .D(n5419), .CK(CLK), .QN(n14042) );
  DFF_X1 \REGISTERS_reg[25][44]  ( .D(n5418), .CK(CLK), .QN(n14043) );
  DFF_X1 \REGISTERS_reg[25][43]  ( .D(n5417), .CK(CLK), .QN(n14044) );
  DFF_X1 \REGISTERS_reg[25][42]  ( .D(n5416), .CK(CLK), .QN(n14045) );
  DFF_X1 \REGISTERS_reg[25][41]  ( .D(n5415), .CK(CLK), .QN(n14046) );
  DFF_X1 \REGISTERS_reg[25][40]  ( .D(n5414), .CK(CLK), .QN(n14047) );
  DFF_X1 \REGISTERS_reg[25][39]  ( .D(n5413), .CK(CLK), .QN(n14048) );
  DFF_X1 \REGISTERS_reg[25][38]  ( .D(n5412), .CK(CLK), .QN(n14049) );
  DFF_X1 \REGISTERS_reg[25][37]  ( .D(n5411), .CK(CLK), .QN(n14050) );
  DFF_X1 \REGISTERS_reg[25][36]  ( .D(n5410), .CK(CLK), .QN(n14051) );
  DFF_X1 \REGISTERS_reg[25][35]  ( .D(n5409), .CK(CLK), .QN(n14052) );
  DFF_X1 \REGISTERS_reg[25][34]  ( .D(n5408), .CK(CLK), .QN(n14053) );
  DFF_X1 \REGISTERS_reg[25][33]  ( .D(n5407), .CK(CLK), .QN(n14054) );
  DFF_X1 \REGISTERS_reg[25][32]  ( .D(n5406), .CK(CLK), .QN(n14055) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n5405), .CK(CLK), .QN(n14056) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n5404), .CK(CLK), .QN(n14057) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n5403), .CK(CLK), .QN(n14058) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n5402), .CK(CLK), .QN(n14059) );
  DFF_X1 \REGISTERS_reg[29][59]  ( .D(n5177), .CK(CLK), .QN(n14087) );
  DFF_X1 \REGISTERS_reg[29][58]  ( .D(n5176), .CK(CLK), .QN(n14088) );
  DFF_X1 \REGISTERS_reg[29][57]  ( .D(n5175), .CK(CLK), .QN(n14089) );
  DFF_X1 \REGISTERS_reg[29][56]  ( .D(n5174), .CK(CLK), .QN(n14090) );
  DFF_X1 \REGISTERS_reg[29][55]  ( .D(n5173), .CK(CLK), .QN(n14091) );
  DFF_X1 \REGISTERS_reg[29][54]  ( .D(n5172), .CK(CLK), .QN(n14092) );
  DFF_X1 \REGISTERS_reg[29][53]  ( .D(n5171), .CK(CLK), .QN(n14093) );
  DFF_X1 \REGISTERS_reg[29][52]  ( .D(n5170), .CK(CLK), .QN(n14094) );
  DFF_X1 \REGISTERS_reg[29][51]  ( .D(n5169), .CK(CLK), .QN(n14095) );
  DFF_X1 \REGISTERS_reg[29][50]  ( .D(n5168), .CK(CLK), .QN(n14096) );
  DFF_X1 \REGISTERS_reg[29][49]  ( .D(n5167), .CK(CLK), .QN(n14097) );
  DFF_X1 \REGISTERS_reg[29][48]  ( .D(n5166), .CK(CLK), .QN(n14098) );
  DFF_X1 \REGISTERS_reg[29][47]  ( .D(n5165), .CK(CLK), .QN(n14099) );
  DFF_X1 \REGISTERS_reg[29][46]  ( .D(n5164), .CK(CLK), .QN(n14100) );
  DFF_X1 \REGISTERS_reg[29][45]  ( .D(n5163), .CK(CLK), .QN(n14101) );
  DFF_X1 \REGISTERS_reg[29][44]  ( .D(n5162), .CK(CLK), .QN(n14102) );
  DFF_X1 \REGISTERS_reg[29][43]  ( .D(n5161), .CK(CLK), .QN(n14103) );
  DFF_X1 \REGISTERS_reg[29][42]  ( .D(n5160), .CK(CLK), .QN(n14104) );
  DFF_X1 \REGISTERS_reg[29][41]  ( .D(n5159), .CK(CLK), .QN(n14105) );
  DFF_X1 \REGISTERS_reg[29][40]  ( .D(n5158), .CK(CLK), .QN(n14106) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n5527), .CK(CLK), .Q(n7199), .QN(n11935)
         );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n5526), .CK(CLK), .Q(n7195), .QN(n11934)
         );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n5525), .CK(CLK), .Q(n7191), .QN(n11842)
         );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n5524), .CK(CLK), .Q(n7187), .QN(n11841)
         );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n5523), .CK(CLK), .Q(n7183), .QN(n11840)
         );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n5522), .CK(CLK), .Q(n7179), .QN(n11839)
         );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n5521), .CK(CLK), .Q(n7175), .QN(n11838)
         );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n5520), .CK(CLK), .Q(n7171), .QN(n11837)
         );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n5519), .CK(CLK), .Q(n7167), .QN(n11836)
         );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n5518), .CK(CLK), .Q(n7163), .QN(n11835)
         );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n5517), .CK(CLK), .Q(n7159), .QN(n11834)
         );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n5516), .CK(CLK), .Q(n7155), .QN(n11833)
         );
  DFF_X1 \REGISTERS_reg[21][34]  ( .D(n5664), .CK(CLK), .QN(n8001) );
  DFF_X1 \REGISTERS_reg[21][33]  ( .D(n5663), .CK(CLK), .QN(n8018) );
  DFF_X1 \REGISTERS_reg[21][32]  ( .D(n5662), .CK(CLK), .QN(n8035) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n5661), .CK(CLK), .QN(n8052) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n5660), .CK(CLK), .QN(n8069) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n5659), .CK(CLK), .QN(n8086) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n5658), .CK(CLK), .QN(n8103) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n5657), .CK(CLK), .QN(n8120) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n5656), .CK(CLK), .QN(n8137) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n5655), .CK(CLK), .QN(n8154) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n5654), .CK(CLK), .QN(n8171) );
  DFF_X1 \REGISTERS_reg[20][59]  ( .D(n5753), .CK(CLK), .QN(n7238) );
  DFF_X1 \REGISTERS_reg[20][58]  ( .D(n5752), .CK(CLK), .QN(n7255) );
  DFF_X1 \REGISTERS_reg[20][57]  ( .D(n5751), .CK(CLK), .QN(n7272) );
  DFF_X1 \REGISTERS_reg[20][56]  ( .D(n5750), .CK(CLK), .QN(n7371) );
  DFF_X1 \REGISTERS_reg[20][55]  ( .D(n5749), .CK(CLK), .QN(n7388) );
  DFF_X1 \REGISTERS_reg[20][54]  ( .D(n5748), .CK(CLK), .QN(n7490) );
  DFF_X1 \REGISTERS_reg[20][53]  ( .D(n5747), .CK(CLK), .QN(n7507) );
  DFF_X1 \REGISTERS_reg[20][52]  ( .D(n5746), .CK(CLK), .QN(n7524) );
  DFF_X1 \REGISTERS_reg[20][51]  ( .D(n5745), .CK(CLK), .QN(n7628) );
  DFF_X1 \REGISTERS_reg[20][50]  ( .D(n5744), .CK(CLK), .QN(n7645) );
  DFF_X1 \REGISTERS_reg[20][49]  ( .D(n5743), .CK(CLK), .QN(n7747) );
  DFF_X1 \REGISTERS_reg[20][48]  ( .D(n5742), .CK(CLK), .QN(n7764) );
  DFF_X1 \REGISTERS_reg[20][47]  ( .D(n5741), .CK(CLK), .QN(n7781) );
  DFF_X1 \REGISTERS_reg[20][46]  ( .D(n5740), .CK(CLK), .QN(n7798) );
  DFF_X1 \REGISTERS_reg[20][45]  ( .D(n5739), .CK(CLK), .QN(n7815) );
  DFF_X1 \REGISTERS_reg[20][44]  ( .D(n5738), .CK(CLK), .QN(n7832) );
  DFF_X1 \REGISTERS_reg[20][43]  ( .D(n5737), .CK(CLK), .QN(n7849) );
  DFF_X1 \REGISTERS_reg[20][42]  ( .D(n5736), .CK(CLK), .QN(n7866) );
  DFF_X1 \REGISTERS_reg[20][41]  ( .D(n5735), .CK(CLK), .QN(n7883) );
  DFF_X1 \REGISTERS_reg[20][40]  ( .D(n5734), .CK(CLK), .QN(n7900) );
  DFF_X1 \REGISTERS_reg[20][39]  ( .D(n5733), .CK(CLK), .QN(n7917) );
  DFF_X1 \REGISTERS_reg[20][38]  ( .D(n5732), .CK(CLK), .QN(n7934) );
  DFF_X1 \REGISTERS_reg[20][37]  ( .D(n5731), .CK(CLK), .QN(n7951) );
  DFF_X1 \REGISTERS_reg[20][36]  ( .D(n5730), .CK(CLK), .QN(n7968) );
  DFF_X1 \REGISTERS_reg[20][35]  ( .D(n5729), .CK(CLK), .QN(n7985) );
  DFF_X1 \REGISTERS_reg[20][34]  ( .D(n5728), .CK(CLK), .QN(n8002) );
  DFF_X1 \REGISTERS_reg[20][33]  ( .D(n5727), .CK(CLK), .QN(n8019) );
  DFF_X1 \REGISTERS_reg[20][32]  ( .D(n5726), .CK(CLK), .QN(n8036) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n5725), .CK(CLK), .QN(n8053) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n5724), .CK(CLK), .QN(n8070) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n5723), .CK(CLK), .QN(n8087) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n5722), .CK(CLK), .QN(n8104) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n5721), .CK(CLK), .QN(n8121) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n5720), .CK(CLK), .QN(n8138) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n5719), .CK(CLK), .QN(n8155) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n5718), .CK(CLK), .QN(n8172) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n5781), .CK(CLK), .Q(n8650), .QN(n11832)
         );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n5780), .CK(CLK), .Q(n8648), .QN(n11831)
         );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n5779), .CK(CLK), .Q(n8646), .QN(n11830)
         );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n5778), .CK(CLK), .Q(n8644), .QN(n11829)
         );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n5777), .CK(CLK), .Q(n8642), .QN(n11828)
         );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n5776), .CK(CLK), .Q(n8640), .QN(n11827)
         );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n5775), .CK(CLK), .Q(n8638), .QN(n11826)
         );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n5773), .CK(CLK), .Q(n8634), .QN(n11825)
         );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n5772), .CK(CLK), .Q(n8632), .QN(n11824)
         );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n5771), .CK(CLK), .Q(n8630), .QN(n11823)
         );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n5770), .CK(CLK), .Q(n8628), .QN(n11822)
         );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n5766), .CK(CLK), .Q(n8620), .QN(n11821)
         );
  DFF_X1 \REGISTERS_reg[17][59]  ( .D(n5945), .CK(CLK), .QN(n7235) );
  DFF_X1 \REGISTERS_reg[17][58]  ( .D(n5944), .CK(CLK), .QN(n7252) );
  DFF_X1 \REGISTERS_reg[17][57]  ( .D(n5943), .CK(CLK), .QN(n7269) );
  DFF_X1 \REGISTERS_reg[17][56]  ( .D(n5942), .CK(CLK), .QN(n7368) );
  DFF_X1 \REGISTERS_reg[17][55]  ( .D(n5941), .CK(CLK), .QN(n7385) );
  DFF_X1 \REGISTERS_reg[17][54]  ( .D(n5940), .CK(CLK), .QN(n7402) );
  DFF_X1 \REGISTERS_reg[17][53]  ( .D(n5939), .CK(CLK), .QN(n7504) );
  DFF_X1 \REGISTERS_reg[17][52]  ( .D(n5938), .CK(CLK), .QN(n7521) );
  DFF_X1 \REGISTERS_reg[17][51]  ( .D(n5937), .CK(CLK), .QN(n7625) );
  DFF_X1 \REGISTERS_reg[17][50]  ( .D(n5936), .CK(CLK), .QN(n7642) );
  DFF_X1 \REGISTERS_reg[17][49]  ( .D(n5935), .CK(CLK), .QN(n7744) );
  DFF_X1 \REGISTERS_reg[17][48]  ( .D(n5934), .CK(CLK), .QN(n7761) );
  DFF_X1 \REGISTERS_reg[17][47]  ( .D(n5933), .CK(CLK), .QN(n7778) );
  DFF_X1 \REGISTERS_reg[17][46]  ( .D(n5932), .CK(CLK), .QN(n7795) );
  DFF_X1 \REGISTERS_reg[17][45]  ( .D(n5931), .CK(CLK), .QN(n7812) );
  DFF_X1 \REGISTERS_reg[17][44]  ( .D(n5930), .CK(CLK), .QN(n7829) );
  DFF_X1 \REGISTERS_reg[17][43]  ( .D(n5929), .CK(CLK), .QN(n7846) );
  DFF_X1 \REGISTERS_reg[17][42]  ( .D(n5928), .CK(CLK), .QN(n7863) );
  DFF_X1 \REGISTERS_reg[17][41]  ( .D(n5927), .CK(CLK), .QN(n7880) );
  DFF_X1 \REGISTERS_reg[17][40]  ( .D(n5926), .CK(CLK), .QN(n7897) );
  DFF_X1 \REGISTERS_reg[17][39]  ( .D(n5925), .CK(CLK), .QN(n7914) );
  DFF_X1 \REGISTERS_reg[17][38]  ( .D(n5924), .CK(CLK), .QN(n7931) );
  DFF_X1 \REGISTERS_reg[17][37]  ( .D(n5923), .CK(CLK), .QN(n7948) );
  DFF_X1 \REGISTERS_reg[17][36]  ( .D(n5922), .CK(CLK), .QN(n7965) );
  DFF_X1 \REGISTERS_reg[17][35]  ( .D(n5921), .CK(CLK), .QN(n7982) );
  DFF_X1 \REGISTERS_reg[17][34]  ( .D(n5920), .CK(CLK), .QN(n7999) );
  DFF_X1 \REGISTERS_reg[17][33]  ( .D(n5919), .CK(CLK), .QN(n8016) );
  DFF_X1 \REGISTERS_reg[17][32]  ( .D(n5918), .CK(CLK), .QN(n8033) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n5917), .CK(CLK), .QN(n8050) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n5916), .CK(CLK), .QN(n8067) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n5915), .CK(CLK), .QN(n8084) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n5914), .CK(CLK), .QN(n8101) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n5913), .CK(CLK), .QN(n8118) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n5912), .CK(CLK), .QN(n8135) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n5911), .CK(CLK), .QN(n8152) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n5910), .CK(CLK), .QN(n8169) );
  DFF_X1 \REGISTERS_reg[16][59]  ( .D(n6009), .CK(CLK), .QN(n7236) );
  DFF_X1 \REGISTERS_reg[16][58]  ( .D(n6008), .CK(CLK), .QN(n7253) );
  DFF_X1 \REGISTERS_reg[16][57]  ( .D(n6007), .CK(CLK), .QN(n7270) );
  DFF_X1 \REGISTERS_reg[16][56]  ( .D(n6006), .CK(CLK), .QN(n7369) );
  DFF_X1 \REGISTERS_reg[16][55]  ( .D(n6005), .CK(CLK), .QN(n7386) );
  DFF_X1 \REGISTERS_reg[16][54]  ( .D(n6004), .CK(CLK), .QN(n7403) );
  DFF_X1 \REGISTERS_reg[16][53]  ( .D(n6003), .CK(CLK), .QN(n7505) );
  DFF_X1 \REGISTERS_reg[16][52]  ( .D(n6002), .CK(CLK), .QN(n7522) );
  DFF_X1 \REGISTERS_reg[16][51]  ( .D(n6001), .CK(CLK), .QN(n7626) );
  DFF_X1 \REGISTERS_reg[16][50]  ( .D(n6000), .CK(CLK), .QN(n7643) );
  DFF_X1 \REGISTERS_reg[16][49]  ( .D(n5999), .CK(CLK), .QN(n7745) );
  DFF_X1 \REGISTERS_reg[16][48]  ( .D(n5998), .CK(CLK), .QN(n7762) );
  DFF_X1 \REGISTERS_reg[16][47]  ( .D(n5997), .CK(CLK), .QN(n7779) );
  DFF_X1 \REGISTERS_reg[16][46]  ( .D(n5996), .CK(CLK), .QN(n7796) );
  DFF_X1 \REGISTERS_reg[16][45]  ( .D(n5995), .CK(CLK), .QN(n7813) );
  DFF_X1 \REGISTERS_reg[16][44]  ( .D(n5994), .CK(CLK), .QN(n7830) );
  DFF_X1 \REGISTERS_reg[16][43]  ( .D(n5993), .CK(CLK), .QN(n7847) );
  DFF_X1 \REGISTERS_reg[16][42]  ( .D(n5992), .CK(CLK), .QN(n7864) );
  DFF_X1 \REGISTERS_reg[16][41]  ( .D(n5991), .CK(CLK), .QN(n7881) );
  DFF_X1 \REGISTERS_reg[16][40]  ( .D(n5990), .CK(CLK), .QN(n7898) );
  DFF_X1 \REGISTERS_reg[16][39]  ( .D(n5989), .CK(CLK), .QN(n7915) );
  DFF_X1 \REGISTERS_reg[16][38]  ( .D(n5988), .CK(CLK), .QN(n7932) );
  DFF_X1 \REGISTERS_reg[16][37]  ( .D(n5987), .CK(CLK), .QN(n7949) );
  DFF_X1 \REGISTERS_reg[16][36]  ( .D(n5986), .CK(CLK), .QN(n7966) );
  DFF_X1 \REGISTERS_reg[16][35]  ( .D(n5985), .CK(CLK), .QN(n7983) );
  DFF_X1 \REGISTERS_reg[16][34]  ( .D(n5984), .CK(CLK), .QN(n8000) );
  DFF_X1 \REGISTERS_reg[16][33]  ( .D(n5983), .CK(CLK), .QN(n8017) );
  DFF_X1 \REGISTERS_reg[16][32]  ( .D(n5982), .CK(CLK), .QN(n8034) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n5981), .CK(CLK), .QN(n8051) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n5980), .CK(CLK), .QN(n8068) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n5979), .CK(CLK), .QN(n8085) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n5978), .CK(CLK), .QN(n8102) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n5977), .CK(CLK), .QN(n8119) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n5976), .CK(CLK), .QN(n8136) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n5975), .CK(CLK), .QN(n8153) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n5974), .CK(CLK), .QN(n8170) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n5515), .CK(CLK), .Q(n7131), .QN(n11820)
         );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n5514), .CK(CLK), .Q(n7105), .QN(n11819)
         );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n5513), .CK(CLK), .Q(n7101), .QN(n11818)
         );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n5512), .CK(CLK), .Q(n7097), .QN(n11817)
         );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n5511), .CK(CLK), .Q(n7093), .QN(n11816)
         );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n5510), .CK(CLK), .Q(n7089), .QN(n11815)
         );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n5509), .CK(CLK), .Q(n7085), .QN(n11814)
         );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n5508), .CK(CLK), .Q(n8614), .QN(n11813)
         );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n5507), .CK(CLK), .Q(n8606), .QN(n11812)
         );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n5506), .CK(CLK), .Q(n7081), .QN(n11811)
         );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n5769), .CK(CLK), .Q(n8626), .QN(n11810)
         );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n5768), .CK(CLK), .Q(n8624), .QN(n11809)
         );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n5767), .CK(CLK), .Q(n8622), .QN(n11808)
         );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n5765), .CK(CLK), .Q(n8618), .QN(n11807)
         );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n5764), .CK(CLK), .Q(n8612), .QN(n11806)
         );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n5763), .CK(CLK), .Q(n8604), .QN(n11805)
         );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n5762), .CK(CLK), .Q(n8600), .QN(n11804)
         );
  DFF_X1 \REGISTERS_reg[23][49]  ( .D(n5551), .CK(CLK), .Q(n7323), .QN(n11933)
         );
  DFF_X1 \REGISTERS_reg[23][48]  ( .D(n5550), .CK(CLK), .Q(n7319), .QN(n11932)
         );
  DFF_X1 \REGISTERS_reg[23][47]  ( .D(n5549), .CK(CLK), .Q(n7315), .QN(n11931)
         );
  DFF_X1 \REGISTERS_reg[23][46]  ( .D(n5548), .CK(CLK), .Q(n7311), .QN(n11930)
         );
  DFF_X1 \REGISTERS_reg[23][45]  ( .D(n5547), .CK(CLK), .Q(n7307), .QN(n11929)
         );
  DFF_X1 \REGISTERS_reg[23][44]  ( .D(n5546), .CK(CLK), .Q(n7303), .QN(n11928)
         );
  DFF_X1 \REGISTERS_reg[23][43]  ( .D(n5545), .CK(CLK), .Q(n7299), .QN(n11927)
         );
  DFF_X1 \REGISTERS_reg[23][42]  ( .D(n5544), .CK(CLK), .Q(n7295), .QN(n11926)
         );
  DFF_X1 \REGISTERS_reg[23][41]  ( .D(n5543), .CK(CLK), .Q(n7291), .QN(n11925)
         );
  DFF_X1 \REGISTERS_reg[23][40]  ( .D(n5542), .CK(CLK), .Q(n7287), .QN(n11924)
         );
  DFF_X1 \REGISTERS_reg[23][39]  ( .D(n5541), .CK(CLK), .Q(n7283), .QN(n11923)
         );
  DFF_X1 \REGISTERS_reg[23][38]  ( .D(n5540), .CK(CLK), .Q(n7279), .QN(n11922)
         );
  DFF_X1 \REGISTERS_reg[23][37]  ( .D(n5539), .CK(CLK), .Q(n8697), .QN(n11921)
         );
  DFF_X1 \REGISTERS_reg[23][36]  ( .D(n5538), .CK(CLK), .Q(n8698), .QN(n11920)
         );
  DFF_X1 \REGISTERS_reg[23][35]  ( .D(n5537), .CK(CLK), .Q(n8699), .QN(n11919)
         );
  DFF_X1 \REGISTERS_reg[23][34]  ( .D(n5536), .CK(CLK), .Q(n8700), .QN(n11918)
         );
  DFF_X1 \REGISTERS_reg[23][33]  ( .D(n5535), .CK(CLK), .Q(n8701), .QN(n11917)
         );
  DFF_X1 \REGISTERS_reg[23][32]  ( .D(n5534), .CK(CLK), .Q(n8702), .QN(n11916)
         );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n5533), .CK(CLK), .Q(n8703), .QN(n11915)
         );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n5532), .CK(CLK), .Q(n8704), .QN(n11914)
         );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n5531), .CK(CLK), .Q(n8705), .QN(n11913)
         );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n5530), .CK(CLK), .Q(n8706), .QN(n11912)
         );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n5529), .CK(CLK), .Q(n8707), .QN(n11911)
         );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n5528), .CK(CLK), .Q(n8708), .QN(n11910)
         );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n5653), .CK(CLK), .QN(n8188) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n5652), .CK(CLK), .QN(n8205) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n5651), .CK(CLK), .QN(n8222) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n5650), .CK(CLK), .QN(n8239) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n5649), .CK(CLK), .QN(n8256) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n5648), .CK(CLK), .QN(n8273) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n5647), .CK(CLK), .QN(n8290) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n5646), .CK(CLK), .QN(n8307) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n5645), .CK(CLK), .QN(n8324) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n5644), .CK(CLK), .QN(n8341) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n5643), .CK(CLK), .QN(n8358) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n5642), .CK(CLK), .QN(n8375) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n5641), .CK(CLK), .QN(n8392) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n5640), .CK(CLK), .QN(n8409) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n5639), .CK(CLK), .QN(n8426) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n5638), .CK(CLK), .QN(n8443) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n5637), .CK(CLK), .QN(n8460) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n5636), .CK(CLK), .QN(n8477) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n5635), .CK(CLK), .QN(n8494) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n5634), .CK(CLK), .QN(n8511) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n5633), .CK(CLK), .QN(n8528) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n5632), .CK(CLK), .QN(n8545) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n5631), .CK(CLK), .QN(n8562) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n5630), .CK(CLK), .QN(n8579) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n5717), .CK(CLK), .QN(n8189) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n5716), .CK(CLK), .QN(n8206) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n5715), .CK(CLK), .QN(n8223) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n5714), .CK(CLK), .QN(n8240) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n5713), .CK(CLK), .QN(n8257) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n5712), .CK(CLK), .QN(n8274) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n5711), .CK(CLK), .QN(n8291) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n5710), .CK(CLK), .QN(n8308) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n5709), .CK(CLK), .QN(n8325) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n5708), .CK(CLK), .QN(n8342) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n5707), .CK(CLK), .QN(n8359) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n5706), .CK(CLK), .QN(n8376) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n5705), .CK(CLK), .QN(n8393) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n5704), .CK(CLK), .QN(n8410) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n5703), .CK(CLK), .QN(n8427) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n5702), .CK(CLK), .QN(n8444) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n5701), .CK(CLK), .QN(n8461) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n5700), .CK(CLK), .QN(n8478) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n5699), .CK(CLK), .QN(n8495) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n5698), .CK(CLK), .QN(n8512) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n5697), .CK(CLK), .QN(n8529) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n5696), .CK(CLK), .QN(n8546) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n5695), .CK(CLK), .QN(n8563) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n5694), .CK(CLK), .QN(n8580) );
  DFF_X1 \REGISTERS_reg[19][46]  ( .D(n5804), .CK(CLK), .Q(n8696), .QN(n11909)
         );
  DFF_X1 \REGISTERS_reg[19][45]  ( .D(n5803), .CK(CLK), .Q(n8694), .QN(n11908)
         );
  DFF_X1 \REGISTERS_reg[19][44]  ( .D(n5802), .CK(CLK), .Q(n8692), .QN(n11907)
         );
  DFF_X1 \REGISTERS_reg[19][43]  ( .D(n5801), .CK(CLK), .Q(n8690), .QN(n11906)
         );
  DFF_X1 \REGISTERS_reg[19][42]  ( .D(n5800), .CK(CLK), .Q(n8688), .QN(n11905)
         );
  DFF_X1 \REGISTERS_reg[19][41]  ( .D(n5799), .CK(CLK), .Q(n8686), .QN(n11904)
         );
  DFF_X1 \REGISTERS_reg[19][40]  ( .D(n5798), .CK(CLK), .Q(n8684), .QN(n11903)
         );
  DFF_X1 \REGISTERS_reg[19][39]  ( .D(n5797), .CK(CLK), .Q(n8682), .QN(n11902)
         );
  DFF_X1 \REGISTERS_reg[19][38]  ( .D(n5796), .CK(CLK), .Q(n8680), .QN(n11901)
         );
  DFF_X1 \REGISTERS_reg[19][37]  ( .D(n5795), .CK(CLK), .Q(n8678), .QN(n11900)
         );
  DFF_X1 \REGISTERS_reg[19][36]  ( .D(n5794), .CK(CLK), .Q(n8676), .QN(n11899)
         );
  DFF_X1 \REGISTERS_reg[19][35]  ( .D(n5793), .CK(CLK), .Q(n8674), .QN(n11898)
         );
  DFF_X1 \REGISTERS_reg[19][34]  ( .D(n5792), .CK(CLK), .Q(n8672), .QN(n11897)
         );
  DFF_X1 \REGISTERS_reg[19][33]  ( .D(n5791), .CK(CLK), .Q(n8670), .QN(n11896)
         );
  DFF_X1 \REGISTERS_reg[19][32]  ( .D(n5790), .CK(CLK), .Q(n8668), .QN(n11895)
         );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n5789), .CK(CLK), .Q(n8666), .QN(n11894)
         );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n5788), .CK(CLK), .Q(n8664), .QN(n11893)
         );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n5787), .CK(CLK), .Q(n8662), .QN(n11892)
         );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n5786), .CK(CLK), .Q(n8660), .QN(n11891)
         );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n5785), .CK(CLK), .Q(n8658), .QN(n11890)
         );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n5784), .CK(CLK), .Q(n8656), .QN(n11889)
         );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n5783), .CK(CLK), .Q(n8654), .QN(n11888)
         );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n5782), .CK(CLK), .Q(n8652), .QN(n11887)
         );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n5774), .CK(CLK), .Q(n8636), .QN(n11803)
         );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n5909), .CK(CLK), .QN(n8186) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n5908), .CK(CLK), .QN(n8203) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n5907), .CK(CLK), .QN(n8220) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n5906), .CK(CLK), .QN(n8237) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n5905), .CK(CLK), .QN(n8254) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n5904), .CK(CLK), .QN(n8271) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n5903), .CK(CLK), .QN(n8288) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n5902), .CK(CLK), .QN(n8305) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n5901), .CK(CLK), .QN(n8322) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n5900), .CK(CLK), .QN(n8339) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n5899), .CK(CLK), .QN(n8356) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n5898), .CK(CLK), .QN(n8373) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n5897), .CK(CLK), .QN(n8390) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n5896), .CK(CLK), .QN(n8407) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n5895), .CK(CLK), .QN(n8424) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n5894), .CK(CLK), .QN(n8441) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n5893), .CK(CLK), .QN(n8458) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n5892), .CK(CLK), .QN(n8475) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n5891), .CK(CLK), .QN(n8492) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n5890), .CK(CLK), .QN(n8509) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n5889), .CK(CLK), .QN(n8526) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n5888), .CK(CLK), .QN(n8543) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n5887), .CK(CLK), .QN(n8560) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n5886), .CK(CLK), .QN(n8577) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n5973), .CK(CLK), .QN(n8187) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n5972), .CK(CLK), .QN(n8204) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n5971), .CK(CLK), .QN(n8221) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n5970), .CK(CLK), .QN(n8238) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n5969), .CK(CLK), .QN(n8255) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n5968), .CK(CLK), .QN(n8272) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n5967), .CK(CLK), .QN(n8289) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n5966), .CK(CLK), .QN(n8306) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n5965), .CK(CLK), .QN(n8323) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n5964), .CK(CLK), .QN(n8340) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n5963), .CK(CLK), .QN(n8357) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n5962), .CK(CLK), .QN(n8374) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n5961), .CK(CLK), .QN(n8391) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n5960), .CK(CLK), .QN(n8408) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n5959), .CK(CLK), .QN(n8425) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n5958), .CK(CLK), .QN(n8442) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n5957), .CK(CLK), .QN(n8459) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n5956), .CK(CLK), .QN(n8476) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n5955), .CK(CLK), .QN(n8493) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n5954), .CK(CLK), .QN(n8510) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n5953), .CK(CLK), .QN(n8527) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n5952), .CK(CLK), .QN(n8544) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n5951), .CK(CLK), .QN(n8561) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n5950), .CK(CLK), .QN(n8578) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n6974), .CK(CLK), .QN(n14216) );
  DFF_X1 \REGISTERS_reg[7][59]  ( .D(n6585), .CK(CLK), .Q(n11765), .QN(n7150)
         );
  DFF_X1 \REGISTERS_reg[7][58]  ( .D(n6584), .CK(CLK), .Q(n11641), .QN(n7247)
         );
  DFF_X1 \REGISTERS_reg[7][57]  ( .D(n6583), .CK(CLK), .Q(n11640), .QN(n7264)
         );
  DFF_X1 \REGISTERS_reg[7][56]  ( .D(n6582), .CK(CLK), .Q(n11639), .QN(n7363)
         );
  DFF_X1 \REGISTERS_reg[7][55]  ( .D(n6581), .CK(CLK), .Q(n11638), .QN(n7380)
         );
  DFF_X1 \REGISTERS_reg[7][54]  ( .D(n6580), .CK(CLK), .Q(n11637), .QN(n7397)
         );
  DFF_X1 \REGISTERS_reg[7][53]  ( .D(n6579), .CK(CLK), .Q(n11636), .QN(n7499)
         );
  DFF_X1 \REGISTERS_reg[7][52]  ( .D(n6578), .CK(CLK), .Q(n11635), .QN(n7516)
         );
  DFF_X1 \REGISTERS_reg[7][51]  ( .D(n6577), .CK(CLK), .Q(n11634), .QN(n7620)
         );
  DFF_X1 \REGISTERS_reg[7][50]  ( .D(n6576), .CK(CLK), .Q(n11633), .QN(n7637)
         );
  DFF_X1 \REGISTERS_reg[7][49]  ( .D(n6575), .CK(CLK), .Q(n11632), .QN(n7654)
         );
  DFF_X1 \REGISTERS_reg[7][48]  ( .D(n6574), .CK(CLK), .Q(n11631), .QN(n7756)
         );
  DFF_X1 \REGISTERS_reg[7][47]  ( .D(n6573), .CK(CLK), .Q(n11630), .QN(n7773)
         );
  DFF_X1 \REGISTERS_reg[7][46]  ( .D(n6572), .CK(CLK), .Q(n11629), .QN(n7790)
         );
  DFF_X1 \REGISTERS_reg[7][45]  ( .D(n6571), .CK(CLK), .Q(n11628), .QN(n7807)
         );
  DFF_X1 \REGISTERS_reg[7][44]  ( .D(n6570), .CK(CLK), .Q(n11627), .QN(n7824)
         );
  DFF_X1 \REGISTERS_reg[7][43]  ( .D(n6569), .CK(CLK), .Q(n11626), .QN(n7841)
         );
  DFF_X1 \REGISTERS_reg[7][42]  ( .D(n6568), .CK(CLK), .Q(n11625), .QN(n7858)
         );
  DFF_X1 \REGISTERS_reg[7][41]  ( .D(n6567), .CK(CLK), .Q(n11624), .QN(n7875)
         );
  DFF_X1 \REGISTERS_reg[7][40]  ( .D(n6566), .CK(CLK), .Q(n11623), .QN(n7892)
         );
  DFF_X1 \REGISTERS_reg[7][39]  ( .D(n6565), .CK(CLK), .Q(n11622), .QN(n7909)
         );
  DFF_X1 \REGISTERS_reg[7][38]  ( .D(n6564), .CK(CLK), .Q(n11621), .QN(n7926)
         );
  DFF_X1 \REGISTERS_reg[7][37]  ( .D(n6563), .CK(CLK), .Q(n11620), .QN(n7943)
         );
  DFF_X1 \REGISTERS_reg[7][36]  ( .D(n6562), .CK(CLK), .Q(n11619), .QN(n7960)
         );
  DFF_X1 \REGISTERS_reg[7][35]  ( .D(n6561), .CK(CLK), .Q(n11618), .QN(n7977)
         );
  DFF_X1 \REGISTERS_reg[7][34]  ( .D(n6560), .CK(CLK), .Q(n11617), .QN(n7994)
         );
  DFF_X1 \REGISTERS_reg[7][33]  ( .D(n6559), .CK(CLK), .Q(n11616), .QN(n8011)
         );
  DFF_X1 \REGISTERS_reg[7][32]  ( .D(n6558), .CK(CLK), .Q(n11615), .QN(n8028)
         );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n6557), .CK(CLK), .Q(n11614), .QN(n8045)
         );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n6556), .CK(CLK), .Q(n11613), .QN(n8062)
         );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n6555), .CK(CLK), .Q(n11612), .QN(n8079)
         );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n6554), .CK(CLK), .Q(n11611), .QN(n8096)
         );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n6553), .CK(CLK), .Q(n11610), .QN(n8113)
         );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n6552), .CK(CLK), .Q(n11609), .QN(n8130)
         );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n6551), .CK(CLK), .Q(n11608), .QN(n8147)
         );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n6550), .CK(CLK), .Q(n11607), .QN(n8164)
         );
  DFF_X1 \REGISTERS_reg[6][59]  ( .D(n6649), .CK(CLK), .Q(n11585), .QN(n7149)
         );
  DFF_X1 \REGISTERS_reg[6][58]  ( .D(n6648), .CK(CLK), .Q(n11461), .QN(n7246)
         );
  DFF_X1 \REGISTERS_reg[6][57]  ( .D(n6647), .CK(CLK), .Q(n11460), .QN(n7263)
         );
  DFF_X1 \REGISTERS_reg[6][56]  ( .D(n6646), .CK(CLK), .Q(n11459), .QN(n7362)
         );
  DFF_X1 \REGISTERS_reg[6][55]  ( .D(n6645), .CK(CLK), .Q(n11458), .QN(n7379)
         );
  DFF_X1 \REGISTERS_reg[6][54]  ( .D(n6644), .CK(CLK), .Q(n11457), .QN(n7396)
         );
  DFF_X1 \REGISTERS_reg[6][53]  ( .D(n6643), .CK(CLK), .Q(n11456), .QN(n7498)
         );
  DFF_X1 \REGISTERS_reg[6][52]  ( .D(n6642), .CK(CLK), .Q(n11455), .QN(n7515)
         );
  DFF_X1 \REGISTERS_reg[6][51]  ( .D(n6641), .CK(CLK), .Q(n11454), .QN(n7619)
         );
  DFF_X1 \REGISTERS_reg[6][50]  ( .D(n6640), .CK(CLK), .Q(n11453), .QN(n7636)
         );
  DFF_X1 \REGISTERS_reg[6][49]  ( .D(n6639), .CK(CLK), .Q(n11452), .QN(n7653)
         );
  DFF_X1 \REGISTERS_reg[6][48]  ( .D(n6638), .CK(CLK), .Q(n11451), .QN(n7755)
         );
  DFF_X1 \REGISTERS_reg[6][47]  ( .D(n6637), .CK(CLK), .Q(n11450), .QN(n7772)
         );
  DFF_X1 \REGISTERS_reg[6][46]  ( .D(n6636), .CK(CLK), .Q(n11449), .QN(n7789)
         );
  DFF_X1 \REGISTERS_reg[6][45]  ( .D(n6635), .CK(CLK), .Q(n11448), .QN(n7806)
         );
  DFF_X1 \REGISTERS_reg[6][44]  ( .D(n6634), .CK(CLK), .Q(n11447), .QN(n7823)
         );
  DFF_X1 \REGISTERS_reg[6][43]  ( .D(n6633), .CK(CLK), .Q(n11446), .QN(n7840)
         );
  DFF_X1 \REGISTERS_reg[6][42]  ( .D(n6632), .CK(CLK), .Q(n11445), .QN(n7857)
         );
  DFF_X1 \REGISTERS_reg[6][41]  ( .D(n6631), .CK(CLK), .Q(n11444), .QN(n7874)
         );
  DFF_X1 \REGISTERS_reg[6][40]  ( .D(n6630), .CK(CLK), .Q(n11443), .QN(n7891)
         );
  DFF_X1 \REGISTERS_reg[6][39]  ( .D(n6629), .CK(CLK), .Q(n11442), .QN(n7908)
         );
  DFF_X1 \REGISTERS_reg[6][38]  ( .D(n6628), .CK(CLK), .Q(n11441), .QN(n7925)
         );
  DFF_X1 \REGISTERS_reg[6][37]  ( .D(n6627), .CK(CLK), .Q(n11440), .QN(n7942)
         );
  DFF_X1 \REGISTERS_reg[6][36]  ( .D(n6626), .CK(CLK), .Q(n11439), .QN(n7959)
         );
  DFF_X1 \REGISTERS_reg[6][35]  ( .D(n6625), .CK(CLK), .Q(n11438), .QN(n7976)
         );
  DFF_X1 \REGISTERS_reg[6][34]  ( .D(n6624), .CK(CLK), .Q(n11437), .QN(n7993)
         );
  DFF_X1 \REGISTERS_reg[6][33]  ( .D(n6623), .CK(CLK), .Q(n11436), .QN(n8010)
         );
  DFF_X1 \REGISTERS_reg[6][32]  ( .D(n6622), .CK(CLK), .Q(n11435), .QN(n8027)
         );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n6621), .CK(CLK), .Q(n11434), .QN(n8044)
         );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n6620), .CK(CLK), .Q(n11433), .QN(n8061)
         );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n6619), .CK(CLK), .Q(n11432), .QN(n8078)
         );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n6618), .CK(CLK), .Q(n11431), .QN(n8095)
         );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n6617), .CK(CLK), .Q(n11430), .QN(n8112)
         );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n6616), .CK(CLK), .Q(n11429), .QN(n8129)
         );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n6615), .CK(CLK), .Q(n11428), .QN(n8146)
         );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n6614), .CK(CLK), .Q(n11427), .QN(n8163)
         );
  DFF_X1 \REGISTERS_reg[5][59]  ( .D(n6713), .CK(CLK), .QN(n14217) );
  DFF_X1 \REGISTERS_reg[5][58]  ( .D(n6712), .CK(CLK), .QN(n14218) );
  DFF_X1 \REGISTERS_reg[5][57]  ( .D(n6711), .CK(CLK), .QN(n14219) );
  DFF_X1 \REGISTERS_reg[5][56]  ( .D(n6710), .CK(CLK), .QN(n14220) );
  DFF_X1 \REGISTERS_reg[5][55]  ( .D(n6709), .CK(CLK), .QN(n14221) );
  DFF_X1 \REGISTERS_reg[5][54]  ( .D(n6708), .CK(CLK), .QN(n14222) );
  DFF_X1 \REGISTERS_reg[5][53]  ( .D(n6707), .CK(CLK), .QN(n14223) );
  DFF_X1 \REGISTERS_reg[5][52]  ( .D(n6706), .CK(CLK), .QN(n14224) );
  DFF_X1 \REGISTERS_reg[5][51]  ( .D(n6705), .CK(CLK), .QN(n14225) );
  DFF_X1 \REGISTERS_reg[5][50]  ( .D(n6704), .CK(CLK), .QN(n14226) );
  DFF_X1 \REGISTERS_reg[5][49]  ( .D(n6703), .CK(CLK), .QN(n14227) );
  DFF_X1 \REGISTERS_reg[5][48]  ( .D(n6702), .CK(CLK), .QN(n14228) );
  DFF_X1 \REGISTERS_reg[5][47]  ( .D(n6701), .CK(CLK), .QN(n14229) );
  DFF_X1 \REGISTERS_reg[5][46]  ( .D(n6700), .CK(CLK), .QN(n14230) );
  DFF_X1 \REGISTERS_reg[5][45]  ( .D(n6699), .CK(CLK), .QN(n14231) );
  DFF_X1 \REGISTERS_reg[5][44]  ( .D(n6698), .CK(CLK), .QN(n14232) );
  DFF_X1 \REGISTERS_reg[5][43]  ( .D(n6697), .CK(CLK), .QN(n14233) );
  DFF_X1 \REGISTERS_reg[5][42]  ( .D(n6696), .CK(CLK), .QN(n14234) );
  DFF_X1 \REGISTERS_reg[5][41]  ( .D(n6695), .CK(CLK), .QN(n14235) );
  DFF_X1 \REGISTERS_reg[5][40]  ( .D(n6694), .CK(CLK), .QN(n14236) );
  DFF_X1 \REGISTERS_reg[5][39]  ( .D(n6693), .CK(CLK), .QN(n14237) );
  DFF_X1 \REGISTERS_reg[5][38]  ( .D(n6692), .CK(CLK), .QN(n14238) );
  DFF_X1 \REGISTERS_reg[5][37]  ( .D(n6691), .CK(CLK), .QN(n14239) );
  DFF_X1 \REGISTERS_reg[5][36]  ( .D(n6690), .CK(CLK), .QN(n14240) );
  DFF_X1 \REGISTERS_reg[5][35]  ( .D(n6689), .CK(CLK), .QN(n14241) );
  DFF_X1 \REGISTERS_reg[5][34]  ( .D(n6688), .CK(CLK), .QN(n14242) );
  DFF_X1 \REGISTERS_reg[5][33]  ( .D(n6687), .CK(CLK), .QN(n14243) );
  DFF_X1 \REGISTERS_reg[5][32]  ( .D(n6686), .CK(CLK), .QN(n14244) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n6685), .CK(CLK), .QN(n14245) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n6684), .CK(CLK), .QN(n14246) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n6683), .CK(CLK), .QN(n14247) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n6682), .CK(CLK), .QN(n14248) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n6681), .CK(CLK), .QN(n14249) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n6680), .CK(CLK), .QN(n14250) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n6679), .CK(CLK), .QN(n14251) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n6678), .CK(CLK), .QN(n14252) );
  DFF_X1 \REGISTERS_reg[4][59]  ( .D(n6777), .CK(CLK), .QN(n14253) );
  DFF_X1 \REGISTERS_reg[4][58]  ( .D(n6776), .CK(CLK), .QN(n14254) );
  DFF_X1 \REGISTERS_reg[4][57]  ( .D(n6775), .CK(CLK), .QN(n14255) );
  DFF_X1 \REGISTERS_reg[4][56]  ( .D(n6774), .CK(CLK), .QN(n14256) );
  DFF_X1 \REGISTERS_reg[4][55]  ( .D(n6773), .CK(CLK), .QN(n14257) );
  DFF_X1 \REGISTERS_reg[4][54]  ( .D(n6772), .CK(CLK), .QN(n14258) );
  DFF_X1 \REGISTERS_reg[4][53]  ( .D(n6771), .CK(CLK), .QN(n14259) );
  DFF_X1 \REGISTERS_reg[4][52]  ( .D(n6770), .CK(CLK), .QN(n14260) );
  DFF_X1 \REGISTERS_reg[4][51]  ( .D(n6769), .CK(CLK), .QN(n14261) );
  DFF_X1 \REGISTERS_reg[4][50]  ( .D(n6768), .CK(CLK), .QN(n14262) );
  DFF_X1 \REGISTERS_reg[4][49]  ( .D(n6767), .CK(CLK), .QN(n14263) );
  DFF_X1 \REGISTERS_reg[4][48]  ( .D(n6766), .CK(CLK), .QN(n14264) );
  DFF_X1 \REGISTERS_reg[4][47]  ( .D(n6765), .CK(CLK), .QN(n14265) );
  DFF_X1 \REGISTERS_reg[4][46]  ( .D(n6764), .CK(CLK), .QN(n14266) );
  DFF_X1 \REGISTERS_reg[4][45]  ( .D(n6763), .CK(CLK), .QN(n14267) );
  DFF_X1 \REGISTERS_reg[4][44]  ( .D(n6762), .CK(CLK), .QN(n14268) );
  DFF_X1 \REGISTERS_reg[4][43]  ( .D(n6761), .CK(CLK), .QN(n14269) );
  DFF_X1 \REGISTERS_reg[4][42]  ( .D(n6760), .CK(CLK), .QN(n14270) );
  DFF_X1 \REGISTERS_reg[4][41]  ( .D(n6759), .CK(CLK), .QN(n14271) );
  DFF_X1 \REGISTERS_reg[4][40]  ( .D(n6758), .CK(CLK), .QN(n14272) );
  DFF_X1 \REGISTERS_reg[4][39]  ( .D(n6757), .CK(CLK), .QN(n14273) );
  DFF_X1 \REGISTERS_reg[4][38]  ( .D(n6756), .CK(CLK), .QN(n14274) );
  DFF_X1 \REGISTERS_reg[4][37]  ( .D(n6755), .CK(CLK), .QN(n14275) );
  DFF_X1 \REGISTERS_reg[4][36]  ( .D(n6754), .CK(CLK), .QN(n14276) );
  DFF_X1 \REGISTERS_reg[4][35]  ( .D(n6753), .CK(CLK), .QN(n14277) );
  DFF_X1 \REGISTERS_reg[4][34]  ( .D(n6752), .CK(CLK), .QN(n14278) );
  DFF_X1 \REGISTERS_reg[4][33]  ( .D(n6751), .CK(CLK), .QN(n14279) );
  DFF_X1 \REGISTERS_reg[4][32]  ( .D(n6750), .CK(CLK), .QN(n14280) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n6749), .CK(CLK), .QN(n14281) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n6748), .CK(CLK), .QN(n14282) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n6747), .CK(CLK), .QN(n14283) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n6746), .CK(CLK), .QN(n14284) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n6745), .CK(CLK), .QN(n14285) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n6744), .CK(CLK), .QN(n14286) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n6743), .CK(CLK), .QN(n14287) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n6742), .CK(CLK), .QN(n14288) );
  DFF_X1 \REGISTERS_reg[3][59]  ( .D(n6841), .CK(CLK), .Q(n9953), .QN(n11994)
         );
  DFF_X1 \REGISTERS_reg[3][58]  ( .D(n6840), .CK(CLK), .Q(n9954), .QN(n11993)
         );
  DFF_X1 \REGISTERS_reg[3][57]  ( .D(n6839), .CK(CLK), .Q(n9955), .QN(n11992)
         );
  DFF_X1 \REGISTERS_reg[3][56]  ( .D(n6838), .CK(CLK), .Q(n9956), .QN(n11991)
         );
  DFF_X1 \REGISTERS_reg[3][55]  ( .D(n6837), .CK(CLK), .Q(n9957), .QN(n11990)
         );
  DFF_X1 \REGISTERS_reg[3][54]  ( .D(n6836), .CK(CLK), .Q(n9958), .QN(n11989)
         );
  DFF_X1 \REGISTERS_reg[3][53]  ( .D(n6835), .CK(CLK), .Q(n9959), .QN(n11988)
         );
  DFF_X1 \REGISTERS_reg[3][52]  ( .D(n6834), .CK(CLK), .Q(n9960), .QN(n11987)
         );
  DFF_X1 \REGISTERS_reg[3][51]  ( .D(n6833), .CK(CLK), .Q(n9961), .QN(n11986)
         );
  DFF_X1 \REGISTERS_reg[3][50]  ( .D(n6832), .CK(CLK), .Q(n9962), .QN(n11985)
         );
  DFF_X1 \REGISTERS_reg[3][49]  ( .D(n6831), .CK(CLK), .Q(n9963), .QN(n11984)
         );
  DFF_X1 \REGISTERS_reg[3][48]  ( .D(n6830), .CK(CLK), .Q(n9964), .QN(n11983)
         );
  DFF_X1 \REGISTERS_reg[3][47]  ( .D(n6829), .CK(CLK), .Q(n9965), .QN(n11982)
         );
  DFF_X1 \REGISTERS_reg[3][46]  ( .D(n6828), .CK(CLK), .Q(n9966), .QN(n11981)
         );
  DFF_X1 \REGISTERS_reg[3][45]  ( .D(n6827), .CK(CLK), .Q(n9967), .QN(n11980)
         );
  DFF_X1 \REGISTERS_reg[3][44]  ( .D(n6826), .CK(CLK), .Q(n9968), .QN(n11979)
         );
  DFF_X1 \REGISTERS_reg[3][43]  ( .D(n6825), .CK(CLK), .Q(n9969), .QN(n11978)
         );
  DFF_X1 \REGISTERS_reg[3][42]  ( .D(n6824), .CK(CLK), .Q(n9970), .QN(n11977)
         );
  DFF_X1 \REGISTERS_reg[3][41]  ( .D(n6823), .CK(CLK), .Q(n9971), .QN(n11976)
         );
  DFF_X1 \REGISTERS_reg[3][40]  ( .D(n6822), .CK(CLK), .Q(n9972), .QN(n11975)
         );
  DFF_X1 \REGISTERS_reg[3][39]  ( .D(n6821), .CK(CLK), .Q(n9973), .QN(n11974)
         );
  DFF_X1 \REGISTERS_reg[3][38]  ( .D(n6820), .CK(CLK), .Q(n9974), .QN(n11973)
         );
  DFF_X1 \REGISTERS_reg[3][37]  ( .D(n6819), .CK(CLK), .Q(n9975), .QN(n11972)
         );
  DFF_X1 \REGISTERS_reg[3][36]  ( .D(n6818), .CK(CLK), .Q(n9976), .QN(n11971)
         );
  DFF_X1 \REGISTERS_reg[3][35]  ( .D(n6817), .CK(CLK), .Q(n9977), .QN(n11970)
         );
  DFF_X1 \REGISTERS_reg[3][34]  ( .D(n6816), .CK(CLK), .Q(n9978), .QN(n11969)
         );
  DFF_X1 \REGISTERS_reg[3][33]  ( .D(n6815), .CK(CLK), .Q(n9979), .QN(n11968)
         );
  DFF_X1 \REGISTERS_reg[3][32]  ( .D(n6814), .CK(CLK), .Q(n9980), .QN(n11967)
         );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n6813), .CK(CLK), .Q(n9981), .QN(n11966)
         );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n6812), .CK(CLK), .Q(n9982), .QN(n11965)
         );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n6811), .CK(CLK), .Q(n9983), .QN(n11964)
         );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n6810), .CK(CLK), .Q(n9984), .QN(n11963)
         );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n6809), .CK(CLK), .Q(n9985), .QN(n11962)
         );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n6808), .CK(CLK), .Q(n9986), .QN(n11961)
         );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n6807), .CK(CLK), .Q(n9987), .QN(n11960)
         );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n6806), .CK(CLK), .Q(n9988), .QN(n11959)
         );
  DFF_X1 \REGISTERS_reg[2][59]  ( .D(n6905), .CK(CLK), .Q(n9889), .QN(n11886)
         );
  DFF_X1 \REGISTERS_reg[2][58]  ( .D(n6904), .CK(CLK), .Q(n9890), .QN(n11885)
         );
  DFF_X1 \REGISTERS_reg[2][57]  ( .D(n6903), .CK(CLK), .Q(n9891), .QN(n11884)
         );
  DFF_X1 \REGISTERS_reg[2][56]  ( .D(n6902), .CK(CLK), .Q(n9892), .QN(n11883)
         );
  DFF_X1 \REGISTERS_reg[2][55]  ( .D(n6901), .CK(CLK), .Q(n9893), .QN(n11882)
         );
  DFF_X1 \REGISTERS_reg[2][54]  ( .D(n6900), .CK(CLK), .Q(n9894), .QN(n11881)
         );
  DFF_X1 \REGISTERS_reg[2][53]  ( .D(n6899), .CK(CLK), .Q(n9895), .QN(n11880)
         );
  DFF_X1 \REGISTERS_reg[2][52]  ( .D(n6898), .CK(CLK), .Q(n9896), .QN(n11879)
         );
  DFF_X1 \REGISTERS_reg[2][51]  ( .D(n6897), .CK(CLK), .Q(n9897), .QN(n11878)
         );
  DFF_X1 \REGISTERS_reg[2][50]  ( .D(n6896), .CK(CLK), .Q(n9898), .QN(n11877)
         );
  DFF_X1 \REGISTERS_reg[2][49]  ( .D(n6895), .CK(CLK), .Q(n9899), .QN(n11876)
         );
  DFF_X1 \REGISTERS_reg[2][48]  ( .D(n6894), .CK(CLK), .Q(n9900), .QN(n11875)
         );
  DFF_X1 \REGISTERS_reg[2][47]  ( .D(n6893), .CK(CLK), .Q(n9901), .QN(n11874)
         );
  DFF_X1 \REGISTERS_reg[2][46]  ( .D(n6892), .CK(CLK), .Q(n9902), .QN(n11873)
         );
  DFF_X1 \REGISTERS_reg[2][45]  ( .D(n6891), .CK(CLK), .Q(n9903), .QN(n11872)
         );
  DFF_X1 \REGISTERS_reg[2][44]  ( .D(n6890), .CK(CLK), .Q(n9904), .QN(n11871)
         );
  DFF_X1 \REGISTERS_reg[2][43]  ( .D(n6889), .CK(CLK), .Q(n9905), .QN(n11870)
         );
  DFF_X1 \REGISTERS_reg[2][42]  ( .D(n6888), .CK(CLK), .Q(n9906), .QN(n11869)
         );
  DFF_X1 \REGISTERS_reg[2][41]  ( .D(n6887), .CK(CLK), .Q(n9907), .QN(n11868)
         );
  DFF_X1 \REGISTERS_reg[2][40]  ( .D(n6886), .CK(CLK), .Q(n9908), .QN(n11867)
         );
  DFF_X1 \REGISTERS_reg[2][39]  ( .D(n6885), .CK(CLK), .Q(n9909), .QN(n11866)
         );
  DFF_X1 \REGISTERS_reg[2][38]  ( .D(n6884), .CK(CLK), .Q(n9910), .QN(n11865)
         );
  DFF_X1 \REGISTERS_reg[2][37]  ( .D(n6883), .CK(CLK), .Q(n9911), .QN(n11864)
         );
  DFF_X1 \REGISTERS_reg[2][36]  ( .D(n6882), .CK(CLK), .Q(n9912), .QN(n11863)
         );
  DFF_X1 \REGISTERS_reg[2][35]  ( .D(n6881), .CK(CLK), .Q(n9913), .QN(n11862)
         );
  DFF_X1 \REGISTERS_reg[2][34]  ( .D(n6880), .CK(CLK), .Q(n9914), .QN(n11861)
         );
  DFF_X1 \REGISTERS_reg[2][33]  ( .D(n6879), .CK(CLK), .Q(n9915), .QN(n11860)
         );
  DFF_X1 \REGISTERS_reg[2][32]  ( .D(n6878), .CK(CLK), .Q(n9916), .QN(n11859)
         );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n6877), .CK(CLK), .Q(n9917), .QN(n11858)
         );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n6876), .CK(CLK), .Q(n9918), .QN(n11857)
         );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n6875), .CK(CLK), .Q(n9919), .QN(n11856)
         );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n6874), .CK(CLK), .Q(n9920), .QN(n11855)
         );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n6873), .CK(CLK), .Q(n9921), .QN(n11854)
         );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n6872), .CK(CLK), .Q(n9922), .QN(n11853)
         );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n6871), .CK(CLK), .Q(n9923), .QN(n11852)
         );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n6870), .CK(CLK), .Q(n9924), .QN(n11851)
         );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n7003), .CK(CLK), .QN(n14289) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n7002), .CK(CLK), .QN(n14290) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n7001), .CK(CLK), .QN(n14291) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n7000), .CK(CLK), .QN(n14292) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n6999), .CK(CLK), .QN(n14293) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n6998), .CK(CLK), .QN(n14294) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n6997), .CK(CLK), .QN(n14295) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n6996), .CK(CLK), .QN(n14296) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n6995), .CK(CLK), .QN(n14297) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n6994), .CK(CLK), .QN(n14298) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n6993), .CK(CLK), .QN(n14299) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n6992), .CK(CLK), .QN(n14300) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n6991), .CK(CLK), .QN(n14301) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n6990), .CK(CLK), .QN(n14302) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n6989), .CK(CLK), .QN(n14303) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n6988), .CK(CLK), .QN(n14304) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n6987), .CK(CLK), .QN(n14305) );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n6986), .CK(CLK), .QN(n14306) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n6985), .CK(CLK), .QN(n14307) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n6984), .CK(CLK), .QN(n14308) );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n6983), .CK(CLK), .QN(n14309) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n6981), .CK(CLK), .QN(n14310) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n6980), .CK(CLK), .QN(n14311) );
  DFF_X1 \REGISTERS_reg[1][39]  ( .D(n6949), .CK(CLK), .QN(n14312) );
  DFF_X1 \REGISTERS_reg[1][38]  ( .D(n6948), .CK(CLK), .QN(n14313) );
  DFF_X1 \REGISTERS_reg[1][37]  ( .D(n6947), .CK(CLK), .QN(n14314) );
  DFF_X1 \REGISTERS_reg[1][36]  ( .D(n6946), .CK(CLK), .QN(n14315) );
  DFF_X1 \REGISTERS_reg[1][35]  ( .D(n6945), .CK(CLK), .QN(n14316) );
  DFF_X1 \REGISTERS_reg[1][34]  ( .D(n6944), .CK(CLK), .QN(n14317) );
  DFF_X1 \REGISTERS_reg[1][33]  ( .D(n6943), .CK(CLK), .QN(n14318) );
  DFF_X1 \REGISTERS_reg[1][32]  ( .D(n6942), .CK(CLK), .QN(n14319) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n6941), .CK(CLK), .QN(n14320) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n6940), .CK(CLK), .QN(n14321) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n6939), .CK(CLK), .QN(n14322) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n6982), .CK(CLK), .QN(n14323) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n6979), .CK(CLK), .QN(n14324) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n6978), .CK(CLK), .QN(n14325) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n6977), .CK(CLK), .QN(n14326) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n6976), .CK(CLK), .QN(n14327) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n6975), .CK(CLK), .QN(n14328) );
  DFF_X1 \REGISTERS_reg[9][59]  ( .D(n6457), .CK(CLK), .Q(n11521), .QN(n7151)
         );
  DFF_X1 \REGISTERS_reg[9][58]  ( .D(n6456), .CK(CLK), .Q(n11520), .QN(n7248)
         );
  DFF_X1 \REGISTERS_reg[9][57]  ( .D(n6455), .CK(CLK), .Q(n11519), .QN(n7265)
         );
  DFF_X1 \REGISTERS_reg[9][56]  ( .D(n6454), .CK(CLK), .Q(n11518), .QN(n7364)
         );
  DFF_X1 \REGISTERS_reg[9][55]  ( .D(n6453), .CK(CLK), .Q(n11517), .QN(n7381)
         );
  DFF_X1 \REGISTERS_reg[9][54]  ( .D(n6452), .CK(CLK), .Q(n11516), .QN(n7398)
         );
  DFF_X1 \REGISTERS_reg[9][53]  ( .D(n6451), .CK(CLK), .Q(n11515), .QN(n7500)
         );
  DFF_X1 \REGISTERS_reg[9][52]  ( .D(n6450), .CK(CLK), .Q(n11514), .QN(n7517)
         );
  DFF_X1 \REGISTERS_reg[9][51]  ( .D(n6449), .CK(CLK), .Q(n11513), .QN(n7621)
         );
  DFF_X1 \REGISTERS_reg[9][50]  ( .D(n6448), .CK(CLK), .Q(n11512), .QN(n7638)
         );
  DFF_X1 \REGISTERS_reg[9][49]  ( .D(n6447), .CK(CLK), .Q(n11511), .QN(n7655)
         );
  DFF_X1 \REGISTERS_reg[9][48]  ( .D(n6446), .CK(CLK), .Q(n11510), .QN(n7757)
         );
  DFF_X1 \REGISTERS_reg[9][47]  ( .D(n6445), .CK(CLK), .Q(n11509), .QN(n7774)
         );
  DFF_X1 \REGISTERS_reg[9][46]  ( .D(n6444), .CK(CLK), .Q(n11508), .QN(n7791)
         );
  DFF_X1 \REGISTERS_reg[9][45]  ( .D(n6443), .CK(CLK), .Q(n11507), .QN(n7808)
         );
  DFF_X1 \REGISTERS_reg[9][44]  ( .D(n6442), .CK(CLK), .Q(n11506), .QN(n7825)
         );
  DFF_X1 \REGISTERS_reg[9][43]  ( .D(n6441), .CK(CLK), .Q(n11505), .QN(n7842)
         );
  DFF_X1 \REGISTERS_reg[9][42]  ( .D(n6440), .CK(CLK), .Q(n11504), .QN(n7859)
         );
  DFF_X1 \REGISTERS_reg[9][41]  ( .D(n6439), .CK(CLK), .Q(n11503), .QN(n7876)
         );
  DFF_X1 \REGISTERS_reg[9][40]  ( .D(n6438), .CK(CLK), .Q(n11502), .QN(n7893)
         );
  DFF_X1 \REGISTERS_reg[9][39]  ( .D(n6437), .CK(CLK), .Q(n11501), .QN(n7910)
         );
  DFF_X1 \REGISTERS_reg[9][38]  ( .D(n6436), .CK(CLK), .Q(n11500), .QN(n7927)
         );
  DFF_X1 \REGISTERS_reg[9][37]  ( .D(n6435), .CK(CLK), .Q(n11499), .QN(n7944)
         );
  DFF_X1 \REGISTERS_reg[9][36]  ( .D(n6434), .CK(CLK), .Q(n11498), .QN(n7961)
         );
  DFF_X1 \REGISTERS_reg[9][35]  ( .D(n6433), .CK(CLK), .Q(n11497), .QN(n7978)
         );
  DFF_X1 \REGISTERS_reg[9][34]  ( .D(n6432), .CK(CLK), .Q(n11496), .QN(n7995)
         );
  DFF_X1 \REGISTERS_reg[9][33]  ( .D(n6431), .CK(CLK), .Q(n11495), .QN(n8012)
         );
  DFF_X1 \REGISTERS_reg[9][32]  ( .D(n6430), .CK(CLK), .Q(n11494), .QN(n8029)
         );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n6429), .CK(CLK), .Q(n11493), .QN(n8046)
         );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n6428), .CK(CLK), .Q(n11492), .QN(n8063)
         );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n6427), .CK(CLK), .Q(n11491), .QN(n8080)
         );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n6426), .CK(CLK), .Q(n11490), .QN(n8097)
         );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n6425), .CK(CLK), .Q(n11489), .QN(n8114)
         );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n6424), .CK(CLK), .Q(n11488), .QN(n8131)
         );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n6423), .CK(CLK), .Q(n11487), .QN(n8148)
         );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n6422), .CK(CLK), .Q(n11486), .QN(n8165)
         );
  DFF_X1 \REGISTERS_reg[8][59]  ( .D(n6521), .CK(CLK), .Q(n11701), .QN(n7152)
         );
  DFF_X1 \REGISTERS_reg[8][58]  ( .D(n6520), .CK(CLK), .Q(n11700), .QN(n7249)
         );
  DFF_X1 \REGISTERS_reg[8][57]  ( .D(n6519), .CK(CLK), .Q(n11699), .QN(n7266)
         );
  DFF_X1 \REGISTERS_reg[8][56]  ( .D(n6518), .CK(CLK), .Q(n11698), .QN(n7365)
         );
  DFF_X1 \REGISTERS_reg[8][55]  ( .D(n6517), .CK(CLK), .Q(n11697), .QN(n7382)
         );
  DFF_X1 \REGISTERS_reg[8][54]  ( .D(n6516), .CK(CLK), .Q(n11696), .QN(n7399)
         );
  DFF_X1 \REGISTERS_reg[8][53]  ( .D(n6515), .CK(CLK), .Q(n11695), .QN(n7501)
         );
  DFF_X1 \REGISTERS_reg[8][52]  ( .D(n6514), .CK(CLK), .Q(n11694), .QN(n7518)
         );
  DFF_X1 \REGISTERS_reg[8][51]  ( .D(n6513), .CK(CLK), .Q(n11693), .QN(n7622)
         );
  DFF_X1 \REGISTERS_reg[8][50]  ( .D(n6512), .CK(CLK), .Q(n11692), .QN(n7639)
         );
  DFF_X1 \REGISTERS_reg[8][49]  ( .D(n6511), .CK(CLK), .Q(n11691), .QN(n7656)
         );
  DFF_X1 \REGISTERS_reg[8][48]  ( .D(n6510), .CK(CLK), .Q(n11690), .QN(n7758)
         );
  DFF_X1 \REGISTERS_reg[8][47]  ( .D(n6509), .CK(CLK), .Q(n11689), .QN(n7775)
         );
  DFF_X1 \REGISTERS_reg[8][46]  ( .D(n6508), .CK(CLK), .Q(n11688), .QN(n7792)
         );
  DFF_X1 \REGISTERS_reg[8][45]  ( .D(n6507), .CK(CLK), .Q(n11687), .QN(n7809)
         );
  DFF_X1 \REGISTERS_reg[8][44]  ( .D(n6506), .CK(CLK), .Q(n11686), .QN(n7826)
         );
  DFF_X1 \REGISTERS_reg[8][43]  ( .D(n6505), .CK(CLK), .Q(n11685), .QN(n7843)
         );
  DFF_X1 \REGISTERS_reg[8][42]  ( .D(n6504), .CK(CLK), .Q(n11684), .QN(n7860)
         );
  DFF_X1 \REGISTERS_reg[8][41]  ( .D(n6503), .CK(CLK), .Q(n11683), .QN(n7877)
         );
  DFF_X1 \REGISTERS_reg[8][40]  ( .D(n6502), .CK(CLK), .Q(n11682), .QN(n7894)
         );
  DFF_X1 \REGISTERS_reg[8][39]  ( .D(n6501), .CK(CLK), .Q(n11681), .QN(n7911)
         );
  DFF_X1 \REGISTERS_reg[8][38]  ( .D(n6500), .CK(CLK), .Q(n11680), .QN(n7928)
         );
  DFF_X1 \REGISTERS_reg[8][37]  ( .D(n6499), .CK(CLK), .Q(n11679), .QN(n7945)
         );
  DFF_X1 \REGISTERS_reg[8][36]  ( .D(n6498), .CK(CLK), .Q(n11678), .QN(n7962)
         );
  DFF_X1 \REGISTERS_reg[8][35]  ( .D(n6497), .CK(CLK), .Q(n11677), .QN(n7979)
         );
  DFF_X1 \REGISTERS_reg[8][34]  ( .D(n6496), .CK(CLK), .Q(n11676), .QN(n7996)
         );
  DFF_X1 \REGISTERS_reg[8][33]  ( .D(n6495), .CK(CLK), .Q(n11675), .QN(n8013)
         );
  DFF_X1 \REGISTERS_reg[8][32]  ( .D(n6494), .CK(CLK), .Q(n11674), .QN(n8030)
         );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n6493), .CK(CLK), .Q(n11673), .QN(n8047)
         );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n6492), .CK(CLK), .Q(n11672), .QN(n8064)
         );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n6491), .CK(CLK), .Q(n11671), .QN(n8081)
         );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n6490), .CK(CLK), .Q(n11670), .QN(n8098)
         );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n6489), .CK(CLK), .Q(n11669), .QN(n8115)
         );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n6488), .CK(CLK), .Q(n11668), .QN(n8132)
         );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n6487), .CK(CLK), .Q(n11667), .QN(n8149)
         );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n6486), .CK(CLK), .Q(n11666), .QN(n8166)
         );
  DFF_X1 \REGISTERS_reg[12][59]  ( .D(n6265), .CK(CLK), .Q(n11761), .QN(n7234)
         );
  DFF_X1 \REGISTERS_reg[12][58]  ( .D(n6264), .CK(CLK), .Q(n11760), .QN(n7251)
         );
  DFF_X1 \REGISTERS_reg[12][57]  ( .D(n6263), .CK(CLK), .Q(n11759), .QN(n7268)
         );
  DFF_X1 \REGISTERS_reg[12][56]  ( .D(n6262), .CK(CLK), .Q(n11758), .QN(n7367)
         );
  DFF_X1 \REGISTERS_reg[12][55]  ( .D(n6261), .CK(CLK), .Q(n11757), .QN(n7384)
         );
  DFF_X1 \REGISTERS_reg[12][54]  ( .D(n6260), .CK(CLK), .Q(n11756), .QN(n7401)
         );
  DFF_X1 \REGISTERS_reg[12][53]  ( .D(n6259), .CK(CLK), .Q(n11755), .QN(n7503)
         );
  DFF_X1 \REGISTERS_reg[12][52]  ( .D(n6258), .CK(CLK), .Q(n11754), .QN(n7520)
         );
  DFF_X1 \REGISTERS_reg[12][51]  ( .D(n6257), .CK(CLK), .Q(n11753), .QN(n7624)
         );
  DFF_X1 \REGISTERS_reg[12][50]  ( .D(n6256), .CK(CLK), .Q(n11752), .QN(n7641)
         );
  DFF_X1 \REGISTERS_reg[12][49]  ( .D(n6255), .CK(CLK), .Q(n11751), .QN(n7743)
         );
  DFF_X1 \REGISTERS_reg[12][48]  ( .D(n6254), .CK(CLK), .Q(n11750), .QN(n7760)
         );
  DFF_X1 \REGISTERS_reg[12][47]  ( .D(n6253), .CK(CLK), .Q(n11749), .QN(n7777)
         );
  DFF_X1 \REGISTERS_reg[12][46]  ( .D(n6252), .CK(CLK), .Q(n11748), .QN(n7794)
         );
  DFF_X1 \REGISTERS_reg[12][45]  ( .D(n6251), .CK(CLK), .Q(n11747), .QN(n7811)
         );
  DFF_X1 \REGISTERS_reg[12][44]  ( .D(n6250), .CK(CLK), .Q(n11746), .QN(n7828)
         );
  DFF_X1 \REGISTERS_reg[12][43]  ( .D(n6249), .CK(CLK), .Q(n11745), .QN(n7845)
         );
  DFF_X1 \REGISTERS_reg[12][42]  ( .D(n6248), .CK(CLK), .Q(n11744), .QN(n7862)
         );
  DFF_X1 \REGISTERS_reg[12][41]  ( .D(n6247), .CK(CLK), .Q(n11743), .QN(n7879)
         );
  DFF_X1 \REGISTERS_reg[12][40]  ( .D(n6246), .CK(CLK), .Q(n11742), .QN(n7896)
         );
  DFF_X1 \REGISTERS_reg[12][39]  ( .D(n6245), .CK(CLK), .Q(n11741), .QN(n7913)
         );
  DFF_X1 \REGISTERS_reg[12][38]  ( .D(n6244), .CK(CLK), .Q(n11740), .QN(n7930)
         );
  DFF_X1 \REGISTERS_reg[12][37]  ( .D(n6243), .CK(CLK), .Q(n11739), .QN(n7947)
         );
  DFF_X1 \REGISTERS_reg[12][36]  ( .D(n6242), .CK(CLK), .Q(n11738), .QN(n7964)
         );
  DFF_X1 \REGISTERS_reg[12][35]  ( .D(n6241), .CK(CLK), .Q(n11737), .QN(n7981)
         );
  DFF_X1 \REGISTERS_reg[12][34]  ( .D(n6240), .CK(CLK), .Q(n11736), .QN(n7998)
         );
  DFF_X1 \REGISTERS_reg[12][33]  ( .D(n6239), .CK(CLK), .Q(n11735), .QN(n8015)
         );
  DFF_X1 \REGISTERS_reg[12][32]  ( .D(n6238), .CK(CLK), .Q(n11734), .QN(n8032)
         );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n6237), .CK(CLK), .Q(n11733), .QN(n8049)
         );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n6236), .CK(CLK), .Q(n11732), .QN(n8066)
         );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n6235), .CK(CLK), .Q(n11731), .QN(n8083)
         );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n6234), .CK(CLK), .Q(n11730), .QN(n8100)
         );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n6233), .CK(CLK), .Q(n11729), .QN(n8117)
         );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n6232), .CK(CLK), .Q(n11728), .QN(n8134)
         );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n6231), .CK(CLK), .Q(n11727), .QN(n8151)
         );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n6230), .CK(CLK), .Q(n11726), .QN(n8168)
         );
  DFF_X1 \REGISTERS_reg[13][59]  ( .D(n6201), .CK(CLK), .Q(n11581), .QN(n7153)
         );
  DFF_X1 \REGISTERS_reg[13][58]  ( .D(n6200), .CK(CLK), .Q(n11580), .QN(n7250)
         );
  DFF_X1 \REGISTERS_reg[13][57]  ( .D(n6199), .CK(CLK), .Q(n11579), .QN(n7267)
         );
  DFF_X1 \REGISTERS_reg[13][56]  ( .D(n6198), .CK(CLK), .Q(n11578), .QN(n7366)
         );
  DFF_X1 \REGISTERS_reg[13][55]  ( .D(n6197), .CK(CLK), .Q(n11577), .QN(n7383)
         );
  DFF_X1 \REGISTERS_reg[13][54]  ( .D(n6196), .CK(CLK), .Q(n11576), .QN(n7400)
         );
  DFF_X1 \REGISTERS_reg[13][53]  ( .D(n6195), .CK(CLK), .Q(n11575), .QN(n7502)
         );
  DFF_X1 \REGISTERS_reg[13][52]  ( .D(n6194), .CK(CLK), .Q(n11574), .QN(n7519)
         );
  DFF_X1 \REGISTERS_reg[13][51]  ( .D(n6193), .CK(CLK), .Q(n11573), .QN(n7623)
         );
  DFF_X1 \REGISTERS_reg[13][50]  ( .D(n6192), .CK(CLK), .Q(n11572), .QN(n7640)
         );
  DFF_X1 \REGISTERS_reg[13][49]  ( .D(n6191), .CK(CLK), .Q(n11571), .QN(n7742)
         );
  DFF_X1 \REGISTERS_reg[13][48]  ( .D(n6190), .CK(CLK), .Q(n11570), .QN(n7759)
         );
  DFF_X1 \REGISTERS_reg[13][47]  ( .D(n6189), .CK(CLK), .Q(n11569), .QN(n7776)
         );
  DFF_X1 \REGISTERS_reg[13][46]  ( .D(n6188), .CK(CLK), .Q(n11568), .QN(n7793)
         );
  DFF_X1 \REGISTERS_reg[13][45]  ( .D(n6187), .CK(CLK), .Q(n11567), .QN(n7810)
         );
  DFF_X1 \REGISTERS_reg[13][44]  ( .D(n6186), .CK(CLK), .Q(n11566), .QN(n7827)
         );
  DFF_X1 \REGISTERS_reg[13][43]  ( .D(n6185), .CK(CLK), .Q(n11565), .QN(n7844)
         );
  DFF_X1 \REGISTERS_reg[13][42]  ( .D(n6184), .CK(CLK), .Q(n11564), .QN(n7861)
         );
  DFF_X1 \REGISTERS_reg[13][41]  ( .D(n6183), .CK(CLK), .Q(n11563), .QN(n7878)
         );
  DFF_X1 \REGISTERS_reg[13][40]  ( .D(n6182), .CK(CLK), .Q(n11562), .QN(n7895)
         );
  DFF_X1 \REGISTERS_reg[13][39]  ( .D(n6181), .CK(CLK), .Q(n11561), .QN(n7912)
         );
  DFF_X1 \REGISTERS_reg[13][38]  ( .D(n6180), .CK(CLK), .Q(n11560), .QN(n7929)
         );
  DFF_X1 \REGISTERS_reg[13][37]  ( .D(n6179), .CK(CLK), .Q(n11559), .QN(n7946)
         );
  DFF_X1 \REGISTERS_reg[13][36]  ( .D(n6178), .CK(CLK), .Q(n11558), .QN(n7963)
         );
  DFF_X1 \REGISTERS_reg[13][35]  ( .D(n6177), .CK(CLK), .Q(n11557), .QN(n7980)
         );
  DFF_X1 \REGISTERS_reg[13][34]  ( .D(n6176), .CK(CLK), .Q(n11556), .QN(n7997)
         );
  DFF_X1 \REGISTERS_reg[13][33]  ( .D(n6175), .CK(CLK), .Q(n11555), .QN(n8014)
         );
  DFF_X1 \REGISTERS_reg[13][32]  ( .D(n6174), .CK(CLK), .Q(n11554), .QN(n8031)
         );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n6173), .CK(CLK), .Q(n11553), .QN(n8048)
         );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n6172), .CK(CLK), .Q(n11552), .QN(n8065)
         );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n6171), .CK(CLK), .Q(n11551), .QN(n8082)
         );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n6170), .CK(CLK), .Q(n11550), .QN(n8099)
         );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n6169), .CK(CLK), .Q(n11549), .QN(n8116)
         );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n6168), .CK(CLK), .Q(n11548), .QN(n8133)
         );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n6167), .CK(CLK), .Q(n11547), .QN(n8150)
         );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n6166), .CK(CLK), .Q(n11546), .QN(n8167)
         );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n6289), .CK(CLK), .QN(n14329) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n6288), .CK(CLK), .QN(n14330) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n6287), .CK(CLK), .QN(n14331) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n6285), .CK(CLK), .QN(n14332) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n6284), .CK(CLK), .QN(n14333) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n6283), .CK(CLK), .QN(n14334) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n6282), .CK(CLK), .QN(n14335) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n6281), .CK(CLK), .QN(n14336) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n6280), .CK(CLK), .QN(n14337) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n6279), .CK(CLK), .QN(n14338) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n6278), .CK(CLK), .QN(n14339) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n6277), .CK(CLK), .QN(n14340) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n6035), .CK(CLK), .QN(n14341) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n6034), .CK(CLK), .QN(n14342) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n6033), .CK(CLK), .QN(n14343) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n6032), .CK(CLK), .QN(n14344) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n6031), .CK(CLK), .QN(n14345) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n6029), .CK(CLK), .QN(n14346) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n6028), .CK(CLK), .QN(n14347) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n6027), .CK(CLK), .QN(n14348) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n6026), .CK(CLK), .QN(n14349) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n6025), .CK(CLK), .QN(n14350) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n6024), .CK(CLK), .QN(n14351) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n6023), .CK(CLK), .QN(n14352) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n6022), .CK(CLK), .QN(n14353) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n6021), .CK(CLK), .QN(n14354) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n6020), .CK(CLK), .QN(n14355) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n6019), .CK(CLK), .QN(n14356) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n6018), .CK(CLK), .QN(n14357) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n6276), .CK(CLK), .QN(n14358) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n6275), .CK(CLK), .QN(n14359) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n6274), .CK(CLK), .QN(n14360) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n6526), .CK(CLK), .Q(n11586), .QN(n8572)
         );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n6590), .CK(CLK), .Q(n11406), .QN(n8571)
         );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n6654), .CK(CLK), .QN(n14361) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n6718), .CK(CLK), .QN(n14362) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n6782), .CK(CLK), .Q(n11766), .QN(n8570)
         );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n6846), .CK(CLK), .Q(n9948), .QN(n11802)
         );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n6549), .CK(CLK), .Q(n11606), .QN(n8181)
         );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n6548), .CK(CLK), .Q(n11605), .QN(n8198)
         );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n6547), .CK(CLK), .Q(n11604), .QN(n8215)
         );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n6546), .CK(CLK), .Q(n11603), .QN(n8232)
         );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n6545), .CK(CLK), .Q(n11602), .QN(n8249)
         );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n6544), .CK(CLK), .Q(n11601), .QN(n8266)
         );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n6543), .CK(CLK), .Q(n11600), .QN(n8283)
         );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n6542), .CK(CLK), .Q(n11599), .QN(n8300)
         );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n6541), .CK(CLK), .Q(n11598), .QN(n8317)
         );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n6540), .CK(CLK), .Q(n11597), .QN(n8334)
         );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n6539), .CK(CLK), .Q(n11596), .QN(n8351)
         );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n6538), .CK(CLK), .Q(n11595), .QN(n8368)
         );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n6537), .CK(CLK), .Q(n11594), .QN(n8385)
         );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n6536), .CK(CLK), .Q(n11593), .QN(n8402)
         );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n6535), .CK(CLK), .Q(n11592), .QN(n8419)
         );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n6534), .CK(CLK), .Q(n11591), .QN(n8436)
         );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n6533), .CK(CLK), .Q(n11590), .QN(n8453)
         );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n6532), .CK(CLK), .Q(n11764), .QN(n8470)
         );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n6531), .CK(CLK), .Q(n11763), .QN(n8487)
         );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n6530), .CK(CLK), .Q(n11589), .QN(n8504)
         );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n6529), .CK(CLK), .Q(n11588), .QN(n8521)
         );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n6528), .CK(CLK), .Q(n11587), .QN(n8538)
         );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n6527), .CK(CLK), .Q(n11762), .QN(n8555)
         );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n6613), .CK(CLK), .Q(n11426), .QN(n8180)
         );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n6612), .CK(CLK), .Q(n11425), .QN(n8197)
         );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n6611), .CK(CLK), .Q(n11424), .QN(n8214)
         );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n6610), .CK(CLK), .Q(n11423), .QN(n8231)
         );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n6609), .CK(CLK), .Q(n11422), .QN(n8248)
         );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n6608), .CK(CLK), .Q(n11421), .QN(n8265)
         );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n6607), .CK(CLK), .Q(n11420), .QN(n8282)
         );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n6606), .CK(CLK), .Q(n11419), .QN(n8299)
         );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n6605), .CK(CLK), .Q(n11418), .QN(n8316)
         );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n6604), .CK(CLK), .Q(n11417), .QN(n8333)
         );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n6603), .CK(CLK), .Q(n11416), .QN(n8350)
         );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n6602), .CK(CLK), .Q(n11415), .QN(n8367)
         );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n6601), .CK(CLK), .Q(n11414), .QN(n8384)
         );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n6600), .CK(CLK), .Q(n11413), .QN(n8401)
         );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n6599), .CK(CLK), .Q(n11412), .QN(n8418)
         );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n6598), .CK(CLK), .Q(n11411), .QN(n8435)
         );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n6597), .CK(CLK), .Q(n11410), .QN(n8452)
         );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n6596), .CK(CLK), .Q(n11584), .QN(n8469)
         );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n6595), .CK(CLK), .Q(n11583), .QN(n8486)
         );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n6594), .CK(CLK), .Q(n11409), .QN(n8503)
         );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n6593), .CK(CLK), .Q(n11408), .QN(n8520)
         );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n6592), .CK(CLK), .Q(n11407), .QN(n8537)
         );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n6591), .CK(CLK), .Q(n11582), .QN(n8554)
         );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n6677), .CK(CLK), .QN(n14363) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n6676), .CK(CLK), .QN(n14364) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n6675), .CK(CLK), .QN(n14365) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n6674), .CK(CLK), .QN(n14366) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n6673), .CK(CLK), .QN(n14367) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n6672), .CK(CLK), .QN(n14368) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n6671), .CK(CLK), .QN(n14369) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n6670), .CK(CLK), .QN(n14370) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n6669), .CK(CLK), .QN(n14371) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n6668), .CK(CLK), .QN(n14372) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n6667), .CK(CLK), .QN(n14373) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n6666), .CK(CLK), .QN(n14374) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n6665), .CK(CLK), .QN(n14375) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n6664), .CK(CLK), .QN(n14376) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n6663), .CK(CLK), .QN(n14377) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n6662), .CK(CLK), .QN(n14378) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n6661), .CK(CLK), .QN(n14379) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n6660), .CK(CLK), .QN(n14380) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n6659), .CK(CLK), .QN(n14381) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n6658), .CK(CLK), .QN(n14382) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n6657), .CK(CLK), .QN(n14383) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n6656), .CK(CLK), .QN(n14384) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n6655), .CK(CLK), .QN(n14385) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n6741), .CK(CLK), .QN(n14386) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n6740), .CK(CLK), .QN(n14387) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n6739), .CK(CLK), .QN(n14388) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n6738), .CK(CLK), .QN(n14389) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n6737), .CK(CLK), .QN(n14390) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n6736), .CK(CLK), .QN(n14391) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n6735), .CK(CLK), .QN(n14392) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n6734), .CK(CLK), .QN(n14393) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n6733), .CK(CLK), .QN(n14394) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n6732), .CK(CLK), .QN(n14395) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n6731), .CK(CLK), .QN(n14396) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n6730), .CK(CLK), .QN(n14397) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n6729), .CK(CLK), .QN(n14398) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n6728), .CK(CLK), .QN(n14399) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n6727), .CK(CLK), .QN(n14400) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n6726), .CK(CLK), .QN(n14401) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n6725), .CK(CLK), .QN(n14402) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n6724), .CK(CLK), .QN(n14403) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n6723), .CK(CLK), .QN(n14404) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n6722), .CK(CLK), .QN(n14405) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n6721), .CK(CLK), .QN(n14406) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n6720), .CK(CLK), .QN(n14407) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n6719), .CK(CLK), .QN(n14408) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n6805), .CK(CLK), .Q(n9989), .QN(n12056)
         );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n6804), .CK(CLK), .Q(n9990), .QN(n12055)
         );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n6803), .CK(CLK), .Q(n9991), .QN(n12054)
         );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n6802), .CK(CLK), .Q(n9992), .QN(n12053)
         );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n6801), .CK(CLK), .Q(n9993), .QN(n12052)
         );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n6800), .CK(CLK), .Q(n9994), .QN(n12051)
         );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n6799), .CK(CLK), .Q(n9995), .QN(n12050)
         );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n6798), .CK(CLK), .Q(n9996), .QN(n12049)
         );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n6797), .CK(CLK), .Q(n9997), .QN(n12048)
         );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n6796), .CK(CLK), .Q(n9998), .QN(n12047)
         );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n6795), .CK(CLK), .Q(n9999), .QN(n12046)
         );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n6794), .CK(CLK), .Q(n11778), .QN(n8366)
         );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n6793), .CK(CLK), .Q(n11777), .QN(n8383)
         );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n6792), .CK(CLK), .Q(n11776), .QN(n8400)
         );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n6791), .CK(CLK), .Q(n11775), .QN(n8417)
         );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n6790), .CK(CLK), .Q(n11774), .QN(n8434)
         );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n6789), .CK(CLK), .Q(n11773), .QN(n8451)
         );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n6788), .CK(CLK), .Q(n11772), .QN(n8468)
         );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n6787), .CK(CLK), .Q(n11771), .QN(n8485)
         );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n6786), .CK(CLK), .Q(n11770), .QN(n8502)
         );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n6785), .CK(CLK), .Q(n11769), .QN(n8519)
         );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n6784), .CK(CLK), .Q(n11768), .QN(n8536)
         );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n6783), .CK(CLK), .Q(n11767), .QN(n8553)
         );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n6869), .CK(CLK), .Q(n9925), .QN(n11801)
         );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n6868), .CK(CLK), .Q(n9926), .QN(n11800)
         );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n6867), .CK(CLK), .Q(n9927), .QN(n11799)
         );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n6866), .CK(CLK), .Q(n9928), .QN(n11798)
         );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n6865), .CK(CLK), .Q(n9929), .QN(n11797)
         );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n6864), .CK(CLK), .Q(n9930), .QN(n11796)
         );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n6863), .CK(CLK), .Q(n9931), .QN(n11795)
         );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n6862), .CK(CLK), .Q(n9932), .QN(n11794)
         );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n6861), .CK(CLK), .Q(n9933), .QN(n11793)
         );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n6860), .CK(CLK), .Q(n9934), .QN(n11792)
         );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n6859), .CK(CLK), .Q(n9935), .QN(n11791)
         );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n6858), .CK(CLK), .Q(n9936), .QN(n11790)
         );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n6857), .CK(CLK), .Q(n9937), .QN(n11789)
         );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n6856), .CK(CLK), .Q(n9938), .QN(n11788)
         );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n6855), .CK(CLK), .Q(n9939), .QN(n11787)
         );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n6854), .CK(CLK), .Q(n9940), .QN(n11786)
         );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n6853), .CK(CLK), .Q(n9941), .QN(n11785)
         );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n6852), .CK(CLK), .Q(n9942), .QN(n11784)
         );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n6851), .CK(CLK), .Q(n9943), .QN(n11783)
         );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n6850), .CK(CLK), .Q(n9944), .QN(n11782)
         );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n6849), .CK(CLK), .Q(n9945), .QN(n11781)
         );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n6848), .CK(CLK), .Q(n9946), .QN(n11780)
         );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n6847), .CK(CLK), .Q(n9947), .QN(n11779)
         );
  DFF_X1 \REGISTERS_reg[1][60]  ( .D(n6970), .CK(CLK), .QN(n14412) );
  DFF_X1 \REGISTERS_reg[1][59]  ( .D(n6969), .CK(CLK), .QN(n14413) );
  DFF_X1 \REGISTERS_reg[1][58]  ( .D(n6968), .CK(CLK), .QN(n14414) );
  DFF_X1 \REGISTERS_reg[1][57]  ( .D(n6967), .CK(CLK), .QN(n14415) );
  DFF_X1 \REGISTERS_reg[1][56]  ( .D(n6966), .CK(CLK), .QN(n14416) );
  DFF_X1 \REGISTERS_reg[1][55]  ( .D(n6965), .CK(CLK), .QN(n14417) );
  DFF_X1 \REGISTERS_reg[1][54]  ( .D(n6964), .CK(CLK), .QN(n14418) );
  DFF_X1 \REGISTERS_reg[1][53]  ( .D(n6963), .CK(CLK), .QN(n14419) );
  DFF_X1 \REGISTERS_reg[1][52]  ( .D(n6962), .CK(CLK), .QN(n14420) );
  DFF_X1 \REGISTERS_reg[1][51]  ( .D(n6961), .CK(CLK), .QN(n14421) );
  DFF_X1 \REGISTERS_reg[1][50]  ( .D(n6960), .CK(CLK), .QN(n14422) );
  DFF_X1 \REGISTERS_reg[1][49]  ( .D(n6959), .CK(CLK), .QN(n14423) );
  DFF_X1 \REGISTERS_reg[1][48]  ( .D(n6958), .CK(CLK), .QN(n14424) );
  DFF_X1 \REGISTERS_reg[1][47]  ( .D(n6957), .CK(CLK), .QN(n14425) );
  DFF_X1 \REGISTERS_reg[1][46]  ( .D(n6956), .CK(CLK), .QN(n14426) );
  DFF_X1 \REGISTERS_reg[1][45]  ( .D(n6955), .CK(CLK), .QN(n14427) );
  DFF_X1 \REGISTERS_reg[1][44]  ( .D(n6954), .CK(CLK), .QN(n14428) );
  DFF_X1 \REGISTERS_reg[1][43]  ( .D(n6953), .CK(CLK), .QN(n14429) );
  DFF_X1 \REGISTERS_reg[1][42]  ( .D(n6952), .CK(CLK), .QN(n14430) );
  DFF_X1 \REGISTERS_reg[1][41]  ( .D(n6951), .CK(CLK), .QN(n14431) );
  DFF_X1 \REGISTERS_reg[1][40]  ( .D(n6950), .CK(CLK), .QN(n14432) );
  DFF_X1 \REGISTERS_reg[0][62]  ( .D(n7036), .CK(CLK), .QN(n14433) );
  DFF_X1 \REGISTERS_reg[0][61]  ( .D(n7035), .CK(CLK), .QN(n14434) );
  DFF_X1 \REGISTERS_reg[0][60]  ( .D(n7034), .CK(CLK), .QN(n14435) );
  DFF_X1 \REGISTERS_reg[0][59]  ( .D(n7033), .CK(CLK), .QN(n14436) );
  DFF_X1 \REGISTERS_reg[0][58]  ( .D(n7032), .CK(CLK), .QN(n14437) );
  DFF_X1 \REGISTERS_reg[0][57]  ( .D(n7031), .CK(CLK), .QN(n14438) );
  DFF_X1 \REGISTERS_reg[0][56]  ( .D(n7030), .CK(CLK), .QN(n14439) );
  DFF_X1 \REGISTERS_reg[0][55]  ( .D(n7029), .CK(CLK), .QN(n14440) );
  DFF_X1 \REGISTERS_reg[0][45]  ( .D(n7019), .CK(CLK), .QN(n14441) );
  DFF_X1 \REGISTERS_reg[0][44]  ( .D(n7018), .CK(CLK), .QN(n14442) );
  DFF_X1 \REGISTERS_reg[0][43]  ( .D(n7017), .CK(CLK), .QN(n14443) );
  DFF_X1 \REGISTERS_reg[0][42]  ( .D(n7016), .CK(CLK), .QN(n14444) );
  DFF_X1 \REGISTERS_reg[0][41]  ( .D(n7015), .CK(CLK), .QN(n14445) );
  DFF_X1 \REGISTERS_reg[0][40]  ( .D(n7014), .CK(CLK), .QN(n14446) );
  DFF_X1 \REGISTERS_reg[0][39]  ( .D(n7013), .CK(CLK), .QN(n14447) );
  DFF_X1 \REGISTERS_reg[0][38]  ( .D(n7012), .CK(CLK), .QN(n14448) );
  DFF_X1 \REGISTERS_reg[0][37]  ( .D(n7011), .CK(CLK), .QN(n14449) );
  DFF_X1 \REGISTERS_reg[0][36]  ( .D(n7010), .CK(CLK), .QN(n14450) );
  DFF_X1 \REGISTERS_reg[0][35]  ( .D(n7009), .CK(CLK), .QN(n14451) );
  DFF_X1 \REGISTERS_reg[0][34]  ( .D(n7008), .CK(CLK), .QN(n14452) );
  DFF_X1 \REGISTERS_reg[0][33]  ( .D(n7007), .CK(CLK), .QN(n14453) );
  DFF_X1 \REGISTERS_reg[0][32]  ( .D(n7006), .CK(CLK), .QN(n14454) );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n7005), .CK(CLK), .QN(n14455) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n7004), .CK(CLK), .QN(n14456) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n6421), .CK(CLK), .Q(n11485), .QN(n8182)
         );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n6420), .CK(CLK), .Q(n11484), .QN(n8199)
         );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n6419), .CK(CLK), .Q(n11483), .QN(n8216)
         );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n6418), .CK(CLK), .Q(n11482), .QN(n8233)
         );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n6417), .CK(CLK), .Q(n11481), .QN(n8250)
         );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n6416), .CK(CLK), .Q(n11480), .QN(n8267)
         );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n6415), .CK(CLK), .Q(n11479), .QN(n8284)
         );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n6414), .CK(CLK), .Q(n11478), .QN(n8301)
         );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n6413), .CK(CLK), .Q(n11477), .QN(n8318)
         );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n6412), .CK(CLK), .Q(n11476), .QN(n8335)
         );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n6411), .CK(CLK), .Q(n11475), .QN(n8352)
         );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n6410), .CK(CLK), .Q(n11474), .QN(n8369)
         );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n6409), .CK(CLK), .Q(n11473), .QN(n8386)
         );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n6408), .CK(CLK), .Q(n11472), .QN(n8403)
         );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n6407), .CK(CLK), .Q(n11471), .QN(n8420)
         );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n6406), .CK(CLK), .Q(n11470), .QN(n8437)
         );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n6405), .CK(CLK), .Q(n11469), .QN(n8454)
         );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n6404), .CK(CLK), .Q(n11468), .QN(n8471)
         );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n6403), .CK(CLK), .Q(n11467), .QN(n8488)
         );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n6402), .CK(CLK), .Q(n11466), .QN(n8505)
         );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n6401), .CK(CLK), .Q(n11465), .QN(n8522)
         );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n6400), .CK(CLK), .Q(n11464), .QN(n8539)
         );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n6399), .CK(CLK), .Q(n11463), .QN(n8556)
         );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n6398), .CK(CLK), .Q(n11462), .QN(n8573)
         );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n6485), .CK(CLK), .Q(n11665), .QN(n8183)
         );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n6484), .CK(CLK), .Q(n11664), .QN(n8200)
         );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n6483), .CK(CLK), .Q(n11663), .QN(n8217)
         );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n6482), .CK(CLK), .Q(n11662), .QN(n8234)
         );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n6481), .CK(CLK), .Q(n11661), .QN(n8251)
         );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n6480), .CK(CLK), .Q(n11660), .QN(n8268)
         );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n6479), .CK(CLK), .Q(n11659), .QN(n8285)
         );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n6478), .CK(CLK), .Q(n11658), .QN(n8302)
         );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n6477), .CK(CLK), .Q(n11657), .QN(n8319)
         );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n6476), .CK(CLK), .Q(n11656), .QN(n8336)
         );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n6475), .CK(CLK), .Q(n11655), .QN(n8353)
         );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n6474), .CK(CLK), .Q(n11654), .QN(n8370)
         );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n6473), .CK(CLK), .Q(n11653), .QN(n8387)
         );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n6472), .CK(CLK), .Q(n11652), .QN(n8404)
         );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n6471), .CK(CLK), .Q(n11651), .QN(n8421)
         );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n6470), .CK(CLK), .Q(n11650), .QN(n8438)
         );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n6469), .CK(CLK), .Q(n11649), .QN(n8455)
         );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n6468), .CK(CLK), .Q(n11648), .QN(n8472)
         );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n6467), .CK(CLK), .Q(n11647), .QN(n8489)
         );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n6466), .CK(CLK), .Q(n11646), .QN(n8506)
         );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n6465), .CK(CLK), .Q(n11645), .QN(n8523)
         );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n6464), .CK(CLK), .Q(n11644), .QN(n8540)
         );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n6463), .CK(CLK), .Q(n11643), .QN(n8557)
         );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n6462), .CK(CLK), .Q(n11642), .QN(n8574)
         );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n6229), .CK(CLK), .Q(n11725), .QN(n8185)
         );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n6228), .CK(CLK), .Q(n11724), .QN(n8202)
         );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n6227), .CK(CLK), .Q(n11723), .QN(n8219)
         );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n6226), .CK(CLK), .Q(n11722), .QN(n8236)
         );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n6225), .CK(CLK), .Q(n11721), .QN(n8253)
         );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n6224), .CK(CLK), .Q(n11720), .QN(n8270)
         );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n6223), .CK(CLK), .Q(n11719), .QN(n8287)
         );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n6222), .CK(CLK), .Q(n11718), .QN(n8304)
         );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n6221), .CK(CLK), .Q(n11717), .QN(n8321)
         );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n6220), .CK(CLK), .Q(n11716), .QN(n8338)
         );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n6219), .CK(CLK), .Q(n11715), .QN(n8355)
         );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n6218), .CK(CLK), .Q(n11714), .QN(n8372)
         );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n6217), .CK(CLK), .Q(n11713), .QN(n8389)
         );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n6216), .CK(CLK), .Q(n11712), .QN(n8406)
         );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n6215), .CK(CLK), .Q(n11711), .QN(n8423)
         );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n6214), .CK(CLK), .Q(n11710), .QN(n8440)
         );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n6213), .CK(CLK), .Q(n11709), .QN(n8457)
         );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n6212), .CK(CLK), .Q(n11708), .QN(n8474)
         );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n6211), .CK(CLK), .Q(n11707), .QN(n8491)
         );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n6210), .CK(CLK), .Q(n11706), .QN(n8508)
         );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n6209), .CK(CLK), .Q(n11705), .QN(n8525)
         );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n6208), .CK(CLK), .Q(n11704), .QN(n8542)
         );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n6207), .CK(CLK), .Q(n11703), .QN(n8559)
         );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n6206), .CK(CLK), .Q(n11702), .QN(n8576)
         );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n6165), .CK(CLK), .Q(n11545), .QN(n8184)
         );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n6164), .CK(CLK), .Q(n11544), .QN(n8201)
         );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n6163), .CK(CLK), .Q(n11543), .QN(n8218)
         );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n6162), .CK(CLK), .Q(n11542), .QN(n8235)
         );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n6161), .CK(CLK), .Q(n11541), .QN(n8252)
         );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n6160), .CK(CLK), .Q(n11540), .QN(n8269)
         );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n6159), .CK(CLK), .Q(n11539), .QN(n8286)
         );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n6158), .CK(CLK), .Q(n11538), .QN(n8303)
         );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n6157), .CK(CLK), .Q(n11537), .QN(n8320)
         );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n6156), .CK(CLK), .Q(n11536), .QN(n8337)
         );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n6155), .CK(CLK), .Q(n11535), .QN(n8354)
         );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n6154), .CK(CLK), .Q(n11534), .QN(n8371)
         );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n6153), .CK(CLK), .Q(n11533), .QN(n8388)
         );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n6152), .CK(CLK), .Q(n11532), .QN(n8405)
         );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n6151), .CK(CLK), .Q(n11531), .QN(n8422)
         );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n6150), .CK(CLK), .Q(n11530), .QN(n8439)
         );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n6149), .CK(CLK), .Q(n11529), .QN(n8456)
         );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n6148), .CK(CLK), .Q(n11528), .QN(n8473)
         );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n6147), .CK(CLK), .Q(n11527), .QN(n8490)
         );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n6146), .CK(CLK), .Q(n11526), .QN(n8507)
         );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n6145), .CK(CLK), .Q(n11525), .QN(n8524)
         );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n6144), .CK(CLK), .Q(n11524), .QN(n8541)
         );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n6143), .CK(CLK), .Q(n11523), .QN(n8558)
         );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n6142), .CK(CLK), .Q(n11522), .QN(n8575)
         );
  DFF_X1 \REGISTERS_reg[11][42]  ( .D(n6312), .CK(CLK), .QN(n14457) );
  DFF_X1 \REGISTERS_reg[11][41]  ( .D(n6311), .CK(CLK), .QN(n14458) );
  DFF_X1 \REGISTERS_reg[11][40]  ( .D(n6310), .CK(CLK), .QN(n14459) );
  DFF_X1 \REGISTERS_reg[11][39]  ( .D(n6309), .CK(CLK), .QN(n14460) );
  NAND3_X1 U6638 ( .A1(n13383), .A2(n13382), .A3(n1922), .ZN(n1906) );
  NAND3_X1 U6640 ( .A1(n1922), .A2(n13383), .A3(ADD_WR[4]), .ZN(n1933) );
  NAND3_X1 U6641 ( .A1(n13385), .A2(n13384), .A3(n13386), .ZN(n1907) );
  NAND3_X1 U6642 ( .A1(n13385), .A2(n13384), .A3(ADD_WR[0]), .ZN(n1909) );
  NAND3_X1 U6643 ( .A1(n13386), .A2(n13384), .A3(ADD_WR[1]), .ZN(n1911) );
  NAND3_X1 U6644 ( .A1(ADD_WR[0]), .A2(n13384), .A3(ADD_WR[1]), .ZN(n1913) );
  NAND3_X1 U6645 ( .A1(n13386), .A2(n13385), .A3(ADD_WR[2]), .ZN(n1915) );
  NAND3_X1 U6646 ( .A1(ADD_WR[0]), .A2(n13385), .A3(ADD_WR[2]), .ZN(n1917) );
  NAND3_X1 U6647 ( .A1(ADD_WR[1]), .A2(n13386), .A3(ADD_WR[2]), .ZN(n1919) );
  NAND3_X1 U6649 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n1921)
         );
  DFF_X1 \REGISTERS_reg[25][63]  ( .D(n5437), .CK(CLK), .QN(n13731) );
  DFF_X1 \REGISTERS_reg[25][62]  ( .D(n5436), .CK(CLK), .QN(n13732) );
  DFF_X1 \REGISTERS_reg[25][61]  ( .D(n5435), .CK(CLK), .QN(n13733) );
  DFF_X1 \REGISTERS_reg[25][60]  ( .D(n5434), .CK(CLK), .QN(n13734) );
  DFF_X1 \REGISTERS_reg[24][63]  ( .D(n5501), .CK(CLK), .QN(n13667) );
  DFF_X1 \REGISTERS_reg[24][62]  ( .D(n5500), .CK(CLK), .QN(n13668) );
  DFF_X1 \REGISTERS_reg[24][61]  ( .D(n5499), .CK(CLK), .QN(n13669) );
  DFF_X1 \REGISTERS_reg[24][60]  ( .D(n5498), .CK(CLK), .QN(n13670) );
  DFF_X1 \REGISTERS_reg[28][63]  ( .D(n5245), .CK(CLK), .QN(n13747) );
  DFF_X1 \REGISTERS_reg[28][62]  ( .D(n5244), .CK(CLK), .QN(n13748) );
  DFF_X1 \REGISTERS_reg[28][61]  ( .D(n5243), .CK(CLK), .QN(n13749) );
  DFF_X1 \REGISTERS_reg[28][60]  ( .D(n5242), .CK(CLK), .QN(n13750) );
  DFF_X1 \REGISTERS_reg[29][63]  ( .D(n5181), .CK(CLK), .QN(n14083) );
  DFF_X1 \REGISTERS_reg[29][62]  ( .D(n5180), .CK(CLK), .QN(n14084) );
  DFF_X1 \REGISTERS_reg[29][61]  ( .D(n5179), .CK(CLK), .QN(n14085) );
  DFF_X1 \REGISTERS_reg[29][60]  ( .D(n5178), .CK(CLK), .QN(n14086) );
  DFF_X1 \REGISTERS_reg[23][63]  ( .D(n5565), .CK(CLK), .Q(n4511), .QN(n13663)
         );
  DFF_X1 \REGISTERS_reg[23][62]  ( .D(n5564), .CK(CLK), .Q(n4509), .QN(n13664)
         );
  DFF_X1 \REGISTERS_reg[23][61]  ( .D(n5563), .CK(CLK), .Q(n4507), .QN(n13665)
         );
  DFF_X1 \REGISTERS_reg[23][60]  ( .D(n5562), .CK(CLK), .Q(n4505), .QN(n13666)
         );
  DFF_X1 \REGISTERS_reg[22][63]  ( .D(n5629), .CK(CLK), .Q(n4510), .QN(n13659)
         );
  DFF_X1 \REGISTERS_reg[22][62]  ( .D(n5628), .CK(CLK), .Q(n4508), .QN(n13660)
         );
  DFF_X1 \REGISTERS_reg[22][61]  ( .D(n5627), .CK(CLK), .Q(n4506), .QN(n13661)
         );
  DFF_X1 \REGISTERS_reg[22][60]  ( .D(n5626), .CK(CLK), .Q(n4504), .QN(n13662)
         );
  DFF_X1 \REGISTERS_reg[19][63]  ( .D(n5821), .CK(CLK), .Q(n4479), .QN(n13655)
         );
  DFF_X1 \REGISTERS_reg[19][62]  ( .D(n5820), .CK(CLK), .Q(n4477), .QN(n13656)
         );
  DFF_X1 \REGISTERS_reg[19][61]  ( .D(n5819), .CK(CLK), .Q(n4475), .QN(n13657)
         );
  DFF_X1 \REGISTERS_reg[19][60]  ( .D(n5818), .CK(CLK), .Q(n4473), .QN(n13658)
         );
  DFF_X1 \REGISTERS_reg[18][63]  ( .D(n5885), .CK(CLK), .Q(n4478), .QN(n13651)
         );
  DFF_X1 \REGISTERS_reg[18][62]  ( .D(n5884), .CK(CLK), .Q(n4476), .QN(n13652)
         );
  DFF_X1 \REGISTERS_reg[18][61]  ( .D(n5883), .CK(CLK), .Q(n4474), .QN(n13653)
         );
  DFF_X1 \REGISTERS_reg[18][60]  ( .D(n5882), .CK(CLK), .Q(n4472), .QN(n13654)
         );
  DFF_X1 \REGISTERS_reg[3][63]  ( .D(n6845), .CK(CLK), .Q(n9949), .QN(n13848)
         );
  DFF_X1 \REGISTERS_reg[10][63]  ( .D(n6397), .CK(CLK), .QN(n13431) );
  DFF_X1 \REGISTERS_reg[10][62]  ( .D(n6396), .CK(CLK), .QN(n13432) );
  DFF_X1 \REGISTERS_reg[10][61]  ( .D(n6395), .CK(CLK), .QN(n13433) );
  DFF_X1 \REGISTERS_reg[10][60]  ( .D(n6394), .CK(CLK), .QN(n13434) );
  DFF_X1 \REGISTERS_reg[11][63]  ( .D(n6333), .CK(CLK), .QN(n13495) );
  DFF_X1 \REGISTERS_reg[11][62]  ( .D(n6332), .CK(CLK), .QN(n13496) );
  DFF_X1 \REGISTERS_reg[11][61]  ( .D(n6331), .CK(CLK), .QN(n13497) );
  DFF_X1 \REGISTERS_reg[11][60]  ( .D(n6330), .CK(CLK), .QN(n13498) );
  DFF_X1 \REGISTERS_reg[15][63]  ( .D(n6077), .CK(CLK), .QN(n13604) );
  DFF_X1 \REGISTERS_reg[15][62]  ( .D(n6076), .CK(CLK), .QN(n13605) );
  DFF_X1 \REGISTERS_reg[15][61]  ( .D(n6075), .CK(CLK), .QN(n13606) );
  DFF_X1 \REGISTERS_reg[15][60]  ( .D(n6074), .CK(CLK), .QN(n13607) );
  DFF_X1 \REGISTERS_reg[14][63]  ( .D(n6141), .CK(CLK), .QN(n13540) );
  DFF_X1 \REGISTERS_reg[14][62]  ( .D(n6140), .CK(CLK), .QN(n13541) );
  DFF_X1 \REGISTERS_reg[14][61]  ( .D(n6139), .CK(CLK), .QN(n13542) );
  DFF_X1 \REGISTERS_reg[14][60]  ( .D(n6138), .CK(CLK), .QN(n13543) );
  DFF_X1 \REGISTERS_reg[5][63]  ( .D(n6717), .CK(CLK), .QN(n13840) );
  DFF_X1 \REGISTERS_reg[5][62]  ( .D(n6716), .CK(CLK), .QN(n13841) );
  DFF_X1 \REGISTERS_reg[5][61]  ( .D(n6715), .CK(CLK), .QN(n13842) );
  DFF_X1 \REGISTERS_reg[5][60]  ( .D(n6714), .CK(CLK), .QN(n13843) );
  DFF_X1 \REGISTERS_reg[4][63]  ( .D(n6781), .CK(CLK), .QN(n13844) );
  DFF_X1 \REGISTERS_reg[4][62]  ( .D(n6780), .CK(CLK), .QN(n13845) );
  DFF_X1 \REGISTERS_reg[4][61]  ( .D(n6779), .CK(CLK), .QN(n13846) );
  DFF_X1 \REGISTERS_reg[4][60]  ( .D(n6778), .CK(CLK), .QN(n13847) );
  DFF_X1 \REGISTERS_reg[2][63]  ( .D(n6909), .CK(CLK), .Q(n9885), .QN(n13849)
         );
  DFF_X1 \REGISTERS_reg[2][62]  ( .D(n6908), .CK(CLK), .Q(n9886), .QN(n13850)
         );
  DFF_X1 \REGISTERS_reg[2][61]  ( .D(n6907), .CK(CLK), .Q(n9887), .QN(n13851)
         );
  DFF_X1 \REGISTERS_reg[2][60]  ( .D(n6906), .CK(CLK), .Q(n9888), .QN(n13852)
         );
  DFF_X1 \REGISTERS_reg[1][63]  ( .D(n6973), .CK(CLK), .QN(n14409) );
  DFF_X1 \REGISTERS_reg[1][62]  ( .D(n6972), .CK(CLK), .QN(n14410) );
  DFF_X1 \REGISTERS_reg[1][61]  ( .D(n6971), .CK(CLK), .QN(n14411) );
  DFF_X1 \REGISTERS_reg[26][63]  ( .D(n5373), .CK(CLK), .Q(n13816), .QN(n4848)
         );
  DFF_X1 \REGISTERS_reg[26][62]  ( .D(n5372), .CK(CLK), .Q(n13817), .QN(n7109)
         );
  DFF_X1 \REGISTERS_reg[26][61]  ( .D(n5371), .CK(CLK), .Q(n13818), .QN(n7126)
         );
  DFF_X1 \REGISTERS_reg[26][60]  ( .D(n5370), .CK(CLK), .Q(n13819), .QN(n7143)
         );
  DFF_X1 \REGISTERS_reg[27][63]  ( .D(n5309), .CK(CLK), .Q(n13820), .QN(n4847)
         );
  DFF_X1 \REGISTERS_reg[27][62]  ( .D(n5308), .CK(CLK), .Q(n13821), .QN(n7108)
         );
  DFF_X1 \REGISTERS_reg[27][61]  ( .D(n5307), .CK(CLK), .Q(n13822), .QN(n7125)
         );
  DFF_X1 \REGISTERS_reg[27][60]  ( .D(n5306), .CK(CLK), .Q(n13823), .QN(n7142)
         );
  DFF_X1 \REGISTERS_reg[30][63]  ( .D(n5117), .CK(CLK), .Q(n13824), .QN(n4850)
         );
  DFF_X1 \REGISTERS_reg[30][62]  ( .D(n5116), .CK(CLK), .Q(n13825), .QN(n7111)
         );
  DFF_X1 \REGISTERS_reg[30][61]  ( .D(n5115), .CK(CLK), .Q(n13826), .QN(n7128)
         );
  DFF_X1 \REGISTERS_reg[30][60]  ( .D(n5114), .CK(CLK), .Q(n13827), .QN(n7145)
         );
  DFF_X1 \REGISTERS_reg[31][63]  ( .D(n5053), .CK(CLK), .Q(n14156), .QN(n4849)
         );
  DFF_X1 \REGISTERS_reg[31][62]  ( .D(n5052), .CK(CLK), .Q(n14157), .QN(n7110)
         );
  DFF_X1 \REGISTERS_reg[31][61]  ( .D(n5051), .CK(CLK), .Q(n14158), .QN(n7127)
         );
  DFF_X1 \REGISTERS_reg[31][60]  ( .D(n5050), .CK(CLK), .Q(n14159), .QN(n7144)
         );
  DFF_X1 \REGISTERS_reg[21][63]  ( .D(n5693), .CK(CLK), .QN(n4845) );
  DFF_X1 \REGISTERS_reg[21][62]  ( .D(n5692), .CK(CLK), .QN(n7106) );
  DFF_X1 \REGISTERS_reg[21][61]  ( .D(n5691), .CK(CLK), .QN(n7123) );
  DFF_X1 \REGISTERS_reg[21][60]  ( .D(n5690), .CK(CLK), .QN(n7140) );
  DFF_X1 \REGISTERS_reg[20][63]  ( .D(n5757), .CK(CLK), .QN(n4846) );
  DFF_X1 \REGISTERS_reg[20][62]  ( .D(n5756), .CK(CLK), .QN(n7107) );
  DFF_X1 \REGISTERS_reg[20][61]  ( .D(n5755), .CK(CLK), .QN(n7124) );
  DFF_X1 \REGISTERS_reg[20][60]  ( .D(n5754), .CK(CLK), .QN(n7141) );
  DFF_X1 \REGISTERS_reg[17][63]  ( .D(n5949), .CK(CLK), .QN(n4843) );
  DFF_X1 \REGISTERS_reg[17][62]  ( .D(n5948), .CK(CLK), .QN(n4860) );
  DFF_X1 \REGISTERS_reg[17][61]  ( .D(n5947), .CK(CLK), .QN(n7121) );
  DFF_X1 \REGISTERS_reg[17][60]  ( .D(n5946), .CK(CLK), .QN(n7138) );
  DFF_X1 \REGISTERS_reg[16][63]  ( .D(n6013), .CK(CLK), .QN(n4844) );
  DFF_X1 \REGISTERS_reg[16][62]  ( .D(n6012), .CK(CLK), .QN(n4861) );
  DFF_X1 \REGISTERS_reg[16][61]  ( .D(n6011), .CK(CLK), .QN(n7122) );
  DFF_X1 \REGISTERS_reg[16][60]  ( .D(n6010), .CK(CLK), .QN(n7139) );
  DFF_X1 \REGISTERS_reg[9][63]  ( .D(n6461), .CK(CLK), .Q(n13853), .QN(n4839)
         );
  DFF_X1 \REGISTERS_reg[9][62]  ( .D(n6460), .CK(CLK), .Q(n13854), .QN(n4856)
         );
  DFF_X1 \REGISTERS_reg[9][61]  ( .D(n6459), .CK(CLK), .Q(n13855), .QN(n7117)
         );
  DFF_X1 \REGISTERS_reg[9][60]  ( .D(n6458), .CK(CLK), .Q(n13856), .QN(n7134)
         );
  DFF_X1 \REGISTERS_reg[8][63]  ( .D(n6525), .CK(CLK), .Q(n13857), .QN(n4840)
         );
  DFF_X1 \REGISTERS_reg[8][62]  ( .D(n6524), .CK(CLK), .Q(n13858), .QN(n4857)
         );
  DFF_X1 \REGISTERS_reg[8][61]  ( .D(n6523), .CK(CLK), .Q(n13859), .QN(n7118)
         );
  DFF_X1 \REGISTERS_reg[8][60]  ( .D(n6522), .CK(CLK), .Q(n13860), .QN(n7135)
         );
  DFF_X1 \REGISTERS_reg[13][63]  ( .D(n6205), .CK(CLK), .Q(n13865), .QN(n4841)
         );
  DFF_X1 \REGISTERS_reg[13][62]  ( .D(n6204), .CK(CLK), .Q(n13866), .QN(n4858)
         );
  DFF_X1 \REGISTERS_reg[13][61]  ( .D(n6203), .CK(CLK), .Q(n13867), .QN(n7119)
         );
  DFF_X1 \REGISTERS_reg[13][60]  ( .D(n6202), .CK(CLK), .Q(n13868), .QN(n7136)
         );
  DFF_X1 \REGISTERS_reg[12][63]  ( .D(n6269), .CK(CLK), .Q(n13861), .QN(n4842)
         );
  DFF_X1 \REGISTERS_reg[12][62]  ( .D(n6268), .CK(CLK), .Q(n13862), .QN(n4859)
         );
  DFF_X1 \REGISTERS_reg[12][61]  ( .D(n6267), .CK(CLK), .Q(n13863), .QN(n7120)
         );
  DFF_X1 \REGISTERS_reg[12][60]  ( .D(n6266), .CK(CLK), .Q(n13864), .QN(n7137)
         );
  DFF_X1 \REGISTERS_reg[7][63]  ( .D(n6589), .CK(CLK), .Q(n13832), .QN(n4838)
         );
  DFF_X1 \REGISTERS_reg[7][62]  ( .D(n6588), .CK(CLK), .Q(n13833), .QN(n4855)
         );
  DFF_X1 \REGISTERS_reg[7][61]  ( .D(n6587), .CK(CLK), .Q(n13834), .QN(n7116)
         );
  DFF_X1 \REGISTERS_reg[7][60]  ( .D(n6586), .CK(CLK), .Q(n13835), .QN(n7133)
         );
  DFF_X1 \REGISTERS_reg[6][63]  ( .D(n6653), .CK(CLK), .Q(n13836), .QN(n4837)
         );
  DFF_X1 \REGISTERS_reg[6][62]  ( .D(n6652), .CK(CLK), .Q(n13837), .QN(n4854)
         );
  DFF_X1 \REGISTERS_reg[6][61]  ( .D(n6651), .CK(CLK), .Q(n13838), .QN(n7115)
         );
  DFF_X1 \REGISTERS_reg[6][60]  ( .D(n6650), .CK(CLK), .Q(n13839), .QN(n7132)
         );
  DFF_X1 \REGISTERS_reg[26][59]  ( .D(n5369), .CK(CLK), .Q(n13893), .QN(n7240)
         );
  DFF_X1 \REGISTERS_reg[26][58]  ( .D(n5368), .CK(CLK), .Q(n13894), .QN(n7257)
         );
  DFF_X1 \REGISTERS_reg[26][57]  ( .D(n5367), .CK(CLK), .Q(n13895), .QN(n7274)
         );
  DFF_X1 \REGISTERS_reg[26][56]  ( .D(n5366), .CK(CLK), .Q(n13896), .QN(n7373)
         );
  DFF_X1 \REGISTERS_reg[26][55]  ( .D(n5365), .CK(CLK), .Q(n13897), .QN(n7390)
         );
  DFF_X1 \REGISTERS_reg[26][54]  ( .D(n5364), .CK(CLK), .Q(n13898), .QN(n7492)
         );
  DFF_X1 \REGISTERS_reg[26][53]  ( .D(n5363), .CK(CLK), .Q(n13899), .QN(n7509)
         );
  DFF_X1 \REGISTERS_reg[26][52]  ( .D(n5362), .CK(CLK), .Q(n13900), .QN(n7526)
         );
  DFF_X1 \REGISTERS_reg[26][51]  ( .D(n5361), .CK(CLK), .Q(n13901), .QN(n7630)
         );
  DFF_X1 \REGISTERS_reg[26][50]  ( .D(n5360), .CK(CLK), .Q(n13902), .QN(n7647)
         );
  DFF_X1 \REGISTERS_reg[26][49]  ( .D(n5359), .CK(CLK), .Q(n13903), .QN(n7749)
         );
  DFF_X1 \REGISTERS_reg[26][48]  ( .D(n5358), .CK(CLK), .Q(n13904), .QN(n7766)
         );
  DFF_X1 \REGISTERS_reg[26][47]  ( .D(n5357), .CK(CLK), .Q(n13905), .QN(n7783)
         );
  DFF_X1 \REGISTERS_reg[26][46]  ( .D(n5356), .CK(CLK), .Q(n13906), .QN(n7800)
         );
  DFF_X1 \REGISTERS_reg[26][45]  ( .D(n5355), .CK(CLK), .Q(n13907), .QN(n7817)
         );
  DFF_X1 \REGISTERS_reg[26][44]  ( .D(n5354), .CK(CLK), .Q(n13908), .QN(n7834)
         );
  DFF_X1 \REGISTERS_reg[26][43]  ( .D(n5353), .CK(CLK), .Q(n13909), .QN(n7851)
         );
  DFF_X1 \REGISTERS_reg[26][42]  ( .D(n5352), .CK(CLK), .Q(n13910), .QN(n7868)
         );
  DFF_X1 \REGISTERS_reg[26][41]  ( .D(n5351), .CK(CLK), .Q(n13911), .QN(n7885)
         );
  DFF_X1 \REGISTERS_reg[26][40]  ( .D(n5350), .CK(CLK), .Q(n13912), .QN(n7902)
         );
  DFF_X1 \REGISTERS_reg[26][39]  ( .D(n5349), .CK(CLK), .Q(n13913), .QN(n7919)
         );
  DFF_X1 \REGISTERS_reg[26][38]  ( .D(n5348), .CK(CLK), .Q(n13914), .QN(n7936)
         );
  DFF_X1 \REGISTERS_reg[26][37]  ( .D(n5347), .CK(CLK), .Q(n13915), .QN(n7953)
         );
  DFF_X1 \REGISTERS_reg[26][36]  ( .D(n5346), .CK(CLK), .Q(n13916), .QN(n7970)
         );
  DFF_X1 \REGISTERS_reg[26][35]  ( .D(n5345), .CK(CLK), .Q(n13917), .QN(n7987)
         );
  DFF_X1 \REGISTERS_reg[26][34]  ( .D(n5344), .CK(CLK), .Q(n13918), .QN(n8004)
         );
  DFF_X1 \REGISTERS_reg[26][33]  ( .D(n5343), .CK(CLK), .Q(n13919), .QN(n8021)
         );
  DFF_X1 \REGISTERS_reg[26][32]  ( .D(n5342), .CK(CLK), .Q(n13920), .QN(n8038)
         );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n5341), .CK(CLK), .Q(n13921), .QN(n8055)
         );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n5340), .CK(CLK), .Q(n13922), .QN(n8072)
         );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n5339), .CK(CLK), .Q(n13923), .QN(n8089)
         );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n5338), .CK(CLK), .Q(n13924), .QN(n8106)
         );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n5337), .CK(CLK), .Q(n13925), .QN(n8123)
         );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n5336), .CK(CLK), .Q(n13926), .QN(n8140)
         );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n5335), .CK(CLK), .Q(n13927), .QN(n8157)
         );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n5334), .CK(CLK), .Q(n13928), .QN(n8174)
         );
  DFF_X1 \REGISTERS_reg[27][59]  ( .D(n5305), .CK(CLK), .Q(n13953), .QN(n7239)
         );
  DFF_X1 \REGISTERS_reg[27][58]  ( .D(n5304), .CK(CLK), .Q(n13954), .QN(n7256)
         );
  DFF_X1 \REGISTERS_reg[27][57]  ( .D(n5303), .CK(CLK), .Q(n13955), .QN(n7273)
         );
  DFF_X1 \REGISTERS_reg[27][56]  ( .D(n5302), .CK(CLK), .Q(n13956), .QN(n7372)
         );
  DFF_X1 \REGISTERS_reg[27][55]  ( .D(n5301), .CK(CLK), .Q(n13957), .QN(n7389)
         );
  DFF_X1 \REGISTERS_reg[27][54]  ( .D(n5300), .CK(CLK), .Q(n13958), .QN(n7491)
         );
  DFF_X1 \REGISTERS_reg[27][53]  ( .D(n5299), .CK(CLK), .Q(n13959), .QN(n7508)
         );
  DFF_X1 \REGISTERS_reg[27][52]  ( .D(n5298), .CK(CLK), .Q(n13960), .QN(n7525)
         );
  DFF_X1 \REGISTERS_reg[27][51]  ( .D(n5297), .CK(CLK), .Q(n13961), .QN(n7629)
         );
  DFF_X1 \REGISTERS_reg[27][50]  ( .D(n5296), .CK(CLK), .Q(n13962), .QN(n7646)
         );
  DFF_X1 \REGISTERS_reg[27][49]  ( .D(n5295), .CK(CLK), .Q(n13963), .QN(n7748)
         );
  DFF_X1 \REGISTERS_reg[27][48]  ( .D(n5294), .CK(CLK), .Q(n13964), .QN(n7765)
         );
  DFF_X1 \REGISTERS_reg[27][47]  ( .D(n5293), .CK(CLK), .Q(n13965), .QN(n7782)
         );
  DFF_X1 \REGISTERS_reg[27][46]  ( .D(n5292), .CK(CLK), .Q(n13966), .QN(n7799)
         );
  DFF_X1 \REGISTERS_reg[27][45]  ( .D(n5291), .CK(CLK), .Q(n13967), .QN(n7816)
         );
  DFF_X1 \REGISTERS_reg[27][44]  ( .D(n5290), .CK(CLK), .Q(n13968), .QN(n7833)
         );
  DFF_X1 \REGISTERS_reg[27][43]  ( .D(n5289), .CK(CLK), .Q(n13969), .QN(n7850)
         );
  DFF_X1 \REGISTERS_reg[27][42]  ( .D(n5288), .CK(CLK), .Q(n13970), .QN(n7867)
         );
  DFF_X1 \REGISTERS_reg[27][41]  ( .D(n5287), .CK(CLK), .Q(n13971), .QN(n7884)
         );
  DFF_X1 \REGISTERS_reg[27][40]  ( .D(n5286), .CK(CLK), .Q(n13972), .QN(n7901)
         );
  DFF_X1 \REGISTERS_reg[27][39]  ( .D(n5285), .CK(CLK), .Q(n13973), .QN(n7918)
         );
  DFF_X1 \REGISTERS_reg[27][38]  ( .D(n5284), .CK(CLK), .Q(n13974), .QN(n7935)
         );
  DFF_X1 \REGISTERS_reg[27][37]  ( .D(n5283), .CK(CLK), .Q(n13975), .QN(n7952)
         );
  DFF_X1 \REGISTERS_reg[27][36]  ( .D(n5282), .CK(CLK), .Q(n13976), .QN(n7969)
         );
  DFF_X1 \REGISTERS_reg[27][35]  ( .D(n5281), .CK(CLK), .Q(n13977), .QN(n7986)
         );
  DFF_X1 \REGISTERS_reg[27][34]  ( .D(n5280), .CK(CLK), .Q(n13978), .QN(n8003)
         );
  DFF_X1 \REGISTERS_reg[27][33]  ( .D(n5279), .CK(CLK), .Q(n13979), .QN(n8020)
         );
  DFF_X1 \REGISTERS_reg[27][32]  ( .D(n5278), .CK(CLK), .Q(n13980), .QN(n8037)
         );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n5277), .CK(CLK), .Q(n13981), .QN(n8054)
         );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n5276), .CK(CLK), .Q(n13982), .QN(n8071)
         );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n5275), .CK(CLK), .Q(n13983), .QN(n8088)
         );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n5274), .CK(CLK), .Q(n13984), .QN(n8105)
         );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n5273), .CK(CLK), .Q(n13985), .QN(n8122)
         );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n5272), .CK(CLK), .Q(n13986), .QN(n8139)
         );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n5271), .CK(CLK), .Q(n13987), .QN(n8156)
         );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n5270), .CK(CLK), .Q(n13988), .QN(n8173)
         );
  DFF_X1 \REGISTERS_reg[30][59]  ( .D(n5113), .CK(CLK), .Q(n13989), .QN(n7242)
         );
  DFF_X1 \REGISTERS_reg[30][58]  ( .D(n5112), .CK(CLK), .Q(n13990), .QN(n7259)
         );
  DFF_X1 \REGISTERS_reg[30][57]  ( .D(n5111), .CK(CLK), .Q(n13991), .QN(n7276)
         );
  DFF_X1 \REGISTERS_reg[30][56]  ( .D(n5110), .CK(CLK), .Q(n13992), .QN(n7375)
         );
  DFF_X1 \REGISTERS_reg[30][55]  ( .D(n5109), .CK(CLK), .Q(n13993), .QN(n7392)
         );
  DFF_X1 \REGISTERS_reg[30][54]  ( .D(n5108), .CK(CLK), .Q(n13994), .QN(n7494)
         );
  DFF_X1 \REGISTERS_reg[30][53]  ( .D(n5107), .CK(CLK), .Q(n13995), .QN(n7511)
         );
  DFF_X1 \REGISTERS_reg[30][52]  ( .D(n5106), .CK(CLK), .Q(n13996), .QN(n7528)
         );
  DFF_X1 \REGISTERS_reg[30][51]  ( .D(n5105), .CK(CLK), .Q(n13997), .QN(n7632)
         );
  DFF_X1 \REGISTERS_reg[30][50]  ( .D(n5104), .CK(CLK), .Q(n13998), .QN(n7649)
         );
  DFF_X1 \REGISTERS_reg[30][49]  ( .D(n5103), .CK(CLK), .Q(n13999), .QN(n7751)
         );
  DFF_X1 \REGISTERS_reg[30][48]  ( .D(n5102), .CK(CLK), .Q(n14000), .QN(n7768)
         );
  DFF_X1 \REGISTERS_reg[30][47]  ( .D(n5101), .CK(CLK), .Q(n14001), .QN(n7785)
         );
  DFF_X1 \REGISTERS_reg[30][46]  ( .D(n5100), .CK(CLK), .Q(n14002), .QN(n7802)
         );
  DFF_X1 \REGISTERS_reg[30][45]  ( .D(n5099), .CK(CLK), .Q(n14003), .QN(n7819)
         );
  DFF_X1 \REGISTERS_reg[30][44]  ( .D(n5098), .CK(CLK), .Q(n14004), .QN(n7836)
         );
  DFF_X1 \REGISTERS_reg[30][43]  ( .D(n5097), .CK(CLK), .Q(n14005), .QN(n7853)
         );
  DFF_X1 \REGISTERS_reg[30][42]  ( .D(n5096), .CK(CLK), .Q(n14006), .QN(n7870)
         );
  DFF_X1 \REGISTERS_reg[30][41]  ( .D(n5095), .CK(CLK), .Q(n14007), .QN(n7887)
         );
  DFF_X1 \REGISTERS_reg[30][40]  ( .D(n5094), .CK(CLK), .Q(n14008), .QN(n7904)
         );
  DFF_X1 \REGISTERS_reg[30][39]  ( .D(n5093), .CK(CLK), .Q(n14009), .QN(n7921)
         );
  DFF_X1 \REGISTERS_reg[30][38]  ( .D(n5092), .CK(CLK), .Q(n14010), .QN(n7938)
         );
  DFF_X1 \REGISTERS_reg[30][37]  ( .D(n5091), .CK(CLK), .Q(n14011), .QN(n7955)
         );
  DFF_X1 \REGISTERS_reg[30][36]  ( .D(n5090), .CK(CLK), .Q(n14012), .QN(n7972)
         );
  DFF_X1 \REGISTERS_reg[30][35]  ( .D(n5089), .CK(CLK), .Q(n14013), .QN(n7989)
         );
  DFF_X1 \REGISTERS_reg[30][34]  ( .D(n5088), .CK(CLK), .Q(n14014), .QN(n8006)
         );
  DFF_X1 \REGISTERS_reg[30][33]  ( .D(n5087), .CK(CLK), .Q(n14015), .QN(n8023)
         );
  DFF_X1 \REGISTERS_reg[30][32]  ( .D(n5086), .CK(CLK), .Q(n14016), .QN(n8040)
         );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n5085), .CK(CLK), .Q(n14017), .QN(n8057)
         );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n5084), .CK(CLK), .Q(n14018), .QN(n8074)
         );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n5083), .CK(CLK), .Q(n14019), .QN(n8091)
         );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n5082), .CK(CLK), .Q(n14020), .QN(n8108)
         );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n5081), .CK(CLK), .Q(n14021), .QN(n8125)
         );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n5080), .CK(CLK), .Q(n14022), .QN(n8142)
         );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n5079), .CK(CLK), .Q(n14023), .QN(n8159)
         );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n5078), .CK(CLK), .Q(n14024), .QN(n8176)
         );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n5333), .CK(CLK), .Q(n14060), .QN(n8191)
         );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n5332), .CK(CLK), .Q(n14061), .QN(n8208)
         );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n5331), .CK(CLK), .Q(n14062), .QN(n8225)
         );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n5330), .CK(CLK), .Q(n14063), .QN(n8242)
         );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n5329), .CK(CLK), .Q(n14064), .QN(n8259)
         );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n5328), .CK(CLK), .Q(n14065), .QN(n8276)
         );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n5327), .CK(CLK), .Q(n14066), .QN(n8293)
         );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n5326), .CK(CLK), .Q(n14067), .QN(n8310)
         );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n5325), .CK(CLK), .Q(n14068), .QN(n8327)
         );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n5324), .CK(CLK), .Q(n14069), .QN(n8344)
         );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n5323), .CK(CLK), .Q(n14070), .QN(n8361)
         );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n5322), .CK(CLK), .Q(n14071), .QN(n8378)
         );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n5321), .CK(CLK), .Q(n14072), .QN(n8395)
         );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n5320), .CK(CLK), .Q(n14073), .QN(n8412)
         );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n5319), .CK(CLK), .Q(n14074), .QN(n8429)
         );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n5318), .CK(CLK), .Q(n14075), .QN(n8446)
         );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n5317), .CK(CLK), .Q(n14076), .QN(n8463)
         );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n5316), .CK(CLK), .Q(n14077), .QN(n8480)
         );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n5315), .CK(CLK), .Q(n14078), .QN(n8497)
         );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n5313), .CK(CLK), .Q(n14079), .QN(n8531)
         );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n5314), .CK(CLK), .Q(n14080), .QN(n8514)
         );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n5312), .CK(CLK), .Q(n14081), .QN(n8548)
         );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n5311), .CK(CLK), .Q(n14082), .QN(n8565)
         );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n5310), .CK(CLK), .Q(n14153), .QN(n8582)
         );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n5269), .CK(CLK), .Q(n14107), .QN(n8190)
         );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n5268), .CK(CLK), .Q(n14108), .QN(n8207)
         );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n5267), .CK(CLK), .Q(n14109), .QN(n8224)
         );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n5266), .CK(CLK), .Q(n14110), .QN(n8241)
         );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n5265), .CK(CLK), .Q(n14111), .QN(n8258)
         );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n5264), .CK(CLK), .Q(n14112), .QN(n8275)
         );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n5263), .CK(CLK), .Q(n14113), .QN(n8292)
         );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n5262), .CK(CLK), .Q(n14114), .QN(n8309)
         );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n5261), .CK(CLK), .Q(n14115), .QN(n8326)
         );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n5260), .CK(CLK), .Q(n14116), .QN(n8343)
         );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n5259), .CK(CLK), .Q(n14117), .QN(n8360)
         );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n5258), .CK(CLK), .Q(n14118), .QN(n8377)
         );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n5257), .CK(CLK), .Q(n14119), .QN(n8394)
         );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n5256), .CK(CLK), .Q(n14120), .QN(n8411)
         );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n5255), .CK(CLK), .Q(n14121), .QN(n8428)
         );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n5254), .CK(CLK), .Q(n14122), .QN(n8445)
         );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n5253), .CK(CLK), .Q(n14123), .QN(n8462)
         );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n5252), .CK(CLK), .Q(n14124), .QN(n8479)
         );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n5251), .CK(CLK), .Q(n14125), .QN(n8496)
         );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n5249), .CK(CLK), .Q(n14126), .QN(n8530)
         );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n5250), .CK(CLK), .Q(n14127), .QN(n8513)
         );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n5248), .CK(CLK), .Q(n14128), .QN(n8547)
         );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n5247), .CK(CLK), .Q(n14129), .QN(n8564)
         );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n5246), .CK(CLK), .Q(n14154), .QN(n8581)
         );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n5077), .CK(CLK), .Q(n14130), .QN(n8193)
         );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n5076), .CK(CLK), .Q(n14131), .QN(n8210)
         );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n5075), .CK(CLK), .Q(n14132), .QN(n8227)
         );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n5074), .CK(CLK), .Q(n14133), .QN(n8244)
         );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n5073), .CK(CLK), .Q(n14134), .QN(n8261)
         );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n5072), .CK(CLK), .Q(n14135), .QN(n8278)
         );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n5071), .CK(CLK), .Q(n14136), .QN(n8295)
         );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n5070), .CK(CLK), .Q(n14137), .QN(n8312)
         );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n5069), .CK(CLK), .Q(n14138), .QN(n8329)
         );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n5068), .CK(CLK), .Q(n14139), .QN(n8346)
         );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n5067), .CK(CLK), .Q(n14140), .QN(n8363)
         );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n5066), .CK(CLK), .Q(n14141), .QN(n8380)
         );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n5065), .CK(CLK), .Q(n14142), .QN(n8397)
         );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n5064), .CK(CLK), .Q(n14143), .QN(n8414)
         );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n5063), .CK(CLK), .Q(n14144), .QN(n8431)
         );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n5062), .CK(CLK), .Q(n14145), .QN(n8448)
         );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n5061), .CK(CLK), .Q(n14146), .QN(n8465)
         );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n5060), .CK(CLK), .Q(n14147), .QN(n8482)
         );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n5059), .CK(CLK), .Q(n14148), .QN(n8499)
         );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n5057), .CK(CLK), .Q(n14149), .QN(n8533)
         );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n5058), .CK(CLK), .Q(n14150), .QN(n8516)
         );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n5056), .CK(CLK), .Q(n14151), .QN(n8550)
         );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n5055), .CK(CLK), .Q(n14152), .QN(n8567)
         );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n5054), .CK(CLK), .Q(n14155), .QN(n8584)
         );
  DFF_X1 \REGISTERS_reg[31][59]  ( .D(n5049), .CK(CLK), .Q(n14160), .QN(n7241)
         );
  DFF_X1 \REGISTERS_reg[31][58]  ( .D(n5048), .CK(CLK), .Q(n14161), .QN(n7258)
         );
  DFF_X1 \REGISTERS_reg[31][57]  ( .D(n5047), .CK(CLK), .Q(n14162), .QN(n7275)
         );
  DFF_X1 \REGISTERS_reg[31][56]  ( .D(n5046), .CK(CLK), .Q(n14163), .QN(n7374)
         );
  DFF_X1 \REGISTERS_reg[31][55]  ( .D(n5045), .CK(CLK), .Q(n14164), .QN(n7391)
         );
  DFF_X1 \REGISTERS_reg[31][54]  ( .D(n5044), .CK(CLK), .Q(n14165), .QN(n7493)
         );
  DFF_X1 \REGISTERS_reg[31][53]  ( .D(n5043), .CK(CLK), .Q(n14166), .QN(n7510)
         );
  DFF_X1 \REGISTERS_reg[31][52]  ( .D(n5042), .CK(CLK), .Q(n14167), .QN(n7527)
         );
  DFF_X1 \REGISTERS_reg[31][51]  ( .D(n5041), .CK(CLK), .Q(n14168), .QN(n7631)
         );
  DFF_X1 \REGISTERS_reg[31][50]  ( .D(n5040), .CK(CLK), .Q(n14169), .QN(n7648)
         );
  DFF_X1 \REGISTERS_reg[31][49]  ( .D(n5039), .CK(CLK), .Q(n14170), .QN(n7750)
         );
  DFF_X1 \REGISTERS_reg[31][48]  ( .D(n5038), .CK(CLK), .Q(n14171), .QN(n7767)
         );
  DFF_X1 \REGISTERS_reg[31][47]  ( .D(n5037), .CK(CLK), .Q(n14172), .QN(n7784)
         );
  DFF_X1 \REGISTERS_reg[31][46]  ( .D(n5036), .CK(CLK), .Q(n14173), .QN(n7801)
         );
  DFF_X1 \REGISTERS_reg[31][45]  ( .D(n5035), .CK(CLK), .Q(n14174), .QN(n7818)
         );
  DFF_X1 \REGISTERS_reg[31][44]  ( .D(n5034), .CK(CLK), .Q(n14175), .QN(n7835)
         );
  DFF_X1 \REGISTERS_reg[31][43]  ( .D(n5033), .CK(CLK), .Q(n14176), .QN(n7852)
         );
  DFF_X1 \REGISTERS_reg[31][42]  ( .D(n5032), .CK(CLK), .Q(n14177), .QN(n7869)
         );
  DFF_X1 \REGISTERS_reg[31][41]  ( .D(n5031), .CK(CLK), .Q(n14178), .QN(n7886)
         );
  DFF_X1 \REGISTERS_reg[31][40]  ( .D(n5030), .CK(CLK), .Q(n14179), .QN(n7903)
         );
  DFF_X1 \REGISTERS_reg[31][39]  ( .D(n5029), .CK(CLK), .Q(n14180), .QN(n7920)
         );
  DFF_X1 \REGISTERS_reg[31][38]  ( .D(n5028), .CK(CLK), .Q(n14181), .QN(n7937)
         );
  DFF_X1 \REGISTERS_reg[31][37]  ( .D(n5027), .CK(CLK), .Q(n14182), .QN(n7954)
         );
  DFF_X1 \REGISTERS_reg[31][36]  ( .D(n5026), .CK(CLK), .Q(n14183), .QN(n7971)
         );
  DFF_X1 \REGISTERS_reg[31][35]  ( .D(n5025), .CK(CLK), .Q(n14184), .QN(n7988)
         );
  DFF_X1 \REGISTERS_reg[31][34]  ( .D(n5024), .CK(CLK), .Q(n14185), .QN(n8005)
         );
  DFF_X1 \REGISTERS_reg[31][33]  ( .D(n5023), .CK(CLK), .Q(n14186), .QN(n8022)
         );
  DFF_X1 \REGISTERS_reg[31][32]  ( .D(n5022), .CK(CLK), .Q(n14187), .QN(n8039)
         );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n5021), .CK(CLK), .Q(n14188), .QN(n8056)
         );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n5020), .CK(CLK), .Q(n14189), .QN(n8073)
         );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n5019), .CK(CLK), .Q(n14190), .QN(n8090)
         );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n5018), .CK(CLK), .Q(n14191), .QN(n8107)
         );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n5017), .CK(CLK), .Q(n14192), .QN(n8124)
         );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n5016), .CK(CLK), .Q(n14193), .QN(n8141)
         );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n5015), .CK(CLK), .Q(n14194), .QN(n8158)
         );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n5014), .CK(CLK), .Q(n14195), .QN(n8175)
         );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n5013), .CK(CLK), .Q(n14196), .QN(n8192)
         );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n5012), .CK(CLK), .Q(n14197), .QN(n8209)
         );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n5011), .CK(CLK), .Q(n14198), .QN(n8226)
         );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n5010), .CK(CLK), .Q(n14199), .QN(n8243)
         );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n5009), .CK(CLK), .Q(n14200), .QN(n8260)
         );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n5008), .CK(CLK), .Q(n14201), .QN(n8277)
         );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n5007), .CK(CLK), .Q(n14202), .QN(n8294)
         );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n5006), .CK(CLK), .Q(n14203), .QN(n8311)
         );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n5005), .CK(CLK), .Q(n14204), .QN(n8328)
         );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n5004), .CK(CLK), .Q(n14205), .QN(n8345)
         );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n5003), .CK(CLK), .Q(n14206), .QN(n8362)
         );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n5002), .CK(CLK), .Q(n14207), .QN(n8379)
         );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n5001), .CK(CLK), .Q(n14208), .QN(n8396)
         );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n5000), .CK(CLK), .Q(n14209), .QN(n8413)
         );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n4999), .CK(CLK), .Q(n14210), .QN(n8430)
         );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n4998), .CK(CLK), .Q(n14211), .QN(n8447)
         );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n4997), .CK(CLK), .Q(n14212), .QN(n8464)
         );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n4996), .CK(CLK), .Q(n14213), .QN(n8481)
         );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n4995), .CK(CLK), .Q(n14214), .QN(n8498)
         );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n4994), .CK(CLK), .Q(n14215), .QN(n8515)
         );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n4993), .CK(CLK), .Q(n13828), .QN(n8532)
         );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n4992), .CK(CLK), .Q(n13829), .QN(n8549)
         );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n4991), .CK(CLK), .Q(n13830), .QN(n8566)
         );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n4990), .CK(CLK), .Q(n13831), .QN(n8583)
         );
  DFF_X1 \REGISTERS_reg[21][59]  ( .D(n5689), .CK(CLK), .QN(n7237) );
  DFF_X1 \REGISTERS_reg[21][58]  ( .D(n5688), .CK(CLK), .QN(n7254) );
  DFF_X1 \REGISTERS_reg[21][57]  ( .D(n5687), .CK(CLK), .QN(n7271) );
  DFF_X1 \REGISTERS_reg[21][56]  ( .D(n5686), .CK(CLK), .QN(n7370) );
  DFF_X1 \REGISTERS_reg[21][55]  ( .D(n5685), .CK(CLK), .QN(n7387) );
  DFF_X1 \REGISTERS_reg[21][54]  ( .D(n5684), .CK(CLK), .QN(n7404) );
  DFF_X1 \REGISTERS_reg[21][53]  ( .D(n5683), .CK(CLK), .QN(n7506) );
  DFF_X1 \REGISTERS_reg[21][52]  ( .D(n5682), .CK(CLK), .QN(n7523) );
  DFF_X1 \REGISTERS_reg[21][51]  ( .D(n5681), .CK(CLK), .QN(n7627) );
  DFF_X1 \REGISTERS_reg[21][50]  ( .D(n5680), .CK(CLK), .QN(n7644) );
  DFF_X1 \REGISTERS_reg[21][49]  ( .D(n5679), .CK(CLK), .QN(n7746) );
  DFF_X1 \REGISTERS_reg[21][48]  ( .D(n5678), .CK(CLK), .QN(n7763) );
  DFF_X1 \REGISTERS_reg[21][47]  ( .D(n5677), .CK(CLK), .QN(n7780) );
  DFF_X1 \REGISTERS_reg[21][46]  ( .D(n5676), .CK(CLK), .QN(n7797) );
  DFF_X1 \REGISTERS_reg[21][45]  ( .D(n5675), .CK(CLK), .QN(n7814) );
  DFF_X1 \REGISTERS_reg[21][44]  ( .D(n5674), .CK(CLK), .QN(n7831) );
  DFF_X1 \REGISTERS_reg[21][43]  ( .D(n5673), .CK(CLK), .QN(n7848) );
  DFF_X1 \REGISTERS_reg[21][42]  ( .D(n5672), .CK(CLK), .QN(n7865) );
  DFF_X1 \REGISTERS_reg[21][41]  ( .D(n5671), .CK(CLK), .QN(n7882) );
  DFF_X1 \REGISTERS_reg[21][40]  ( .D(n5670), .CK(CLK), .QN(n7899) );
  DFF_X1 \REGISTERS_reg[21][39]  ( .D(n5669), .CK(CLK), .QN(n7916) );
  DFF_X1 \REGISTERS_reg[21][38]  ( .D(n5668), .CK(CLK), .QN(n7933) );
  DFF_X1 \REGISTERS_reg[21][37]  ( .D(n5667), .CK(CLK), .QN(n7950) );
  DFF_X1 \REGISTERS_reg[21][36]  ( .D(n5666), .CK(CLK), .QN(n7967) );
  DFF_X1 \REGISTERS_reg[21][35]  ( .D(n5665), .CK(CLK), .QN(n7984) );
  NOR2_X1 U3 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n4450) );
  NOR2_X1 U4 ( .A1(n13389), .A2(ADD_RD2[1]), .ZN(n4454) );
  AND3_X1 U5 ( .A1(ENABLE), .A2(n12139), .A3(RD2), .ZN(n3211) );
  NAND2_X1 U6 ( .A1(n3209), .A2(n3189), .ZN(n1995) );
  CLKBUF_X1 U7 ( .A(n12614), .Z(n12612) );
  CLKBUF_X1 U8 ( .A(n12690), .Z(n12688) );
  CLKBUF_X1 U9 ( .A(n12633), .Z(n12631) );
  CLKBUF_X1 U10 ( .A(n12709), .Z(n12707) );
  CLKBUF_X1 U11 ( .A(n12595), .Z(n12593) );
  CLKBUF_X1 U12 ( .A(n12652), .Z(n12650) );
  CLKBUF_X1 U13 ( .A(n12671), .Z(n12669) );
  BUF_X1 U14 ( .A(n1910), .Z(n13130) );
  BUF_X1 U15 ( .A(n1912), .Z(n13110) );
  BUF_X1 U16 ( .A(n1914), .Z(n13090) );
  BUF_X1 U17 ( .A(n1916), .Z(n13070) );
  BUF_X1 U18 ( .A(n1918), .Z(n13050) );
  BUF_X1 U19 ( .A(n1920), .Z(n13030) );
  BUF_X1 U20 ( .A(n1908), .Z(n13150) );
  BUF_X1 U21 ( .A(n1842), .Z(n13359) );
  BUF_X1 U22 ( .A(n1932), .Z(n12850) );
  BUF_X1 U23 ( .A(n1934), .Z(n12830) );
  BUF_X1 U24 ( .A(n1937), .Z(n12770) );
  BUF_X1 U25 ( .A(n1938), .Z(n12750) );
  BUF_X1 U26 ( .A(n1940), .Z(n12710) );
  BUF_X1 U27 ( .A(n1939), .Z(n12730) );
  BUF_X1 U28 ( .A(n1936), .Z(n12790) );
  BUF_X1 U29 ( .A(n1935), .Z(n12810) );
  BUF_X1 U30 ( .A(n1928), .Z(n12930) );
  BUF_X1 U31 ( .A(n1923), .Z(n13010) );
  BUF_X1 U32 ( .A(n1925), .Z(n12990) );
  BUF_X1 U33 ( .A(n1929), .Z(n12910) );
  BUF_X1 U34 ( .A(n1948), .Z(n12577) );
  BUF_X1 U35 ( .A(n1945), .Z(n12634) );
  BUF_X1 U36 ( .A(n1947), .Z(n12596) );
  BUF_X1 U37 ( .A(n1931), .Z(n12870) );
  BUF_X1 U38 ( .A(n1930), .Z(n12890) );
  BUF_X1 U39 ( .A(n1927), .Z(n12950) );
  BUF_X1 U40 ( .A(n1944), .Z(n12653) );
  BUF_X1 U41 ( .A(n1946), .Z(n12615) );
  BUF_X1 U42 ( .A(n1943), .Z(n12672) );
  BUF_X1 U43 ( .A(n1941), .Z(n12691) );
  BUF_X1 U44 ( .A(n1926), .Z(n12970) );
  INV_X1 U45 ( .A(n12573), .ZN(n12552) );
  INV_X1 U46 ( .A(n12573), .ZN(n12553) );
  INV_X1 U47 ( .A(n12573), .ZN(n12554) );
  INV_X1 U48 ( .A(n12573), .ZN(n12555) );
  INV_X1 U49 ( .A(n12573), .ZN(n12551) );
  INV_X1 U50 ( .A(n13128), .ZN(n13112) );
  INV_X1 U51 ( .A(n13128), .ZN(n13113) );
  INV_X1 U52 ( .A(n13128), .ZN(n13114) );
  INV_X1 U53 ( .A(n13007), .ZN(n12991) );
  INV_X1 U54 ( .A(n12847), .ZN(n12831) );
  INV_X1 U55 ( .A(n12787), .ZN(n12771) );
  INV_X1 U56 ( .A(n12767), .ZN(n12751) );
  INV_X1 U57 ( .A(n12927), .ZN(n12911) );
  INV_X1 U58 ( .A(n13027), .ZN(n13011) );
  INV_X1 U59 ( .A(n13067), .ZN(n13051) );
  INV_X1 U60 ( .A(n13047), .ZN(n13031) );
  INV_X1 U61 ( .A(n12928), .ZN(n12912) );
  INV_X1 U62 ( .A(n12928), .ZN(n12913) );
  INV_X1 U63 ( .A(n12928), .ZN(n12914) );
  INV_X1 U64 ( .A(n12948), .ZN(n12932) );
  INV_X1 U65 ( .A(n12948), .ZN(n12933) );
  INV_X1 U66 ( .A(n12948), .ZN(n12934) );
  INV_X1 U67 ( .A(n13028), .ZN(n13012) );
  INV_X1 U68 ( .A(n13028), .ZN(n13013) );
  INV_X1 U69 ( .A(n13028), .ZN(n13014) );
  INV_X1 U70 ( .A(n13008), .ZN(n12992) );
  INV_X1 U71 ( .A(n13008), .ZN(n12993) );
  INV_X1 U72 ( .A(n13008), .ZN(n12994) );
  INV_X1 U73 ( .A(n13068), .ZN(n13052) );
  INV_X1 U74 ( .A(n13068), .ZN(n13053) );
  INV_X1 U75 ( .A(n13068), .ZN(n13054) );
  INV_X1 U76 ( .A(n13048), .ZN(n13032) );
  INV_X1 U77 ( .A(n13048), .ZN(n13033) );
  INV_X1 U78 ( .A(n13048), .ZN(n13034) );
  INV_X1 U79 ( .A(n12867), .ZN(n12851) );
  INV_X1 U80 ( .A(n12868), .ZN(n12852) );
  INV_X1 U81 ( .A(n12868), .ZN(n12853) );
  INV_X1 U82 ( .A(n12868), .ZN(n12854) );
  INV_X1 U83 ( .A(n12848), .ZN(n12832) );
  INV_X1 U84 ( .A(n12848), .ZN(n12833) );
  INV_X1 U85 ( .A(n12848), .ZN(n12834) );
  INV_X1 U86 ( .A(n12788), .ZN(n12772) );
  INV_X1 U87 ( .A(n12788), .ZN(n12773) );
  INV_X1 U88 ( .A(n12788), .ZN(n12774) );
  INV_X1 U89 ( .A(n12768), .ZN(n12752) );
  INV_X1 U90 ( .A(n12768), .ZN(n12753) );
  INV_X1 U91 ( .A(n12768), .ZN(n12754) );
  INV_X1 U92 ( .A(n12594), .ZN(n12578) );
  INV_X1 U93 ( .A(n12594), .ZN(n12579) );
  INV_X1 U94 ( .A(n12594), .ZN(n12580) );
  INV_X1 U95 ( .A(n12651), .ZN(n12635) );
  INV_X1 U96 ( .A(n12651), .ZN(n12636) );
  INV_X1 U97 ( .A(n12651), .ZN(n12637) );
  INV_X1 U98 ( .A(n12670), .ZN(n12654) );
  INV_X1 U99 ( .A(n12670), .ZN(n12655) );
  INV_X1 U100 ( .A(n12670), .ZN(n12656) );
  INV_X1 U101 ( .A(n13127), .ZN(n13111) );
  INV_X1 U102 ( .A(n13147), .ZN(n13131) );
  INV_X1 U103 ( .A(n13107), .ZN(n13091) );
  INV_X1 U104 ( .A(n13087), .ZN(n13071) );
  INV_X1 U105 ( .A(n13376), .ZN(n13360) );
  INV_X1 U106 ( .A(n12807), .ZN(n12791) );
  INV_X1 U107 ( .A(n12727), .ZN(n12711) );
  INV_X1 U108 ( .A(n12747), .ZN(n12731) );
  INV_X1 U109 ( .A(n12827), .ZN(n12811) );
  INV_X1 U110 ( .A(n12887), .ZN(n12871) );
  INV_X1 U111 ( .A(n12907), .ZN(n12891) );
  INV_X1 U112 ( .A(n12967), .ZN(n12951) );
  INV_X1 U113 ( .A(n12987), .ZN(n12971) );
  INV_X1 U114 ( .A(n13167), .ZN(n13151) );
  INV_X1 U115 ( .A(n13168), .ZN(n13154) );
  INV_X1 U116 ( .A(n13168), .ZN(n13153) );
  INV_X1 U117 ( .A(n13377), .ZN(n13361) );
  INV_X1 U118 ( .A(n13148), .ZN(n13132) );
  INV_X1 U119 ( .A(n13148), .ZN(n13133) );
  INV_X1 U120 ( .A(n13148), .ZN(n13134) );
  INV_X1 U121 ( .A(n13108), .ZN(n13092) );
  INV_X1 U122 ( .A(n13108), .ZN(n13093) );
  INV_X1 U123 ( .A(n13108), .ZN(n13094) );
  INV_X1 U124 ( .A(n13088), .ZN(n13072) );
  INV_X1 U125 ( .A(n13088), .ZN(n13073) );
  INV_X1 U126 ( .A(n13088), .ZN(n13074) );
  INV_X1 U127 ( .A(n12808), .ZN(n12792) );
  INV_X1 U128 ( .A(n12728), .ZN(n12713) );
  INV_X1 U129 ( .A(n12728), .ZN(n12712) );
  INV_X1 U130 ( .A(n12613), .ZN(n12599) );
  INV_X1 U131 ( .A(n12689), .ZN(n12674) );
  INV_X1 U132 ( .A(n12613), .ZN(n12597) );
  INV_X1 U133 ( .A(n12613), .ZN(n12598) );
  INV_X1 U134 ( .A(n12689), .ZN(n12673) );
  INV_X1 U135 ( .A(n12632), .ZN(n12616) );
  INV_X1 U136 ( .A(n12632), .ZN(n12617) );
  INV_X1 U137 ( .A(n12632), .ZN(n12618) );
  INV_X1 U138 ( .A(n12689), .ZN(n12675) );
  INV_X1 U139 ( .A(n12708), .ZN(n12692) );
  INV_X1 U140 ( .A(n12708), .ZN(n12693) );
  INV_X1 U141 ( .A(n12708), .ZN(n12694) );
  INV_X1 U142 ( .A(n12728), .ZN(n12714) );
  INV_X1 U143 ( .A(n12748), .ZN(n12732) );
  INV_X1 U144 ( .A(n12748), .ZN(n12733) );
  INV_X1 U145 ( .A(n12748), .ZN(n12734) );
  INV_X1 U146 ( .A(n12808), .ZN(n12793) );
  INV_X1 U147 ( .A(n12808), .ZN(n12794) );
  INV_X1 U148 ( .A(n12828), .ZN(n12812) );
  INV_X1 U149 ( .A(n12828), .ZN(n12813) );
  INV_X1 U150 ( .A(n12828), .ZN(n12814) );
  INV_X1 U151 ( .A(n12888), .ZN(n12872) );
  INV_X1 U152 ( .A(n12888), .ZN(n12873) );
  INV_X1 U153 ( .A(n12888), .ZN(n12874) );
  INV_X1 U154 ( .A(n12908), .ZN(n12892) );
  INV_X1 U155 ( .A(n12908), .ZN(n12893) );
  INV_X1 U156 ( .A(n12908), .ZN(n12894) );
  INV_X1 U157 ( .A(n12968), .ZN(n12952) );
  INV_X1 U158 ( .A(n12968), .ZN(n12953) );
  INV_X1 U159 ( .A(n12968), .ZN(n12954) );
  INV_X1 U160 ( .A(n12988), .ZN(n12972) );
  INV_X1 U161 ( .A(n12988), .ZN(n12973) );
  INV_X1 U162 ( .A(n12988), .ZN(n12974) );
  INV_X1 U163 ( .A(n13168), .ZN(n13152) );
  INV_X1 U164 ( .A(n13377), .ZN(n13362) );
  INV_X1 U165 ( .A(n13377), .ZN(n13363) );
  INV_X1 U166 ( .A(n12947), .ZN(n12931) );
  BUF_X1 U167 ( .A(n12575), .Z(n12573) );
  BUF_X1 U168 ( .A(n12576), .Z(n12571) );
  BUF_X1 U169 ( .A(n12574), .Z(n12570) );
  BUF_X1 U170 ( .A(n12575), .Z(n12569) );
  BUF_X1 U171 ( .A(n12574), .Z(n12568) );
  BUF_X1 U172 ( .A(n12574), .Z(n12567) );
  BUF_X1 U173 ( .A(n12574), .Z(n12566) );
  BUF_X1 U174 ( .A(n12574), .Z(n12565) );
  BUF_X1 U175 ( .A(n12575), .Z(n12564) );
  BUF_X1 U176 ( .A(n12575), .Z(n12563) );
  BUF_X1 U177 ( .A(n12575), .Z(n12562) );
  BUF_X1 U178 ( .A(n12576), .Z(n12561) );
  BUF_X1 U179 ( .A(n12576), .Z(n12560) );
  BUF_X1 U180 ( .A(n12576), .Z(n12559) );
  BUF_X1 U181 ( .A(n12574), .Z(n12572) );
  BUF_X1 U182 ( .A(n12576), .Z(n12558) );
  BUF_X1 U183 ( .A(n12576), .Z(n12557) );
  BUF_X1 U184 ( .A(n1998), .Z(n12357) );
  BUF_X1 U185 ( .A(n1998), .Z(n12358) );
  BUF_X1 U186 ( .A(n1998), .Z(n12359) );
  BUF_X1 U187 ( .A(n1998), .Z(n12360) );
  BUF_X1 U188 ( .A(n1998), .Z(n12361) );
  BUF_X1 U189 ( .A(n12929), .Z(n12927) );
  BUF_X1 U190 ( .A(n12949), .Z(n12947) );
  BUF_X1 U191 ( .A(n13009), .Z(n13007) );
  BUF_X1 U192 ( .A(n13149), .Z(n13147) );
  BUF_X1 U193 ( .A(n13109), .Z(n13107) );
  BUF_X1 U194 ( .A(n13089), .Z(n13087) );
  BUF_X1 U195 ( .A(n13378), .Z(n13376) );
  BUF_X1 U196 ( .A(n12849), .Z(n12847) );
  BUF_X1 U197 ( .A(n12789), .Z(n12787) );
  BUF_X1 U198 ( .A(n12769), .Z(n12767) );
  BUF_X1 U199 ( .A(n12729), .Z(n12727) );
  BUF_X1 U200 ( .A(n12749), .Z(n12747) );
  BUF_X1 U201 ( .A(n12809), .Z(n12807) );
  BUF_X1 U202 ( .A(n12829), .Z(n12827) );
  BUF_X1 U203 ( .A(n12889), .Z(n12887) );
  BUF_X1 U204 ( .A(n12909), .Z(n12907) );
  BUF_X1 U205 ( .A(n12969), .Z(n12967) );
  BUF_X1 U206 ( .A(n12989), .Z(n12987) );
  BUF_X1 U207 ( .A(n13169), .Z(n13167) );
  BUF_X1 U208 ( .A(n13021), .Z(n13024) );
  BUF_X1 U209 ( .A(n13020), .Z(n13023) );
  BUF_X1 U210 ( .A(n13041), .Z(n13044) );
  BUF_X1 U211 ( .A(n13040), .Z(n13043) );
  BUF_X1 U212 ( .A(n13015), .Z(n13022) );
  BUF_X1 U213 ( .A(n13029), .Z(n13021) );
  BUF_X1 U214 ( .A(n13029), .Z(n13020) );
  BUF_X1 U215 ( .A(n13029), .Z(n13019) );
  BUF_X1 U216 ( .A(n13029), .Z(n13018) );
  BUF_X1 U217 ( .A(n13029), .Z(n13017) );
  BUF_X1 U218 ( .A(n13029), .Z(n13016) );
  BUF_X1 U219 ( .A(n13035), .Z(n13042) );
  BUF_X1 U220 ( .A(n13049), .Z(n13041) );
  BUF_X1 U221 ( .A(n13049), .Z(n13040) );
  BUF_X1 U222 ( .A(n13049), .Z(n13039) );
  BUF_X1 U223 ( .A(n13049), .Z(n13038) );
  BUF_X1 U224 ( .A(n13049), .Z(n13037) );
  BUF_X1 U225 ( .A(n13049), .Z(n13036) );
  BUF_X1 U226 ( .A(n13029), .Z(n13015) );
  BUF_X1 U227 ( .A(n13049), .Z(n13035) );
  BUF_X1 U228 ( .A(n12929), .Z(n12926) );
  BUF_X1 U229 ( .A(n12929), .Z(n12925) );
  BUF_X1 U230 ( .A(n12929), .Z(n12924) );
  BUF_X1 U231 ( .A(n12929), .Z(n12923) );
  BUF_X1 U232 ( .A(n12941), .Z(n12944) );
  BUF_X1 U233 ( .A(n13009), .Z(n13006) );
  BUF_X1 U234 ( .A(n13009), .Z(n13005) );
  BUF_X1 U235 ( .A(n13009), .Z(n13004) );
  BUF_X1 U236 ( .A(n13009), .Z(n13003) );
  BUF_X1 U237 ( .A(n13371), .Z(n13369) );
  BUF_X1 U238 ( .A(n13375), .Z(n13368) );
  BUF_X1 U239 ( .A(n13162), .Z(n13158) );
  BUF_X1 U240 ( .A(n13166), .Z(n13157) );
  BUF_X1 U241 ( .A(n13165), .Z(n13156) );
  BUF_X1 U242 ( .A(n13164), .Z(n13155) );
  BUF_X1 U243 ( .A(n13149), .Z(n13146) );
  BUF_X1 U244 ( .A(n13149), .Z(n13145) );
  BUF_X1 U245 ( .A(n13149), .Z(n13144) );
  BUF_X1 U246 ( .A(n13149), .Z(n13143) );
  BUF_X1 U247 ( .A(n13121), .Z(n13124) );
  BUF_X1 U248 ( .A(n13120), .Z(n13123) );
  BUF_X1 U249 ( .A(n13109), .Z(n13106) );
  BUF_X1 U250 ( .A(n13109), .Z(n13105) );
  BUF_X1 U251 ( .A(n13109), .Z(n13104) );
  BUF_X1 U252 ( .A(n13109), .Z(n13103) );
  BUF_X1 U253 ( .A(n13089), .Z(n13086) );
  BUF_X1 U254 ( .A(n13089), .Z(n13085) );
  BUF_X1 U255 ( .A(n13089), .Z(n13084) );
  BUF_X1 U256 ( .A(n13089), .Z(n13083) );
  BUF_X1 U257 ( .A(n13061), .Z(n13064) );
  BUF_X1 U258 ( .A(n13060), .Z(n13063) );
  BUF_X1 U259 ( .A(n12889), .Z(n12886) );
  BUF_X1 U260 ( .A(n12889), .Z(n12885) );
  BUF_X1 U261 ( .A(n12969), .Z(n12966) );
  BUF_X1 U262 ( .A(n12969), .Z(n12965) );
  BUF_X1 U263 ( .A(n12929), .Z(n12922) );
  BUF_X1 U264 ( .A(n12922), .Z(n12921) );
  BUF_X1 U265 ( .A(n12926), .Z(n12920) );
  BUF_X1 U266 ( .A(n12925), .Z(n12919) );
  BUF_X1 U267 ( .A(n12924), .Z(n12918) );
  BUF_X1 U268 ( .A(n12923), .Z(n12917) );
  BUF_X1 U269 ( .A(n12922), .Z(n12916) );
  BUF_X1 U270 ( .A(n12940), .Z(n12942) );
  BUF_X1 U271 ( .A(n12949), .Z(n12941) );
  BUF_X1 U272 ( .A(n12949), .Z(n12940) );
  BUF_X1 U273 ( .A(n12949), .Z(n12939) );
  BUF_X1 U274 ( .A(n12949), .Z(n12938) );
  BUF_X1 U275 ( .A(n12949), .Z(n12937) );
  BUF_X1 U276 ( .A(n12949), .Z(n12936) );
  BUF_X1 U277 ( .A(n13009), .Z(n13002) );
  BUF_X1 U278 ( .A(n13002), .Z(n13001) );
  BUF_X1 U279 ( .A(n13006), .Z(n13000) );
  BUF_X1 U280 ( .A(n13005), .Z(n12999) );
  BUF_X1 U281 ( .A(n13004), .Z(n12998) );
  BUF_X1 U282 ( .A(n13003), .Z(n12997) );
  BUF_X1 U283 ( .A(n13002), .Z(n12996) );
  BUF_X1 U284 ( .A(n13163), .Z(n13161) );
  BUF_X1 U285 ( .A(n13162), .Z(n13160) );
  BUF_X1 U286 ( .A(n13166), .Z(n13159) );
  BUF_X1 U287 ( .A(n13378), .Z(n13375) );
  BUF_X1 U288 ( .A(n13378), .Z(n13374) );
  BUF_X1 U289 ( .A(n13378), .Z(n13373) );
  BUF_X1 U290 ( .A(n13378), .Z(n13372) );
  BUF_X1 U291 ( .A(n13378), .Z(n13371) );
  BUF_X1 U292 ( .A(n13374), .Z(n13370) );
  BUF_X1 U293 ( .A(n13149), .Z(n13142) );
  BUF_X1 U294 ( .A(n13142), .Z(n13141) );
  BUF_X1 U295 ( .A(n13146), .Z(n13140) );
  BUF_X1 U296 ( .A(n13145), .Z(n13139) );
  BUF_X1 U297 ( .A(n13144), .Z(n13138) );
  BUF_X1 U298 ( .A(n13143), .Z(n13137) );
  BUF_X1 U299 ( .A(n13142), .Z(n13136) );
  BUF_X1 U300 ( .A(n13119), .Z(n13122) );
  BUF_X1 U301 ( .A(n13129), .Z(n13121) );
  BUF_X1 U302 ( .A(n13129), .Z(n13120) );
  BUF_X1 U303 ( .A(n13129), .Z(n13119) );
  BUF_X1 U304 ( .A(n13129), .Z(n13118) );
  BUF_X1 U305 ( .A(n13129), .Z(n13117) );
  BUF_X1 U306 ( .A(n13129), .Z(n13116) );
  BUF_X1 U307 ( .A(n13109), .Z(n13102) );
  BUF_X1 U308 ( .A(n13102), .Z(n13101) );
  BUF_X1 U309 ( .A(n13106), .Z(n13100) );
  BUF_X1 U310 ( .A(n13105), .Z(n13099) );
  BUF_X1 U311 ( .A(n13104), .Z(n13098) );
  BUF_X1 U312 ( .A(n13103), .Z(n13097) );
  BUF_X1 U313 ( .A(n13102), .Z(n13096) );
  BUF_X1 U314 ( .A(n13089), .Z(n13082) );
  BUF_X1 U315 ( .A(n13082), .Z(n13081) );
  BUF_X1 U316 ( .A(n13086), .Z(n13080) );
  BUF_X1 U317 ( .A(n13085), .Z(n13079) );
  BUF_X1 U318 ( .A(n13084), .Z(n13078) );
  BUF_X1 U319 ( .A(n13083), .Z(n13077) );
  BUF_X1 U320 ( .A(n13082), .Z(n13076) );
  BUF_X1 U321 ( .A(n13055), .Z(n13062) );
  BUF_X1 U322 ( .A(n13069), .Z(n13061) );
  BUF_X1 U323 ( .A(n13069), .Z(n13060) );
  BUF_X1 U324 ( .A(n13069), .Z(n13059) );
  BUF_X1 U325 ( .A(n13069), .Z(n13058) );
  BUF_X1 U326 ( .A(n13069), .Z(n13057) );
  BUF_X1 U327 ( .A(n13069), .Z(n13056) );
  BUF_X1 U328 ( .A(n12861), .Z(n12864) );
  BUF_X1 U329 ( .A(n12860), .Z(n12863) );
  BUF_X1 U330 ( .A(n12849), .Z(n12846) );
  BUF_X1 U331 ( .A(n12849), .Z(n12845) );
  BUF_X1 U332 ( .A(n12849), .Z(n12844) );
  BUF_X1 U333 ( .A(n12849), .Z(n12843) );
  BUF_X1 U334 ( .A(n12809), .Z(n12802) );
  BUF_X1 U335 ( .A(n12802), .Z(n12801) );
  BUF_X1 U336 ( .A(n12806), .Z(n12800) );
  BUF_X1 U337 ( .A(n12805), .Z(n12799) );
  BUF_X1 U338 ( .A(n12789), .Z(n12786) );
  BUF_X1 U339 ( .A(n12789), .Z(n12785) );
  BUF_X1 U340 ( .A(n12789), .Z(n12784) );
  BUF_X1 U341 ( .A(n12789), .Z(n12783) );
  BUF_X1 U342 ( .A(n12769), .Z(n12766) );
  BUF_X1 U343 ( .A(n12769), .Z(n12765) );
  BUF_X1 U344 ( .A(n12769), .Z(n12764) );
  BUF_X1 U345 ( .A(n12769), .Z(n12763) );
  BUF_X1 U346 ( .A(n12722), .Z(n12721) );
  BUF_X1 U347 ( .A(n12726), .Z(n12720) );
  BUF_X1 U348 ( .A(n12725), .Z(n12719) );
  BUF_X1 U349 ( .A(n12724), .Z(n12718) );
  BUF_X1 U350 ( .A(n12729), .Z(n12726) );
  BUF_X1 U351 ( .A(n12729), .Z(n12725) );
  BUF_X1 U352 ( .A(n12855), .Z(n12862) );
  BUF_X1 U353 ( .A(n12869), .Z(n12861) );
  BUF_X1 U354 ( .A(n12869), .Z(n12860) );
  BUF_X1 U355 ( .A(n12869), .Z(n12859) );
  BUF_X1 U356 ( .A(n12869), .Z(n12858) );
  BUF_X1 U357 ( .A(n12869), .Z(n12857) );
  BUF_X1 U358 ( .A(n12869), .Z(n12856) );
  BUF_X1 U359 ( .A(n12849), .Z(n12842) );
  BUF_X1 U360 ( .A(n12842), .Z(n12841) );
  BUF_X1 U361 ( .A(n12846), .Z(n12840) );
  BUF_X1 U362 ( .A(n12845), .Z(n12839) );
  BUF_X1 U363 ( .A(n12844), .Z(n12838) );
  BUF_X1 U364 ( .A(n12843), .Z(n12837) );
  BUF_X1 U365 ( .A(n12845), .Z(n12836) );
  BUF_X1 U366 ( .A(n12809), .Z(n12806) );
  BUF_X1 U367 ( .A(n12809), .Z(n12805) );
  BUF_X1 U368 ( .A(n12809), .Z(n12804) );
  BUF_X1 U369 ( .A(n12809), .Z(n12803) );
  BUF_X1 U370 ( .A(n12789), .Z(n12782) );
  BUF_X1 U371 ( .A(n12782), .Z(n12781) );
  BUF_X1 U372 ( .A(n12786), .Z(n12780) );
  BUF_X1 U373 ( .A(n12785), .Z(n12779) );
  BUF_X1 U374 ( .A(n12784), .Z(n12778) );
  BUF_X1 U375 ( .A(n12783), .Z(n12777) );
  BUF_X1 U376 ( .A(n12785), .Z(n12776) );
  BUF_X1 U377 ( .A(n12769), .Z(n12762) );
  BUF_X1 U378 ( .A(n12762), .Z(n12761) );
  BUF_X1 U379 ( .A(n12766), .Z(n12760) );
  BUF_X1 U380 ( .A(n12765), .Z(n12759) );
  BUF_X1 U381 ( .A(n12764), .Z(n12758) );
  BUF_X1 U382 ( .A(n12763), .Z(n12757) );
  BUF_X1 U383 ( .A(n12765), .Z(n12756) );
  BUF_X1 U384 ( .A(n12729), .Z(n12724) );
  BUF_X1 U385 ( .A(n12729), .Z(n12723) );
  BUF_X1 U386 ( .A(n12729), .Z(n12722) );
  BUF_X1 U387 ( .A(n12595), .Z(n12592) );
  BUF_X1 U388 ( .A(n12595), .Z(n12591) );
  BUF_X1 U389 ( .A(n12595), .Z(n12590) );
  BUF_X1 U390 ( .A(n12595), .Z(n12589) );
  BUF_X1 U391 ( .A(n12652), .Z(n12649) );
  BUF_X1 U392 ( .A(n12652), .Z(n12648) );
  BUF_X1 U393 ( .A(n12652), .Z(n12647) );
  BUF_X1 U394 ( .A(n12652), .Z(n12646) );
  BUF_X1 U395 ( .A(n12611), .Z(n12603) );
  BUF_X1 U396 ( .A(n12610), .Z(n12602) );
  BUF_X1 U397 ( .A(n12609), .Z(n12601) );
  BUF_X1 U398 ( .A(n12608), .Z(n12600) );
  BUF_X1 U399 ( .A(n12671), .Z(n12668) );
  BUF_X1 U400 ( .A(n12671), .Z(n12667) );
  BUF_X1 U401 ( .A(n12671), .Z(n12666) );
  BUF_X1 U402 ( .A(n12671), .Z(n12665) );
  BUF_X1 U403 ( .A(n12687), .Z(n12682) );
  BUF_X1 U404 ( .A(n12686), .Z(n12681) );
  BUF_X1 U405 ( .A(n12685), .Z(n12680) );
  BUF_X1 U406 ( .A(n12684), .Z(n12679) );
  BUF_X1 U407 ( .A(n12614), .Z(n12610) );
  BUF_X1 U408 ( .A(n12595), .Z(n12588) );
  BUF_X1 U409 ( .A(n12588), .Z(n12587) );
  BUF_X1 U410 ( .A(n12592), .Z(n12586) );
  BUF_X1 U411 ( .A(n12590), .Z(n12585) );
  BUF_X1 U412 ( .A(n12589), .Z(n12584) );
  BUF_X1 U413 ( .A(n12590), .Z(n12583) );
  BUF_X1 U414 ( .A(n12589), .Z(n12582) );
  BUF_X1 U415 ( .A(n12652), .Z(n12645) );
  BUF_X1 U416 ( .A(n12645), .Z(n12644) );
  BUF_X1 U417 ( .A(n12649), .Z(n12643) );
  BUF_X1 U418 ( .A(n12647), .Z(n12642) );
  BUF_X1 U419 ( .A(n12646), .Z(n12641) );
  BUF_X1 U420 ( .A(n12647), .Z(n12640) );
  BUF_X1 U421 ( .A(n12646), .Z(n12639) );
  BUF_X1 U422 ( .A(n12614), .Z(n12609) );
  BUF_X1 U423 ( .A(n12614), .Z(n12608) );
  BUF_X1 U424 ( .A(n12614), .Z(n12607) );
  BUF_X1 U425 ( .A(n12607), .Z(n12606) );
  BUF_X1 U426 ( .A(n12607), .Z(n12605) );
  BUF_X1 U427 ( .A(n12611), .Z(n12604) );
  BUF_X1 U428 ( .A(n12671), .Z(n12664) );
  BUF_X1 U429 ( .A(n12664), .Z(n12663) );
  BUF_X1 U430 ( .A(n12668), .Z(n12662) );
  BUF_X1 U431 ( .A(n12666), .Z(n12661) );
  BUF_X1 U432 ( .A(n12665), .Z(n12660) );
  BUF_X1 U433 ( .A(n12666), .Z(n12659) );
  BUF_X1 U434 ( .A(n12665), .Z(n12658) );
  BUF_X1 U435 ( .A(n12690), .Z(n12687) );
  BUF_X1 U436 ( .A(n12690), .Z(n12686) );
  BUF_X1 U437 ( .A(n12690), .Z(n12685) );
  BUF_X1 U438 ( .A(n12690), .Z(n12684) );
  BUF_X1 U439 ( .A(n12690), .Z(n12683) );
  BUF_X1 U440 ( .A(n12926), .Z(n12915) );
  BUF_X1 U441 ( .A(n12949), .Z(n12935) );
  BUF_X1 U442 ( .A(n13006), .Z(n12995) );
  BUF_X1 U443 ( .A(n13146), .Z(n13135) );
  BUF_X1 U444 ( .A(n13129), .Z(n13115) );
  BUF_X1 U445 ( .A(n13106), .Z(n13095) );
  BUF_X1 U446 ( .A(n13086), .Z(n13075) );
  BUF_X1 U447 ( .A(n13069), .Z(n13055) );
  BUF_X1 U448 ( .A(n12869), .Z(n12855) );
  BUF_X1 U449 ( .A(n12842), .Z(n12835) );
  BUF_X1 U450 ( .A(n12782), .Z(n12775) );
  BUF_X1 U451 ( .A(n12762), .Z(n12755) );
  BUF_X1 U452 ( .A(n12591), .Z(n12581) );
  BUF_X1 U453 ( .A(n12648), .Z(n12638) );
  BUF_X1 U454 ( .A(n12667), .Z(n12657) );
  BUF_X1 U455 ( .A(n12614), .Z(n12611) );
  BUF_X1 U456 ( .A(n12633), .Z(n12630) );
  BUF_X1 U457 ( .A(n12633), .Z(n12629) );
  BUF_X1 U458 ( .A(n12633), .Z(n12628) );
  BUF_X1 U459 ( .A(n12633), .Z(n12627) );
  BUF_X1 U460 ( .A(n12633), .Z(n12626) );
  BUF_X1 U461 ( .A(n12630), .Z(n12625) );
  BUF_X1 U462 ( .A(n12629), .Z(n12624) );
  BUF_X1 U463 ( .A(n12628), .Z(n12623) );
  BUF_X1 U464 ( .A(n12627), .Z(n12622) );
  BUF_X1 U465 ( .A(n12626), .Z(n12621) );
  BUF_X1 U466 ( .A(n12628), .Z(n12620) );
  BUF_X1 U467 ( .A(n12630), .Z(n12619) );
  BUF_X1 U468 ( .A(n12683), .Z(n12678) );
  BUF_X1 U469 ( .A(n12687), .Z(n12677) );
  BUF_X1 U470 ( .A(n12686), .Z(n12676) );
  BUF_X1 U471 ( .A(n12709), .Z(n12706) );
  BUF_X1 U472 ( .A(n12709), .Z(n12705) );
  BUF_X1 U473 ( .A(n12709), .Z(n12704) );
  BUF_X1 U474 ( .A(n12709), .Z(n12703) );
  BUF_X1 U475 ( .A(n12709), .Z(n12702) );
  BUF_X1 U476 ( .A(n12706), .Z(n12701) );
  BUF_X1 U477 ( .A(n12705), .Z(n12700) );
  BUF_X1 U478 ( .A(n12704), .Z(n12699) );
  BUF_X1 U479 ( .A(n12703), .Z(n12698) );
  BUF_X1 U480 ( .A(n12702), .Z(n12697) );
  BUF_X1 U481 ( .A(n12704), .Z(n12696) );
  BUF_X1 U482 ( .A(n12706), .Z(n12695) );
  BUF_X1 U483 ( .A(n12723), .Z(n12717) );
  BUF_X1 U484 ( .A(n12722), .Z(n12716) );
  BUF_X1 U485 ( .A(n12726), .Z(n12715) );
  BUF_X1 U486 ( .A(n12749), .Z(n12746) );
  BUF_X1 U487 ( .A(n12749), .Z(n12745) );
  BUF_X1 U488 ( .A(n12749), .Z(n12744) );
  BUF_X1 U489 ( .A(n12749), .Z(n12743) );
  BUF_X1 U490 ( .A(n12749), .Z(n12742) );
  BUF_X1 U491 ( .A(n12742), .Z(n12741) );
  BUF_X1 U492 ( .A(n12746), .Z(n12740) );
  BUF_X1 U493 ( .A(n12745), .Z(n12739) );
  BUF_X1 U494 ( .A(n12744), .Z(n12738) );
  BUF_X1 U495 ( .A(n12743), .Z(n12737) );
  BUF_X1 U496 ( .A(n12745), .Z(n12736) );
  BUF_X1 U497 ( .A(n12742), .Z(n12735) );
  BUF_X1 U498 ( .A(n12804), .Z(n12798) );
  BUF_X1 U499 ( .A(n12803), .Z(n12797) );
  BUF_X1 U500 ( .A(n12805), .Z(n12796) );
  BUF_X1 U501 ( .A(n12802), .Z(n12795) );
  BUF_X1 U502 ( .A(n12829), .Z(n12826) );
  BUF_X1 U503 ( .A(n12829), .Z(n12825) );
  BUF_X1 U504 ( .A(n12829), .Z(n12824) );
  BUF_X1 U505 ( .A(n12829), .Z(n12823) );
  BUF_X1 U506 ( .A(n12829), .Z(n12822) );
  BUF_X1 U507 ( .A(n12822), .Z(n12821) );
  BUF_X1 U508 ( .A(n12826), .Z(n12820) );
  BUF_X1 U509 ( .A(n12825), .Z(n12819) );
  BUF_X1 U510 ( .A(n12824), .Z(n12818) );
  BUF_X1 U511 ( .A(n12823), .Z(n12817) );
  BUF_X1 U512 ( .A(n12825), .Z(n12816) );
  BUF_X1 U513 ( .A(n12822), .Z(n12815) );
  BUF_X1 U514 ( .A(n12889), .Z(n12884) );
  BUF_X1 U515 ( .A(n12889), .Z(n12883) );
  BUF_X1 U516 ( .A(n12889), .Z(n12882) );
  BUF_X1 U517 ( .A(n12882), .Z(n12881) );
  BUF_X1 U518 ( .A(n12886), .Z(n12880) );
  BUF_X1 U519 ( .A(n12885), .Z(n12879) );
  BUF_X1 U520 ( .A(n12884), .Z(n12878) );
  BUF_X1 U521 ( .A(n12883), .Z(n12877) );
  BUF_X1 U522 ( .A(n12882), .Z(n12876) );
  BUF_X1 U523 ( .A(n12886), .Z(n12875) );
  BUF_X1 U524 ( .A(n12909), .Z(n12906) );
  BUF_X1 U525 ( .A(n12909), .Z(n12905) );
  BUF_X1 U526 ( .A(n12909), .Z(n12904) );
  BUF_X1 U527 ( .A(n12909), .Z(n12903) );
  BUF_X1 U528 ( .A(n12909), .Z(n12902) );
  BUF_X1 U529 ( .A(n12902), .Z(n12901) );
  BUF_X1 U530 ( .A(n12906), .Z(n12900) );
  BUF_X1 U531 ( .A(n12905), .Z(n12899) );
  BUF_X1 U532 ( .A(n12904), .Z(n12898) );
  BUF_X1 U533 ( .A(n12903), .Z(n12897) );
  BUF_X1 U534 ( .A(n12902), .Z(n12896) );
  BUF_X1 U535 ( .A(n12906), .Z(n12895) );
  BUF_X1 U536 ( .A(n12969), .Z(n12964) );
  BUF_X1 U537 ( .A(n12969), .Z(n12963) );
  BUF_X1 U538 ( .A(n12969), .Z(n12962) );
  BUF_X1 U539 ( .A(n12962), .Z(n12961) );
  BUF_X1 U540 ( .A(n12966), .Z(n12960) );
  BUF_X1 U541 ( .A(n12965), .Z(n12959) );
  BUF_X1 U542 ( .A(n12964), .Z(n12958) );
  BUF_X1 U543 ( .A(n12963), .Z(n12957) );
  BUF_X1 U544 ( .A(n12962), .Z(n12956) );
  BUF_X1 U545 ( .A(n12966), .Z(n12955) );
  BUF_X1 U546 ( .A(n12989), .Z(n12986) );
  BUF_X1 U547 ( .A(n12989), .Z(n12985) );
  BUF_X1 U548 ( .A(n12989), .Z(n12984) );
  BUF_X1 U549 ( .A(n12989), .Z(n12983) );
  BUF_X1 U550 ( .A(n12989), .Z(n12982) );
  BUF_X1 U551 ( .A(n12982), .Z(n12981) );
  BUF_X1 U552 ( .A(n12986), .Z(n12980) );
  BUF_X1 U553 ( .A(n12985), .Z(n12979) );
  BUF_X1 U554 ( .A(n12984), .Z(n12978) );
  BUF_X1 U555 ( .A(n12983), .Z(n12977) );
  BUF_X1 U556 ( .A(n12982), .Z(n12976) );
  BUF_X1 U557 ( .A(n12986), .Z(n12975) );
  BUF_X1 U558 ( .A(n13169), .Z(n13166) );
  BUF_X1 U559 ( .A(n13169), .Z(n13165) );
  BUF_X1 U560 ( .A(n13169), .Z(n13164) );
  BUF_X1 U561 ( .A(n13169), .Z(n13163) );
  BUF_X1 U562 ( .A(n13169), .Z(n13162) );
  BUF_X1 U563 ( .A(n13373), .Z(n13367) );
  BUF_X1 U564 ( .A(n13372), .Z(n13366) );
  BUF_X1 U565 ( .A(n13371), .Z(n13365) );
  BUF_X1 U566 ( .A(n13375), .Z(n13364) );
  BUF_X1 U567 ( .A(n13029), .Z(n13027) );
  BUF_X1 U568 ( .A(n13049), .Z(n13047) );
  BUF_X1 U569 ( .A(n13129), .Z(n13127) );
  BUF_X1 U570 ( .A(n13069), .Z(n13067) );
  BUF_X1 U571 ( .A(n12869), .Z(n12867) );
  BUF_X1 U572 ( .A(n13019), .Z(n13025) );
  BUF_X1 U573 ( .A(n13039), .Z(n13045) );
  BUF_X1 U574 ( .A(n12935), .Z(n12946) );
  BUF_X1 U575 ( .A(n13118), .Z(n13125) );
  BUF_X1 U576 ( .A(n13059), .Z(n13065) );
  BUF_X1 U577 ( .A(n12859), .Z(n12865) );
  BUF_X1 U578 ( .A(n13029), .Z(n13028) );
  BUF_X1 U579 ( .A(n13049), .Z(n13048) );
  BUF_X1 U580 ( .A(n12614), .Z(n12613) );
  BUF_X1 U581 ( .A(n12929), .Z(n12928) );
  BUF_X1 U582 ( .A(n12949), .Z(n12948) );
  BUF_X1 U583 ( .A(n13009), .Z(n13008) );
  BUF_X1 U584 ( .A(n13149), .Z(n13148) );
  BUF_X1 U585 ( .A(n13129), .Z(n13128) );
  BUF_X1 U586 ( .A(n13109), .Z(n13108) );
  BUF_X1 U587 ( .A(n13089), .Z(n13088) );
  BUF_X1 U588 ( .A(n13069), .Z(n13068) );
  BUF_X1 U589 ( .A(n12869), .Z(n12868) );
  BUF_X1 U590 ( .A(n12849), .Z(n12848) );
  BUF_X1 U591 ( .A(n12789), .Z(n12788) );
  BUF_X1 U592 ( .A(n12769), .Z(n12768) );
  BUF_X1 U593 ( .A(n12595), .Z(n12594) );
  BUF_X1 U594 ( .A(n12652), .Z(n12651) );
  BUF_X1 U595 ( .A(n12671), .Z(n12670) );
  BUF_X1 U596 ( .A(n12633), .Z(n12632) );
  BUF_X1 U597 ( .A(n12690), .Z(n12689) );
  BUF_X1 U598 ( .A(n12709), .Z(n12708) );
  BUF_X1 U599 ( .A(n12729), .Z(n12728) );
  BUF_X1 U600 ( .A(n12749), .Z(n12748) );
  BUF_X1 U601 ( .A(n12809), .Z(n12808) );
  BUF_X1 U602 ( .A(n12829), .Z(n12828) );
  BUF_X1 U603 ( .A(n12889), .Z(n12888) );
  BUF_X1 U604 ( .A(n12909), .Z(n12908) );
  BUF_X1 U605 ( .A(n12969), .Z(n12968) );
  BUF_X1 U606 ( .A(n12989), .Z(n12988) );
  BUF_X1 U607 ( .A(n13169), .Z(n13168) );
  BUF_X1 U608 ( .A(n13378), .Z(n13377) );
  BUF_X1 U609 ( .A(n12939), .Z(n12945) );
  BUF_X1 U610 ( .A(n13018), .Z(n13026) );
  BUF_X1 U611 ( .A(n13038), .Z(n13046) );
  BUF_X1 U612 ( .A(n12938), .Z(n12943) );
  BUF_X1 U613 ( .A(n13117), .Z(n13126) );
  BUF_X1 U614 ( .A(n13058), .Z(n13066) );
  BUF_X1 U615 ( .A(n12858), .Z(n12866) );
  INV_X1 U616 ( .A(n12550), .ZN(n12574) );
  INV_X1 U617 ( .A(n12550), .ZN(n12575) );
  INV_X1 U618 ( .A(n12550), .ZN(n12576) );
  BUF_X1 U619 ( .A(n1982), .Z(n12435) );
  BUF_X1 U620 ( .A(n1987), .Z(n12411) );
  BUF_X1 U621 ( .A(n1982), .Z(n12436) );
  BUF_X1 U622 ( .A(n1987), .Z(n12412) );
  BUF_X1 U623 ( .A(n1982), .Z(n12437) );
  BUF_X1 U624 ( .A(n1987), .Z(n12413) );
  BUF_X1 U625 ( .A(n1982), .Z(n12438) );
  BUF_X1 U626 ( .A(n1987), .Z(n12414) );
  BUF_X1 U627 ( .A(n1982), .Z(n12439) );
  BUF_X1 U628 ( .A(n1987), .Z(n12415) );
  BUF_X1 U629 ( .A(n1992), .Z(n12387) );
  BUF_X1 U630 ( .A(n1997), .Z(n12363) );
  BUF_X1 U631 ( .A(n1958), .Z(n12531) );
  BUF_X1 U632 ( .A(n1963), .Z(n12507) );
  BUF_X1 U633 ( .A(n1968), .Z(n12483) );
  BUF_X1 U634 ( .A(n1973), .Z(n12459) );
  BUF_X1 U635 ( .A(n1992), .Z(n12388) );
  BUF_X1 U636 ( .A(n1997), .Z(n12364) );
  BUF_X1 U637 ( .A(n1958), .Z(n12532) );
  BUF_X1 U638 ( .A(n1963), .Z(n12508) );
  BUF_X1 U639 ( .A(n1968), .Z(n12484) );
  BUF_X1 U640 ( .A(n1973), .Z(n12460) );
  BUF_X1 U641 ( .A(n1992), .Z(n12389) );
  BUF_X1 U642 ( .A(n1997), .Z(n12365) );
  BUF_X1 U643 ( .A(n1958), .Z(n12533) );
  BUF_X1 U644 ( .A(n1963), .Z(n12509) );
  BUF_X1 U645 ( .A(n1968), .Z(n12485) );
  BUF_X1 U646 ( .A(n1973), .Z(n12461) );
  BUF_X1 U647 ( .A(n1992), .Z(n12390) );
  BUF_X1 U648 ( .A(n1997), .Z(n12366) );
  BUF_X1 U649 ( .A(n1958), .Z(n12534) );
  BUF_X1 U650 ( .A(n1963), .Z(n12510) );
  BUF_X1 U651 ( .A(n1968), .Z(n12486) );
  BUF_X1 U652 ( .A(n1973), .Z(n12462) );
  BUF_X1 U653 ( .A(n1992), .Z(n12391) );
  BUF_X1 U654 ( .A(n1997), .Z(n12367) );
  BUF_X1 U655 ( .A(n1958), .Z(n12535) );
  BUF_X1 U656 ( .A(n1963), .Z(n12511) );
  BUF_X1 U657 ( .A(n1968), .Z(n12487) );
  BUF_X1 U658 ( .A(n1973), .Z(n12463) );
  BUF_X1 U659 ( .A(n1983), .Z(n12429) );
  BUF_X1 U660 ( .A(n1988), .Z(n12405) );
  BUF_X1 U661 ( .A(n1993), .Z(n12381) );
  BUF_X1 U662 ( .A(n1959), .Z(n12525) );
  BUF_X1 U663 ( .A(n1964), .Z(n12501) );
  BUF_X1 U664 ( .A(n1969), .Z(n12477) );
  BUF_X1 U665 ( .A(n1974), .Z(n12453) );
  BUF_X1 U666 ( .A(n1983), .Z(n12430) );
  BUF_X1 U667 ( .A(n1988), .Z(n12406) );
  BUF_X1 U668 ( .A(n1993), .Z(n12382) );
  BUF_X1 U669 ( .A(n1959), .Z(n12526) );
  BUF_X1 U670 ( .A(n1964), .Z(n12502) );
  BUF_X1 U671 ( .A(n1969), .Z(n12478) );
  BUF_X1 U672 ( .A(n1974), .Z(n12454) );
  BUF_X1 U673 ( .A(n1983), .Z(n12431) );
  BUF_X1 U674 ( .A(n1988), .Z(n12407) );
  BUF_X1 U675 ( .A(n1993), .Z(n12383) );
  BUF_X1 U676 ( .A(n1959), .Z(n12527) );
  BUF_X1 U677 ( .A(n1964), .Z(n12503) );
  BUF_X1 U678 ( .A(n1969), .Z(n12479) );
  BUF_X1 U679 ( .A(n1974), .Z(n12455) );
  BUF_X1 U680 ( .A(n1983), .Z(n12432) );
  BUF_X1 U681 ( .A(n1988), .Z(n12408) );
  BUF_X1 U682 ( .A(n1993), .Z(n12384) );
  BUF_X1 U683 ( .A(n1959), .Z(n12528) );
  BUF_X1 U684 ( .A(n1964), .Z(n12504) );
  BUF_X1 U685 ( .A(n1969), .Z(n12480) );
  BUF_X1 U686 ( .A(n1974), .Z(n12456) );
  BUF_X1 U687 ( .A(n1983), .Z(n12433) );
  BUF_X1 U688 ( .A(n1988), .Z(n12409) );
  BUF_X1 U689 ( .A(n1993), .Z(n12385) );
  BUF_X1 U690 ( .A(n1959), .Z(n12529) );
  BUF_X1 U691 ( .A(n1964), .Z(n12505) );
  BUF_X1 U692 ( .A(n1969), .Z(n12481) );
  BUF_X1 U693 ( .A(n1974), .Z(n12457) );
  BUF_X1 U694 ( .A(n1995), .Z(n12375) );
  BUF_X1 U695 ( .A(n2000), .Z(n12351) );
  BUF_X1 U696 ( .A(n1961), .Z(n12519) );
  BUF_X1 U697 ( .A(n1966), .Z(n12495) );
  BUF_X1 U698 ( .A(n1995), .Z(n12376) );
  BUF_X1 U699 ( .A(n2000), .Z(n12352) );
  BUF_X1 U700 ( .A(n1961), .Z(n12520) );
  BUF_X1 U701 ( .A(n1966), .Z(n12496) );
  BUF_X1 U702 ( .A(n1995), .Z(n12377) );
  BUF_X1 U703 ( .A(n2000), .Z(n12353) );
  BUF_X1 U704 ( .A(n1961), .Z(n12521) );
  BUF_X1 U705 ( .A(n1966), .Z(n12497) );
  BUF_X1 U706 ( .A(n1995), .Z(n12378) );
  BUF_X1 U707 ( .A(n2000), .Z(n12354) );
  BUF_X1 U708 ( .A(n1961), .Z(n12522) );
  BUF_X1 U709 ( .A(n1966), .Z(n12498) );
  BUF_X1 U710 ( .A(n1995), .Z(n12379) );
  BUF_X1 U711 ( .A(n2000), .Z(n12355) );
  BUF_X1 U712 ( .A(n1961), .Z(n12523) );
  BUF_X1 U713 ( .A(n1966), .Z(n12499) );
  BUF_X1 U714 ( .A(n1985), .Z(n12423) );
  BUF_X1 U715 ( .A(n1990), .Z(n12399) );
  BUF_X1 U716 ( .A(n1971), .Z(n12471) );
  BUF_X1 U717 ( .A(n1976), .Z(n12447) );
  BUF_X1 U718 ( .A(n1985), .Z(n12424) );
  BUF_X1 U719 ( .A(n1990), .Z(n12400) );
  BUF_X1 U720 ( .A(n1971), .Z(n12472) );
  BUF_X1 U721 ( .A(n1976), .Z(n12448) );
  BUF_X1 U722 ( .A(n1985), .Z(n12425) );
  BUF_X1 U723 ( .A(n1990), .Z(n12401) );
  BUF_X1 U724 ( .A(n1971), .Z(n12473) );
  BUF_X1 U725 ( .A(n1976), .Z(n12449) );
  BUF_X1 U726 ( .A(n1985), .Z(n12426) );
  BUF_X1 U727 ( .A(n1990), .Z(n12402) );
  BUF_X1 U728 ( .A(n1971), .Z(n12474) );
  BUF_X1 U729 ( .A(n1976), .Z(n12450) );
  BUF_X1 U730 ( .A(n1985), .Z(n12427) );
  BUF_X1 U731 ( .A(n1990), .Z(n12403) );
  BUF_X1 U732 ( .A(n1971), .Z(n12475) );
  BUF_X1 U733 ( .A(n1976), .Z(n12451) );
  BUF_X1 U734 ( .A(n1986), .Z(n12417) );
  BUF_X1 U735 ( .A(n1991), .Z(n12393) );
  BUF_X1 U736 ( .A(n1986), .Z(n12418) );
  BUF_X1 U737 ( .A(n1991), .Z(n12394) );
  BUF_X1 U738 ( .A(n1986), .Z(n12419) );
  BUF_X1 U739 ( .A(n1991), .Z(n12395) );
  BUF_X1 U740 ( .A(n1986), .Z(n12420) );
  BUF_X1 U741 ( .A(n1991), .Z(n12396) );
  BUF_X1 U742 ( .A(n1986), .Z(n12421) );
  BUF_X1 U743 ( .A(n1991), .Z(n12397) );
  BUF_X1 U744 ( .A(n1996), .Z(n12369) );
  BUF_X1 U745 ( .A(n2001), .Z(n12345) );
  BUF_X1 U746 ( .A(n1962), .Z(n12513) );
  BUF_X1 U747 ( .A(n1967), .Z(n12489) );
  BUF_X1 U748 ( .A(n1996), .Z(n12370) );
  BUF_X1 U749 ( .A(n2001), .Z(n12346) );
  BUF_X1 U750 ( .A(n1962), .Z(n12514) );
  BUF_X1 U751 ( .A(n1967), .Z(n12490) );
  BUF_X1 U752 ( .A(n1996), .Z(n12371) );
  BUF_X1 U753 ( .A(n2001), .Z(n12347) );
  BUF_X1 U754 ( .A(n1962), .Z(n12515) );
  BUF_X1 U755 ( .A(n1967), .Z(n12491) );
  BUF_X1 U756 ( .A(n1996), .Z(n12372) );
  BUF_X1 U757 ( .A(n2001), .Z(n12348) );
  BUF_X1 U758 ( .A(n1962), .Z(n12516) );
  BUF_X1 U759 ( .A(n1967), .Z(n12492) );
  BUF_X1 U760 ( .A(n1996), .Z(n12373) );
  BUF_X1 U761 ( .A(n2001), .Z(n12349) );
  BUF_X1 U762 ( .A(n1962), .Z(n12517) );
  BUF_X1 U763 ( .A(n1967), .Z(n12493) );
  BUF_X1 U764 ( .A(n1972), .Z(n12465) );
  BUF_X1 U765 ( .A(n1977), .Z(n12441) );
  BUF_X1 U766 ( .A(n1972), .Z(n12466) );
  BUF_X1 U767 ( .A(n1977), .Z(n12442) );
  BUF_X1 U768 ( .A(n1972), .Z(n12467) );
  BUF_X1 U769 ( .A(n1977), .Z(n12443) );
  BUF_X1 U770 ( .A(n1972), .Z(n12468) );
  BUF_X1 U771 ( .A(n1977), .Z(n12444) );
  BUF_X1 U772 ( .A(n1972), .Z(n12469) );
  BUF_X1 U773 ( .A(n1977), .Z(n12445) );
  AND2_X1 U774 ( .A1(n3209), .A2(n3194), .ZN(n1998) );
  BUF_X1 U775 ( .A(n1949), .Z(n12550) );
  INV_X1 U776 ( .A(n13030), .ZN(n13049) );
  INV_X1 U777 ( .A(n13010), .ZN(n13029) );
  INV_X1 U778 ( .A(n12577), .ZN(n12595) );
  INV_X1 U779 ( .A(n12910), .ZN(n12929) );
  INV_X1 U780 ( .A(n12830), .ZN(n12849) );
  INV_X1 U781 ( .A(n12790), .ZN(n12809) );
  INV_X1 U782 ( .A(n12770), .ZN(n12789) );
  INV_X1 U783 ( .A(n12750), .ZN(n12769) );
  INV_X1 U784 ( .A(n12710), .ZN(n12729) );
  INV_X1 U785 ( .A(n12730), .ZN(n12749) );
  INV_X1 U786 ( .A(n12810), .ZN(n12829) );
  INV_X1 U787 ( .A(n12850), .ZN(n12869) );
  INV_X1 U788 ( .A(n13359), .ZN(n13378) );
  INV_X1 U789 ( .A(n13130), .ZN(n13149) );
  INV_X1 U790 ( .A(n13090), .ZN(n13109) );
  INV_X1 U791 ( .A(n13070), .ZN(n13089) );
  INV_X1 U792 ( .A(n13150), .ZN(n13169) );
  INV_X1 U793 ( .A(n13110), .ZN(n13129) );
  INV_X1 U794 ( .A(n13050), .ZN(n13069) );
  INV_X1 U795 ( .A(n12990), .ZN(n13009) );
  INV_X1 U796 ( .A(n12930), .ZN(n12949) );
  INV_X1 U797 ( .A(n12634), .ZN(n12652) );
  INV_X1 U798 ( .A(n12653), .ZN(n12671) );
  INV_X1 U799 ( .A(n12672), .ZN(n12690) );
  INV_X1 U800 ( .A(n12596), .ZN(n12614) );
  INV_X1 U801 ( .A(n12615), .ZN(n12633) );
  INV_X1 U802 ( .A(n12691), .ZN(n12709) );
  INV_X1 U803 ( .A(n12870), .ZN(n12889) );
  INV_X1 U804 ( .A(n12890), .ZN(n12909) );
  INV_X1 U805 ( .A(n12950), .ZN(n12969) );
  INV_X1 U806 ( .A(n12970), .ZN(n12989) );
  BUF_X1 U807 ( .A(n3259), .Z(n12152) );
  BUF_X1 U808 ( .A(n3259), .Z(n12153) );
  BUF_X1 U809 ( .A(n3259), .Z(n12154) );
  BUF_X1 U810 ( .A(n3259), .Z(n12155) );
  BUF_X1 U811 ( .A(n3259), .Z(n12156) );
  NOR2_X1 U812 ( .A1(n14463), .A2(n14464), .ZN(n3194) );
  NOR3_X1 U813 ( .A1(n14465), .A2(n14461), .A3(n14462), .ZN(n3209) );
  NAND2_X1 U814 ( .A1(n3189), .A2(n3205), .ZN(n1985) );
  NAND2_X1 U815 ( .A1(n3193), .A2(n3205), .ZN(n1990) );
  NAND2_X1 U816 ( .A1(n3208), .A2(n3189), .ZN(n1996) );
  NAND2_X1 U817 ( .A1(n3190), .A2(n3189), .ZN(n1961) );
  NAND2_X1 U818 ( .A1(n3188), .A2(n3189), .ZN(n1962) );
  NAND2_X1 U819 ( .A1(n3209), .A2(n3193), .ZN(n2000) );
  NAND2_X1 U820 ( .A1(n3208), .A2(n3193), .ZN(n2001) );
  NAND2_X1 U821 ( .A1(n3190), .A2(n3193), .ZN(n1966) );
  NAND2_X1 U822 ( .A1(n3188), .A2(n3193), .ZN(n1967) );
  NAND2_X1 U823 ( .A1(n3197), .A2(n3194), .ZN(n1976) );
  NAND2_X1 U824 ( .A1(n3196), .A2(n3194), .ZN(n1977) );
  NAND2_X1 U825 ( .A1(n3197), .A2(n3191), .ZN(n1971) );
  NAND2_X1 U826 ( .A1(n3196), .A2(n3191), .ZN(n1972) );
  OAI21_X1 U827 ( .B1(n1921), .B2(n1942), .A(n12137), .ZN(n1949) );
  AND2_X1 U828 ( .A1(n3205), .A2(n3191), .ZN(n1983) );
  AND2_X1 U829 ( .A1(n3194), .A2(n3205), .ZN(n1988) );
  AND2_X1 U830 ( .A1(n3208), .A2(n3191), .ZN(n1992) );
  AND2_X1 U831 ( .A1(n3208), .A2(n3194), .ZN(n1997) );
  AND2_X1 U832 ( .A1(n3188), .A2(n3191), .ZN(n1958) );
  AND2_X1 U833 ( .A1(n3190), .A2(n3191), .ZN(n1959) );
  AND2_X1 U834 ( .A1(n3188), .A2(n3194), .ZN(n1963) );
  AND2_X1 U835 ( .A1(n3190), .A2(n3194), .ZN(n1964) );
  AND2_X1 U836 ( .A1(n3196), .A2(n3189), .ZN(n1968) );
  AND2_X1 U837 ( .A1(n3197), .A2(n3189), .ZN(n1969) );
  AND2_X1 U838 ( .A1(n3196), .A2(n3193), .ZN(n1973) );
  AND2_X1 U839 ( .A1(n3197), .A2(n3193), .ZN(n1974) );
  AND2_X1 U840 ( .A1(n3209), .A2(n3191), .ZN(n1993) );
  OAI21_X1 U841 ( .B1(n1919), .B2(n1942), .A(n12137), .ZN(n1948) );
  OAI21_X1 U842 ( .B1(n1913), .B2(n1942), .A(n12137), .ZN(n1945) );
  OAI21_X1 U843 ( .B1(n1911), .B2(n1942), .A(n12137), .ZN(n1944) );
  OAI21_X1 U844 ( .B1(n1917), .B2(n1942), .A(n12137), .ZN(n1947) );
  OAI21_X1 U845 ( .B1(n1915), .B2(n1942), .A(n12137), .ZN(n1946) );
  OAI21_X1 U846 ( .B1(n1909), .B2(n1942), .A(n12137), .ZN(n1943) );
  OAI21_X1 U847 ( .B1(n1907), .B2(n1942), .A(n12137), .ZN(n1941) );
  OAI21_X1 U848 ( .B1(n1917), .B2(n1924), .A(n12138), .ZN(n1929) );
  OAI21_X1 U849 ( .B1(n1921), .B2(n1924), .A(n12138), .ZN(n1931) );
  OAI21_X1 U850 ( .B1(n1919), .B2(n1924), .A(n12138), .ZN(n1930) );
  OAI21_X1 U851 ( .B1(n1913), .B2(n1924), .A(n12138), .ZN(n1927) );
  OAI21_X1 U852 ( .B1(n1911), .B2(n1924), .A(n12139), .ZN(n1926) );
  BUF_X1 U853 ( .A(n3219), .Z(n12326) );
  BUF_X1 U854 ( .A(n3224), .Z(n12302) );
  BUF_X1 U855 ( .A(n3229), .Z(n12278) );
  BUF_X1 U856 ( .A(n3234), .Z(n12254) );
  BUF_X1 U857 ( .A(n3243), .Z(n12230) );
  BUF_X1 U858 ( .A(n3248), .Z(n12206) );
  BUF_X1 U859 ( .A(n3253), .Z(n12182) );
  BUF_X1 U860 ( .A(n3258), .Z(n12158) );
  BUF_X1 U861 ( .A(n3219), .Z(n12327) );
  BUF_X1 U862 ( .A(n3224), .Z(n12303) );
  BUF_X1 U863 ( .A(n3229), .Z(n12279) );
  BUF_X1 U864 ( .A(n3234), .Z(n12255) );
  BUF_X1 U865 ( .A(n3243), .Z(n12231) );
  BUF_X1 U866 ( .A(n3248), .Z(n12207) );
  BUF_X1 U867 ( .A(n3253), .Z(n12183) );
  BUF_X1 U868 ( .A(n3258), .Z(n12159) );
  BUF_X1 U869 ( .A(n3219), .Z(n12328) );
  BUF_X1 U870 ( .A(n3224), .Z(n12304) );
  BUF_X1 U871 ( .A(n3229), .Z(n12280) );
  BUF_X1 U872 ( .A(n3234), .Z(n12256) );
  BUF_X1 U873 ( .A(n3243), .Z(n12232) );
  BUF_X1 U874 ( .A(n3248), .Z(n12208) );
  BUF_X1 U875 ( .A(n3253), .Z(n12184) );
  BUF_X1 U876 ( .A(n3258), .Z(n12160) );
  BUF_X1 U877 ( .A(n3219), .Z(n12329) );
  BUF_X1 U878 ( .A(n3224), .Z(n12305) );
  BUF_X1 U879 ( .A(n3229), .Z(n12281) );
  BUF_X1 U880 ( .A(n3234), .Z(n12257) );
  BUF_X1 U881 ( .A(n3243), .Z(n12233) );
  BUF_X1 U882 ( .A(n3248), .Z(n12209) );
  BUF_X1 U883 ( .A(n3253), .Z(n12185) );
  BUF_X1 U884 ( .A(n3258), .Z(n12161) );
  BUF_X1 U885 ( .A(n3219), .Z(n12330) );
  BUF_X1 U886 ( .A(n3224), .Z(n12306) );
  BUF_X1 U887 ( .A(n3229), .Z(n12282) );
  BUF_X1 U888 ( .A(n3234), .Z(n12258) );
  BUF_X1 U889 ( .A(n3243), .Z(n12234) );
  BUF_X1 U890 ( .A(n3248), .Z(n12210) );
  BUF_X1 U891 ( .A(n3253), .Z(n12186) );
  BUF_X1 U892 ( .A(n3258), .Z(n12162) );
  BUF_X1 U893 ( .A(n3220), .Z(n12320) );
  BUF_X1 U894 ( .A(n3225), .Z(n12296) );
  BUF_X1 U895 ( .A(n3230), .Z(n12272) );
  BUF_X1 U896 ( .A(n3235), .Z(n12248) );
  BUF_X1 U897 ( .A(n3244), .Z(n12224) );
  BUF_X1 U898 ( .A(n3249), .Z(n12200) );
  BUF_X1 U899 ( .A(n3254), .Z(n12176) );
  BUF_X1 U900 ( .A(n3220), .Z(n12321) );
  BUF_X1 U901 ( .A(n3225), .Z(n12297) );
  BUF_X1 U902 ( .A(n3230), .Z(n12273) );
  BUF_X1 U903 ( .A(n3235), .Z(n12249) );
  BUF_X1 U904 ( .A(n3244), .Z(n12225) );
  BUF_X1 U905 ( .A(n3249), .Z(n12201) );
  BUF_X1 U906 ( .A(n3254), .Z(n12177) );
  BUF_X1 U907 ( .A(n3220), .Z(n12322) );
  BUF_X1 U908 ( .A(n3225), .Z(n12298) );
  BUF_X1 U909 ( .A(n3230), .Z(n12274) );
  BUF_X1 U910 ( .A(n3235), .Z(n12250) );
  BUF_X1 U911 ( .A(n3244), .Z(n12226) );
  BUF_X1 U912 ( .A(n3249), .Z(n12202) );
  BUF_X1 U913 ( .A(n3254), .Z(n12178) );
  BUF_X1 U914 ( .A(n3220), .Z(n12323) );
  BUF_X1 U915 ( .A(n3225), .Z(n12299) );
  BUF_X1 U916 ( .A(n3230), .Z(n12275) );
  BUF_X1 U917 ( .A(n3235), .Z(n12251) );
  BUF_X1 U918 ( .A(n3244), .Z(n12227) );
  BUF_X1 U919 ( .A(n3249), .Z(n12203) );
  BUF_X1 U920 ( .A(n3254), .Z(n12179) );
  BUF_X1 U921 ( .A(n3220), .Z(n12324) );
  BUF_X1 U922 ( .A(n3225), .Z(n12300) );
  BUF_X1 U923 ( .A(n3230), .Z(n12276) );
  BUF_X1 U924 ( .A(n3235), .Z(n12252) );
  BUF_X1 U925 ( .A(n3244), .Z(n12228) );
  BUF_X1 U926 ( .A(n3249), .Z(n12204) );
  BUF_X1 U927 ( .A(n3254), .Z(n12180) );
  BUF_X1 U928 ( .A(n3222), .Z(n12314) );
  BUF_X1 U929 ( .A(n3227), .Z(n12290) );
  BUF_X1 U930 ( .A(n3256), .Z(n12170) );
  BUF_X1 U931 ( .A(n3261), .Z(n12146) );
  BUF_X1 U932 ( .A(n3222), .Z(n12315) );
  BUF_X1 U933 ( .A(n3227), .Z(n12291) );
  BUF_X1 U934 ( .A(n3256), .Z(n12171) );
  BUF_X1 U935 ( .A(n3261), .Z(n12147) );
  BUF_X1 U936 ( .A(n3222), .Z(n12316) );
  BUF_X1 U937 ( .A(n3227), .Z(n12292) );
  BUF_X1 U938 ( .A(n3256), .Z(n12172) );
  BUF_X1 U939 ( .A(n3261), .Z(n12148) );
  BUF_X1 U940 ( .A(n3222), .Z(n12317) );
  BUF_X1 U941 ( .A(n3227), .Z(n12293) );
  BUF_X1 U942 ( .A(n3256), .Z(n12173) );
  BUF_X1 U943 ( .A(n3261), .Z(n12149) );
  BUF_X1 U944 ( .A(n3222), .Z(n12318) );
  BUF_X1 U945 ( .A(n3227), .Z(n12294) );
  BUF_X1 U946 ( .A(n3256), .Z(n12174) );
  BUF_X1 U947 ( .A(n3261), .Z(n12150) );
  BUF_X1 U948 ( .A(n3232), .Z(n12266) );
  BUF_X1 U949 ( .A(n3246), .Z(n12218) );
  BUF_X1 U950 ( .A(n3251), .Z(n12194) );
  BUF_X1 U951 ( .A(n3232), .Z(n12267) );
  BUF_X1 U952 ( .A(n3246), .Z(n12219) );
  BUF_X1 U953 ( .A(n3251), .Z(n12195) );
  BUF_X1 U954 ( .A(n3232), .Z(n12268) );
  BUF_X1 U955 ( .A(n3246), .Z(n12220) );
  BUF_X1 U956 ( .A(n3251), .Z(n12196) );
  BUF_X1 U957 ( .A(n3232), .Z(n12269) );
  BUF_X1 U958 ( .A(n3246), .Z(n12221) );
  BUF_X1 U959 ( .A(n3251), .Z(n12197) );
  BUF_X1 U960 ( .A(n3232), .Z(n12270) );
  BUF_X1 U961 ( .A(n3246), .Z(n12222) );
  BUF_X1 U962 ( .A(n3251), .Z(n12198) );
  BUF_X1 U963 ( .A(n3237), .Z(n12242) );
  BUF_X1 U964 ( .A(n3237), .Z(n12243) );
  BUF_X1 U965 ( .A(n3237), .Z(n12244) );
  BUF_X1 U966 ( .A(n3237), .Z(n12245) );
  BUF_X1 U967 ( .A(n3237), .Z(n12246) );
  BUF_X1 U968 ( .A(n3223), .Z(n12308) );
  BUF_X1 U969 ( .A(n3228), .Z(n12284) );
  BUF_X1 U970 ( .A(n3257), .Z(n12164) );
  BUF_X1 U971 ( .A(n3262), .Z(n12140) );
  BUF_X1 U972 ( .A(n3223), .Z(n12309) );
  BUF_X1 U973 ( .A(n3228), .Z(n12285) );
  BUF_X1 U974 ( .A(n3257), .Z(n12165) );
  BUF_X1 U975 ( .A(n3262), .Z(n12141) );
  BUF_X1 U976 ( .A(n3223), .Z(n12310) );
  BUF_X1 U977 ( .A(n3228), .Z(n12286) );
  BUF_X1 U978 ( .A(n3257), .Z(n12166) );
  BUF_X1 U979 ( .A(n3262), .Z(n12142) );
  BUF_X1 U980 ( .A(n3223), .Z(n12311) );
  BUF_X1 U981 ( .A(n3228), .Z(n12287) );
  BUF_X1 U982 ( .A(n3257), .Z(n12167) );
  BUF_X1 U983 ( .A(n3262), .Z(n12143) );
  BUF_X1 U984 ( .A(n3223), .Z(n12312) );
  BUF_X1 U985 ( .A(n3228), .Z(n12288) );
  BUF_X1 U986 ( .A(n3257), .Z(n12168) );
  BUF_X1 U987 ( .A(n3262), .Z(n12144) );
  BUF_X1 U988 ( .A(n3233), .Z(n12260) );
  BUF_X1 U989 ( .A(n3247), .Z(n12212) );
  BUF_X1 U990 ( .A(n3252), .Z(n12188) );
  BUF_X1 U991 ( .A(n3233), .Z(n12261) );
  BUF_X1 U992 ( .A(n3247), .Z(n12213) );
  BUF_X1 U993 ( .A(n3252), .Z(n12189) );
  BUF_X1 U994 ( .A(n3233), .Z(n12262) );
  BUF_X1 U995 ( .A(n3247), .Z(n12214) );
  BUF_X1 U996 ( .A(n3252), .Z(n12190) );
  BUF_X1 U997 ( .A(n3233), .Z(n12263) );
  BUF_X1 U998 ( .A(n3247), .Z(n12215) );
  BUF_X1 U999 ( .A(n3252), .Z(n12191) );
  BUF_X1 U1000 ( .A(n3233), .Z(n12264) );
  BUF_X1 U1001 ( .A(n3247), .Z(n12216) );
  BUF_X1 U1002 ( .A(n3252), .Z(n12192) );
  BUF_X1 U1003 ( .A(n3238), .Z(n12236) );
  BUF_X1 U1004 ( .A(n3238), .Z(n12237) );
  BUF_X1 U1005 ( .A(n3238), .Z(n12238) );
  BUF_X1 U1006 ( .A(n3238), .Z(n12239) );
  BUF_X1 U1007 ( .A(n3238), .Z(n12240) );
  BUF_X1 U1008 ( .A(n12332), .Z(n12338) );
  BUF_X1 U1009 ( .A(n12332), .Z(n12337) );
  BUF_X1 U1010 ( .A(n12332), .Z(n12335) );
  BUF_X1 U1011 ( .A(n12332), .Z(n12334) );
  BUF_X1 U1012 ( .A(n12332), .Z(n12336) );
  BUF_X1 U1013 ( .A(n12332), .Z(n12339) );
  BUF_X1 U1014 ( .A(n12333), .Z(n12340) );
  BUF_X1 U1015 ( .A(n12333), .Z(n12341) );
  BUF_X1 U1016 ( .A(n12333), .Z(n12342) );
  BUF_X1 U1017 ( .A(n12333), .Z(n12343) );
  AND2_X1 U1018 ( .A1(n4470), .A2(n4455), .ZN(n3259) );
  BUF_X1 U1019 ( .A(n12130), .Z(n12137) );
  BUF_X1 U1020 ( .A(n12130), .Z(n12136) );
  BUF_X1 U1021 ( .A(n12129), .Z(n12134) );
  BUF_X1 U1022 ( .A(n12130), .Z(n12135) );
  BUF_X1 U1023 ( .A(n12129), .Z(n12133) );
  BUF_X1 U1024 ( .A(n12129), .Z(n12132) );
  BUF_X1 U1025 ( .A(n12537), .Z(n12543) );
  BUF_X1 U1026 ( .A(n12537), .Z(n12542) );
  BUF_X1 U1027 ( .A(n12537), .Z(n12540) );
  BUF_X1 U1028 ( .A(n12537), .Z(n12539) );
  BUF_X1 U1029 ( .A(n12537), .Z(n12541) );
  BUF_X1 U1030 ( .A(n12537), .Z(n12544) );
  BUF_X1 U1031 ( .A(n12538), .Z(n12545) );
  BUF_X1 U1032 ( .A(n12538), .Z(n12546) );
  BUF_X1 U1033 ( .A(n12538), .Z(n12547) );
  BUF_X1 U1034 ( .A(n12538), .Z(n12548) );
  BUF_X1 U1035 ( .A(n12131), .Z(n12138) );
  BUF_X1 U1036 ( .A(n12131), .Z(n12139) );
  NOR2_X1 U1037 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n3189) );
  NOR2_X1 U1038 ( .A1(n14463), .A2(ADD_RD1[1]), .ZN(n3193) );
  NOR3_X1 U1039 ( .A1(n14461), .A2(ADD_RD1[3]), .A3(n14465), .ZN(n3205) );
  NOR2_X1 U1040 ( .A1(n14464), .A2(ADD_RD1[2]), .ZN(n3191) );
  NOR3_X1 U1041 ( .A1(n14461), .A2(ADD_RD1[0]), .A3(n14462), .ZN(n3208) );
  NOR3_X1 U1042 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n14465), .ZN(n3188) );
  NOR3_X1 U1043 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(n3190) );
  NOR3_X1 U1044 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n14462), .ZN(n3196) );
  NOR3_X1 U1045 ( .A1(n14465), .A2(ADD_RD1[4]), .A3(n14462), .ZN(n3197) );
  AOI221_X1 U1046 ( .B1(n12507), .B2(n11586), .C1(n12501), .C2(n11406), .A(
        n3192), .ZN(n3185) );
  OAI22_X1 U1047 ( .A1(n14362), .A2(n12495), .B1(n14361), .B2(n12489), .ZN(
        n3192) );
  AOI221_X1 U1048 ( .B1(n12507), .B2(n11762), .C1(n12501), .C2(n11582), .A(
        n3169), .ZN(n3166) );
  OAI22_X1 U1049 ( .A1(n14408), .A2(n12495), .B1(n14385), .B2(n12489), .ZN(
        n3169) );
  AOI221_X1 U1050 ( .B1(n12507), .B2(n11587), .C1(n12501), .C2(n11407), .A(
        n3150), .ZN(n3147) );
  OAI22_X1 U1051 ( .A1(n14407), .A2(n12495), .B1(n14384), .B2(n12489), .ZN(
        n3150) );
  AOI221_X1 U1052 ( .B1(n12507), .B2(n11588), .C1(n12501), .C2(n11408), .A(
        n3131), .ZN(n3128) );
  OAI22_X1 U1053 ( .A1(n14406), .A2(n12495), .B1(n14383), .B2(n12489), .ZN(
        n3131) );
  AOI221_X1 U1054 ( .B1(n12507), .B2(n11589), .C1(n12501), .C2(n11409), .A(
        n3112), .ZN(n3109) );
  OAI22_X1 U1055 ( .A1(n14405), .A2(n12495), .B1(n14382), .B2(n12489), .ZN(
        n3112) );
  AOI221_X1 U1056 ( .B1(n12507), .B2(n11763), .C1(n12501), .C2(n11583), .A(
        n3093), .ZN(n3090) );
  OAI22_X1 U1057 ( .A1(n14404), .A2(n12495), .B1(n14381), .B2(n12489), .ZN(
        n3093) );
  AOI221_X1 U1058 ( .B1(n12507), .B2(n11764), .C1(n12501), .C2(n11584), .A(
        n3074), .ZN(n3071) );
  OAI22_X1 U1059 ( .A1(n14403), .A2(n12495), .B1(n14380), .B2(n12489), .ZN(
        n3074) );
  AOI221_X1 U1060 ( .B1(n12507), .B2(n11590), .C1(n12501), .C2(n11410), .A(
        n3055), .ZN(n3052) );
  OAI22_X1 U1061 ( .A1(n14402), .A2(n12495), .B1(n14379), .B2(n12489), .ZN(
        n3055) );
  AOI221_X1 U1062 ( .B1(n12507), .B2(n11591), .C1(n12501), .C2(n11411), .A(
        n3036), .ZN(n3033) );
  OAI22_X1 U1063 ( .A1(n14401), .A2(n12495), .B1(n14378), .B2(n12489), .ZN(
        n3036) );
  AOI221_X1 U1064 ( .B1(n12507), .B2(n11592), .C1(n12501), .C2(n11412), .A(
        n3017), .ZN(n3014) );
  OAI22_X1 U1065 ( .A1(n14400), .A2(n12495), .B1(n14377), .B2(n12489), .ZN(
        n3017) );
  AOI221_X1 U1066 ( .B1(n12507), .B2(n11593), .C1(n12501), .C2(n11413), .A(
        n2998), .ZN(n2995) );
  OAI22_X1 U1067 ( .A1(n14399), .A2(n12495), .B1(n14376), .B2(n12489), .ZN(
        n2998) );
  AOI221_X1 U1068 ( .B1(n12507), .B2(n11594), .C1(n12501), .C2(n11414), .A(
        n2979), .ZN(n2976) );
  OAI22_X1 U1069 ( .A1(n14398), .A2(n12495), .B1(n14375), .B2(n12489), .ZN(
        n2979) );
  AOI221_X1 U1070 ( .B1(n12508), .B2(n11595), .C1(n12502), .C2(n11415), .A(
        n2960), .ZN(n2957) );
  OAI22_X1 U1071 ( .A1(n14397), .A2(n12496), .B1(n14374), .B2(n12490), .ZN(
        n2960) );
  AOI221_X1 U1072 ( .B1(n12508), .B2(n11596), .C1(n12502), .C2(n11416), .A(
        n2941), .ZN(n2938) );
  OAI22_X1 U1073 ( .A1(n14396), .A2(n12496), .B1(n14373), .B2(n12490), .ZN(
        n2941) );
  AOI221_X1 U1074 ( .B1(n12508), .B2(n11597), .C1(n12502), .C2(n11417), .A(
        n2922), .ZN(n2919) );
  OAI22_X1 U1075 ( .A1(n14395), .A2(n12496), .B1(n14372), .B2(n12490), .ZN(
        n2922) );
  AOI221_X1 U1076 ( .B1(n12508), .B2(n11598), .C1(n12502), .C2(n11418), .A(
        n2903), .ZN(n2900) );
  OAI22_X1 U1077 ( .A1(n14394), .A2(n12496), .B1(n14371), .B2(n12490), .ZN(
        n2903) );
  AOI221_X1 U1078 ( .B1(n12508), .B2(n11599), .C1(n12502), .C2(n11419), .A(
        n2884), .ZN(n2881) );
  OAI22_X1 U1079 ( .A1(n14393), .A2(n12496), .B1(n14370), .B2(n12490), .ZN(
        n2884) );
  AOI221_X1 U1080 ( .B1(n12508), .B2(n11600), .C1(n12502), .C2(n11420), .A(
        n2865), .ZN(n2862) );
  OAI22_X1 U1081 ( .A1(n14392), .A2(n12496), .B1(n14369), .B2(n12490), .ZN(
        n2865) );
  AOI221_X1 U1082 ( .B1(n12508), .B2(n11601), .C1(n12502), .C2(n11421), .A(
        n2846), .ZN(n2843) );
  OAI22_X1 U1083 ( .A1(n14391), .A2(n12496), .B1(n14368), .B2(n12490), .ZN(
        n2846) );
  AOI221_X1 U1084 ( .B1(n12508), .B2(n11602), .C1(n12502), .C2(n11422), .A(
        n2827), .ZN(n2824) );
  OAI22_X1 U1085 ( .A1(n14390), .A2(n12496), .B1(n14367), .B2(n12490), .ZN(
        n2827) );
  AOI221_X1 U1086 ( .B1(n12508), .B2(n11603), .C1(n12502), .C2(n11423), .A(
        n2808), .ZN(n2805) );
  OAI22_X1 U1087 ( .A1(n14389), .A2(n12496), .B1(n14366), .B2(n12490), .ZN(
        n2808) );
  AOI221_X1 U1088 ( .B1(n12508), .B2(n11604), .C1(n12502), .C2(n11424), .A(
        n2789), .ZN(n2786) );
  OAI22_X1 U1089 ( .A1(n14388), .A2(n12496), .B1(n14365), .B2(n12490), .ZN(
        n2789) );
  AOI221_X1 U1090 ( .B1(n12508), .B2(n11605), .C1(n12502), .C2(n11425), .A(
        n2770), .ZN(n2767) );
  OAI22_X1 U1091 ( .A1(n14387), .A2(n12496), .B1(n14364), .B2(n12490), .ZN(
        n2770) );
  AOI221_X1 U1092 ( .B1(n12508), .B2(n11606), .C1(n12502), .C2(n11426), .A(
        n2751), .ZN(n2748) );
  OAI22_X1 U1093 ( .A1(n14386), .A2(n12496), .B1(n14363), .B2(n12490), .ZN(
        n2751) );
  AOI221_X1 U1094 ( .B1(n12509), .B2(n11607), .C1(n12503), .C2(n11427), .A(
        n2732), .ZN(n2729) );
  OAI22_X1 U1095 ( .A1(n14288), .A2(n12497), .B1(n14252), .B2(n12491), .ZN(
        n2732) );
  AOI221_X1 U1096 ( .B1(n12509), .B2(n11608), .C1(n12503), .C2(n11428), .A(
        n2713), .ZN(n2710) );
  OAI22_X1 U1097 ( .A1(n14287), .A2(n12497), .B1(n14251), .B2(n12491), .ZN(
        n2713) );
  AOI221_X1 U1098 ( .B1(n12509), .B2(n11609), .C1(n12503), .C2(n11429), .A(
        n2694), .ZN(n2691) );
  OAI22_X1 U1099 ( .A1(n14286), .A2(n12497), .B1(n14250), .B2(n12491), .ZN(
        n2694) );
  AOI221_X1 U1100 ( .B1(n12509), .B2(n11610), .C1(n12503), .C2(n11430), .A(
        n2675), .ZN(n2672) );
  OAI22_X1 U1101 ( .A1(n14285), .A2(n12497), .B1(n14249), .B2(n12491), .ZN(
        n2675) );
  AOI221_X1 U1102 ( .B1(n12509), .B2(n11611), .C1(n12503), .C2(n11431), .A(
        n2656), .ZN(n2653) );
  OAI22_X1 U1103 ( .A1(n14284), .A2(n12497), .B1(n14248), .B2(n12491), .ZN(
        n2656) );
  AOI221_X1 U1104 ( .B1(n12509), .B2(n11612), .C1(n12503), .C2(n11432), .A(
        n2637), .ZN(n2634) );
  OAI22_X1 U1105 ( .A1(n14283), .A2(n12497), .B1(n14247), .B2(n12491), .ZN(
        n2637) );
  AOI221_X1 U1106 ( .B1(n12509), .B2(n11613), .C1(n12503), .C2(n11433), .A(
        n2618), .ZN(n2615) );
  OAI22_X1 U1107 ( .A1(n14282), .A2(n12497), .B1(n14246), .B2(n12491), .ZN(
        n2618) );
  AOI221_X1 U1108 ( .B1(n12509), .B2(n11614), .C1(n12503), .C2(n11434), .A(
        n2599), .ZN(n2596) );
  OAI22_X1 U1109 ( .A1(n14281), .A2(n12497), .B1(n14245), .B2(n12491), .ZN(
        n2599) );
  AOI221_X1 U1110 ( .B1(n12509), .B2(n11615), .C1(n12503), .C2(n11435), .A(
        n2580), .ZN(n2577) );
  OAI22_X1 U1111 ( .A1(n14280), .A2(n12497), .B1(n14244), .B2(n12491), .ZN(
        n2580) );
  AOI221_X1 U1112 ( .B1(n12509), .B2(n11616), .C1(n12503), .C2(n11436), .A(
        n2561), .ZN(n2558) );
  OAI22_X1 U1113 ( .A1(n14279), .A2(n12497), .B1(n14243), .B2(n12491), .ZN(
        n2561) );
  AOI221_X1 U1114 ( .B1(n12509), .B2(n11617), .C1(n12503), .C2(n11437), .A(
        n2542), .ZN(n2539) );
  OAI22_X1 U1115 ( .A1(n14278), .A2(n12497), .B1(n14242), .B2(n12491), .ZN(
        n2542) );
  AOI221_X1 U1116 ( .B1(n12509), .B2(n11618), .C1(n12503), .C2(n11438), .A(
        n2523), .ZN(n2520) );
  OAI22_X1 U1117 ( .A1(n14277), .A2(n12497), .B1(n14241), .B2(n12491), .ZN(
        n2523) );
  AOI221_X1 U1118 ( .B1(n12510), .B2(n11619), .C1(n12504), .C2(n11439), .A(
        n2504), .ZN(n2501) );
  OAI22_X1 U1119 ( .A1(n14276), .A2(n12498), .B1(n14240), .B2(n12492), .ZN(
        n2504) );
  AOI221_X1 U1120 ( .B1(n12510), .B2(n11620), .C1(n12504), .C2(n11440), .A(
        n2485), .ZN(n2482) );
  OAI22_X1 U1121 ( .A1(n14275), .A2(n12498), .B1(n14239), .B2(n12492), .ZN(
        n2485) );
  AOI221_X1 U1122 ( .B1(n12510), .B2(n11621), .C1(n12504), .C2(n11441), .A(
        n2466), .ZN(n2463) );
  OAI22_X1 U1123 ( .A1(n14274), .A2(n12498), .B1(n14238), .B2(n12492), .ZN(
        n2466) );
  AOI221_X1 U1124 ( .B1(n12510), .B2(n11622), .C1(n12504), .C2(n11442), .A(
        n2447), .ZN(n2444) );
  OAI22_X1 U1125 ( .A1(n14273), .A2(n12498), .B1(n14237), .B2(n12492), .ZN(
        n2447) );
  AOI221_X1 U1126 ( .B1(n12510), .B2(n11623), .C1(n12504), .C2(n11443), .A(
        n2428), .ZN(n2425) );
  OAI22_X1 U1127 ( .A1(n14272), .A2(n12498), .B1(n14236), .B2(n12492), .ZN(
        n2428) );
  AOI221_X1 U1128 ( .B1(n12510), .B2(n11624), .C1(n12504), .C2(n11444), .A(
        n2409), .ZN(n2406) );
  OAI22_X1 U1129 ( .A1(n14271), .A2(n12498), .B1(n14235), .B2(n12492), .ZN(
        n2409) );
  AOI221_X1 U1130 ( .B1(n12510), .B2(n11625), .C1(n12504), .C2(n11445), .A(
        n2390), .ZN(n2387) );
  OAI22_X1 U1131 ( .A1(n14270), .A2(n12498), .B1(n14234), .B2(n12492), .ZN(
        n2390) );
  AOI221_X1 U1132 ( .B1(n12510), .B2(n11626), .C1(n12504), .C2(n11446), .A(
        n2371), .ZN(n2368) );
  OAI22_X1 U1133 ( .A1(n14269), .A2(n12498), .B1(n14233), .B2(n12492), .ZN(
        n2371) );
  AOI221_X1 U1134 ( .B1(n12510), .B2(n11627), .C1(n12504), .C2(n11447), .A(
        n2352), .ZN(n2349) );
  OAI22_X1 U1135 ( .A1(n14268), .A2(n12498), .B1(n14232), .B2(n12492), .ZN(
        n2352) );
  AOI221_X1 U1136 ( .B1(n12510), .B2(n11628), .C1(n12504), .C2(n11448), .A(
        n2333), .ZN(n2330) );
  OAI22_X1 U1137 ( .A1(n14267), .A2(n12498), .B1(n14231), .B2(n12492), .ZN(
        n2333) );
  AOI221_X1 U1138 ( .B1(n12510), .B2(n11629), .C1(n12504), .C2(n11449), .A(
        n2314), .ZN(n2311) );
  OAI22_X1 U1139 ( .A1(n14266), .A2(n12498), .B1(n14230), .B2(n12492), .ZN(
        n2314) );
  AOI221_X1 U1140 ( .B1(n12510), .B2(n11630), .C1(n12504), .C2(n11450), .A(
        n2295), .ZN(n2292) );
  OAI22_X1 U1141 ( .A1(n14265), .A2(n12498), .B1(n14229), .B2(n12492), .ZN(
        n2295) );
  AOI221_X1 U1142 ( .B1(n12511), .B2(n11631), .C1(n12505), .C2(n11451), .A(
        n2276), .ZN(n2273) );
  OAI22_X1 U1143 ( .A1(n14264), .A2(n12499), .B1(n14228), .B2(n12493), .ZN(
        n2276) );
  AOI221_X1 U1144 ( .B1(n12511), .B2(n11632), .C1(n12505), .C2(n11452), .A(
        n2257), .ZN(n2254) );
  OAI22_X1 U1145 ( .A1(n14263), .A2(n12499), .B1(n14227), .B2(n12493), .ZN(
        n2257) );
  AOI221_X1 U1146 ( .B1(n12511), .B2(n11633), .C1(n12505), .C2(n11453), .A(
        n2238), .ZN(n2235) );
  OAI22_X1 U1147 ( .A1(n14262), .A2(n12499), .B1(n14226), .B2(n12493), .ZN(
        n2238) );
  AOI221_X1 U1148 ( .B1(n12511), .B2(n11634), .C1(n12505), .C2(n11454), .A(
        n2219), .ZN(n2216) );
  OAI22_X1 U1149 ( .A1(n14261), .A2(n12499), .B1(n14225), .B2(n12493), .ZN(
        n2219) );
  AOI221_X1 U1150 ( .B1(n12511), .B2(n11635), .C1(n12505), .C2(n11455), .A(
        n2200), .ZN(n2197) );
  OAI22_X1 U1151 ( .A1(n14260), .A2(n12499), .B1(n14224), .B2(n12493), .ZN(
        n2200) );
  AOI221_X1 U1152 ( .B1(n12511), .B2(n11636), .C1(n12505), .C2(n11456), .A(
        n2181), .ZN(n2178) );
  OAI22_X1 U1153 ( .A1(n14259), .A2(n12499), .B1(n14223), .B2(n12493), .ZN(
        n2181) );
  AOI221_X1 U1154 ( .B1(n12511), .B2(n11637), .C1(n12505), .C2(n11457), .A(
        n2162), .ZN(n2159) );
  OAI22_X1 U1155 ( .A1(n14258), .A2(n12499), .B1(n14222), .B2(n12493), .ZN(
        n2162) );
  AOI221_X1 U1156 ( .B1(n12511), .B2(n11638), .C1(n12505), .C2(n11458), .A(
        n2143), .ZN(n2140) );
  OAI22_X1 U1157 ( .A1(n14257), .A2(n12499), .B1(n14221), .B2(n12493), .ZN(
        n2143) );
  AOI221_X1 U1158 ( .B1(n12511), .B2(n11639), .C1(n12505), .C2(n11459), .A(
        n2124), .ZN(n2121) );
  OAI22_X1 U1159 ( .A1(n14256), .A2(n12499), .B1(n14220), .B2(n12493), .ZN(
        n2124) );
  AOI221_X1 U1160 ( .B1(n12511), .B2(n11640), .C1(n12505), .C2(n11460), .A(
        n2105), .ZN(n2102) );
  OAI22_X1 U1161 ( .A1(n14255), .A2(n12499), .B1(n14219), .B2(n12493), .ZN(
        n2105) );
  AOI221_X1 U1162 ( .B1(n12511), .B2(n11641), .C1(n12505), .C2(n11461), .A(
        n2086), .ZN(n2083) );
  OAI22_X1 U1163 ( .A1(n14254), .A2(n12499), .B1(n14218), .B2(n12493), .ZN(
        n2086) );
  AOI221_X1 U1164 ( .B1(n12511), .B2(n11765), .C1(n12505), .C2(n11585), .A(
        n2067), .ZN(n2064) );
  OAI22_X1 U1165 ( .A1(n14253), .A2(n12499), .B1(n14217), .B2(n12493), .ZN(
        n2067) );
  AOI221_X1 U1166 ( .B1(n12512), .B2(n13835), .C1(n12506), .C2(n13839), .A(
        n2048), .ZN(n2045) );
  OAI22_X1 U1167 ( .A1(n13847), .A2(n12500), .B1(n13843), .B2(n12494), .ZN(
        n2048) );
  AOI221_X1 U1168 ( .B1(n12512), .B2(n13834), .C1(n12506), .C2(n13838), .A(
        n2029), .ZN(n2026) );
  OAI22_X1 U1169 ( .A1(n13846), .A2(n12500), .B1(n13842), .B2(n12494), .ZN(
        n2029) );
  AOI221_X1 U1170 ( .B1(n12512), .B2(n13833), .C1(n12506), .C2(n13837), .A(
        n2010), .ZN(n2007) );
  OAI22_X1 U1171 ( .A1(n13845), .A2(n12500), .B1(n13841), .B2(n12494), .ZN(
        n2010) );
  AOI221_X1 U1172 ( .B1(n12512), .B2(n13832), .C1(n12506), .C2(n13836), .A(
        n1965), .ZN(n1956) );
  OAI22_X1 U1173 ( .A1(n13844), .A2(n12500), .B1(n13840), .B2(n12494), .ZN(
        n1965) );
  AOI221_X1 U1174 ( .B1(n12387), .B2(n14153), .C1(n12381), .C2(n14154), .A(
        n3207), .ZN(n3200) );
  OAI22_X1 U1175 ( .A1(n13746), .A2(n12375), .B1(n13730), .B2(n12369), .ZN(
        n3207) );
  AOI221_X1 U1176 ( .B1(n12483), .B2(n11642), .C1(n12477), .C2(n11462), .A(
        n3195), .ZN(n3184) );
  OAI22_X1 U1177 ( .A1(n13539), .A2(n12471), .B1(n13494), .B2(n12465), .ZN(
        n3195) );
  AOI221_X1 U1178 ( .B1(n12387), .B2(n14082), .C1(n12381), .C2(n14129), .A(
        n3178), .ZN(n3173) );
  OAI22_X1 U1179 ( .A1(n13745), .A2(n12375), .B1(n13729), .B2(n12369), .ZN(
        n3178) );
  AOI221_X1 U1180 ( .B1(n12483), .B2(n11643), .C1(n12477), .C2(n11463), .A(
        n3170), .ZN(n3165) );
  OAI22_X1 U1181 ( .A1(n13538), .A2(n12471), .B1(n13493), .B2(n12465), .ZN(
        n3170) );
  AOI221_X1 U1182 ( .B1(n12387), .B2(n14081), .C1(n12381), .C2(n14128), .A(
        n3159), .ZN(n3154) );
  OAI22_X1 U1183 ( .A1(n13744), .A2(n12375), .B1(n13728), .B2(n12369), .ZN(
        n3159) );
  AOI221_X1 U1184 ( .B1(n12483), .B2(n11644), .C1(n12477), .C2(n11464), .A(
        n3151), .ZN(n3146) );
  OAI22_X1 U1185 ( .A1(n13537), .A2(n12471), .B1(n13492), .B2(n12465), .ZN(
        n3151) );
  AOI221_X1 U1186 ( .B1(n12483), .B2(n11645), .C1(n12477), .C2(n11465), .A(
        n3132), .ZN(n3127) );
  OAI22_X1 U1187 ( .A1(n13536), .A2(n12471), .B1(n13491), .B2(n12465), .ZN(
        n3132) );
  AOI221_X1 U1188 ( .B1(n12483), .B2(n11646), .C1(n12477), .C2(n11466), .A(
        n3113), .ZN(n3108) );
  OAI22_X1 U1189 ( .A1(n14360), .A2(n12471), .B1(n13490), .B2(n12465), .ZN(
        n3113) );
  AOI221_X1 U1190 ( .B1(n12387), .B2(n14078), .C1(n12381), .C2(n14125), .A(
        n3102), .ZN(n3097) );
  OAI22_X1 U1191 ( .A1(n13891), .A2(n12375), .B1(n13725), .B2(n12369), .ZN(
        n3102) );
  AOI221_X1 U1192 ( .B1(n12483), .B2(n11647), .C1(n12477), .C2(n11467), .A(
        n3094), .ZN(n3089) );
  OAI22_X1 U1193 ( .A1(n14359), .A2(n12471), .B1(n13489), .B2(n12465), .ZN(
        n3094) );
  AOI221_X1 U1194 ( .B1(n12387), .B2(n14077), .C1(n12381), .C2(n14124), .A(
        n3083), .ZN(n3078) );
  OAI22_X1 U1195 ( .A1(n13890), .A2(n12375), .B1(n13724), .B2(n12369), .ZN(
        n3083) );
  AOI221_X1 U1196 ( .B1(n12483), .B2(n11648), .C1(n12477), .C2(n11468), .A(
        n3075), .ZN(n3070) );
  OAI22_X1 U1197 ( .A1(n14358), .A2(n12471), .B1(n13488), .B2(n12465), .ZN(
        n3075) );
  AOI221_X1 U1198 ( .B1(n12483), .B2(n11649), .C1(n12477), .C2(n11469), .A(
        n3056), .ZN(n3051) );
  OAI22_X1 U1199 ( .A1(n14340), .A2(n12471), .B1(n13487), .B2(n12465), .ZN(
        n3056) );
  AOI221_X1 U1200 ( .B1(n12483), .B2(n11650), .C1(n12477), .C2(n11470), .A(
        n3037), .ZN(n3032) );
  OAI22_X1 U1201 ( .A1(n14339), .A2(n12471), .B1(n13486), .B2(n12465), .ZN(
        n3037) );
  AOI221_X1 U1202 ( .B1(n12483), .B2(n11651), .C1(n12477), .C2(n11471), .A(
        n3018), .ZN(n3013) );
  OAI22_X1 U1203 ( .A1(n14338), .A2(n12471), .B1(n13485), .B2(n12465), .ZN(
        n3018) );
  AOI221_X1 U1204 ( .B1(n12483), .B2(n11652), .C1(n12477), .C2(n11472), .A(
        n2999), .ZN(n2994) );
  OAI22_X1 U1205 ( .A1(n14337), .A2(n12471), .B1(n13484), .B2(n12465), .ZN(
        n2999) );
  AOI221_X1 U1206 ( .B1(n12483), .B2(n11653), .C1(n12477), .C2(n11473), .A(
        n2980), .ZN(n2975) );
  OAI22_X1 U1207 ( .A1(n14336), .A2(n12471), .B1(n13483), .B2(n12465), .ZN(
        n2980) );
  AOI221_X1 U1208 ( .B1(n12484), .B2(n11654), .C1(n12478), .C2(n11474), .A(
        n2961), .ZN(n2956) );
  OAI22_X1 U1209 ( .A1(n14335), .A2(n12472), .B1(n13482), .B2(n12466), .ZN(
        n2961) );
  AOI221_X1 U1210 ( .B1(n12484), .B2(n11655), .C1(n12478), .C2(n11475), .A(
        n2942), .ZN(n2937) );
  OAI22_X1 U1211 ( .A1(n14334), .A2(n12472), .B1(n13481), .B2(n12466), .ZN(
        n2942) );
  AOI221_X1 U1212 ( .B1(n12484), .B2(n11656), .C1(n12478), .C2(n11476), .A(
        n2923), .ZN(n2918) );
  OAI22_X1 U1213 ( .A1(n14333), .A2(n12472), .B1(n13480), .B2(n12466), .ZN(
        n2923) );
  AOI221_X1 U1214 ( .B1(n12484), .B2(n11657), .C1(n12478), .C2(n11477), .A(
        n2904), .ZN(n2899) );
  OAI22_X1 U1215 ( .A1(n14332), .A2(n12472), .B1(n13479), .B2(n12466), .ZN(
        n2904) );
  AOI221_X1 U1216 ( .B1(n12484), .B2(n11658), .C1(n12478), .C2(n11478), .A(
        n2885), .ZN(n2880) );
  OAI22_X1 U1217 ( .A1(n13535), .A2(n12472), .B1(n13478), .B2(n12466), .ZN(
        n2885) );
  AOI221_X1 U1218 ( .B1(n12484), .B2(n11659), .C1(n12478), .C2(n11479), .A(
        n2866), .ZN(n2861) );
  OAI22_X1 U1219 ( .A1(n14331), .A2(n12472), .B1(n13477), .B2(n12466), .ZN(
        n2866) );
  AOI221_X1 U1220 ( .B1(n12484), .B2(n11660), .C1(n12478), .C2(n11480), .A(
        n2847), .ZN(n2842) );
  OAI22_X1 U1221 ( .A1(n14330), .A2(n12472), .B1(n13476), .B2(n12466), .ZN(
        n2847) );
  AOI221_X1 U1222 ( .B1(n12484), .B2(n11661), .C1(n12478), .C2(n11481), .A(
        n2828), .ZN(n2823) );
  OAI22_X1 U1223 ( .A1(n14329), .A2(n12472), .B1(n13475), .B2(n12466), .ZN(
        n2828) );
  AOI221_X1 U1224 ( .B1(n12484), .B2(n11662), .C1(n12478), .C2(n11482), .A(
        n2809), .ZN(n2804) );
  OAI22_X1 U1225 ( .A1(n13534), .A2(n12472), .B1(n13474), .B2(n12466), .ZN(
        n2809) );
  AOI221_X1 U1226 ( .B1(n12484), .B2(n11663), .C1(n12478), .C2(n11483), .A(
        n2790), .ZN(n2785) );
  OAI22_X1 U1227 ( .A1(n13533), .A2(n12472), .B1(n13473), .B2(n12466), .ZN(
        n2790) );
  AOI221_X1 U1228 ( .B1(n12484), .B2(n11664), .C1(n12478), .C2(n11484), .A(
        n2771), .ZN(n2766) );
  OAI22_X1 U1229 ( .A1(n13532), .A2(n12472), .B1(n13472), .B2(n12466), .ZN(
        n2771) );
  AOI221_X1 U1230 ( .B1(n12484), .B2(n11665), .C1(n12478), .C2(n11485), .A(
        n2752), .ZN(n2747) );
  OAI22_X1 U1231 ( .A1(n13531), .A2(n12472), .B1(n13471), .B2(n12466), .ZN(
        n2752) );
  AOI221_X1 U1232 ( .B1(n12485), .B2(n11666), .C1(n12479), .C2(n11486), .A(
        n2733), .ZN(n2728) );
  OAI22_X1 U1233 ( .A1(n13530), .A2(n12473), .B1(n13470), .B2(n12467), .ZN(
        n2733) );
  AOI221_X1 U1234 ( .B1(n12485), .B2(n11667), .C1(n12479), .C2(n11487), .A(
        n2714), .ZN(n2709) );
  OAI22_X1 U1235 ( .A1(n13529), .A2(n12473), .B1(n13469), .B2(n12467), .ZN(
        n2714) );
  AOI221_X1 U1236 ( .B1(n12485), .B2(n11668), .C1(n12479), .C2(n11488), .A(
        n2695), .ZN(n2690) );
  OAI22_X1 U1237 ( .A1(n13528), .A2(n12473), .B1(n13468), .B2(n12467), .ZN(
        n2695) );
  AOI221_X1 U1238 ( .B1(n12485), .B2(n11669), .C1(n12479), .C2(n11489), .A(
        n2676), .ZN(n2671) );
  OAI22_X1 U1239 ( .A1(n13527), .A2(n12473), .B1(n13467), .B2(n12467), .ZN(
        n2676) );
  AOI221_X1 U1240 ( .B1(n12485), .B2(n11670), .C1(n12479), .C2(n11490), .A(
        n2657), .ZN(n2652) );
  OAI22_X1 U1241 ( .A1(n13526), .A2(n12473), .B1(n13466), .B2(n12467), .ZN(
        n2657) );
  AOI221_X1 U1242 ( .B1(n12485), .B2(n11671), .C1(n12479), .C2(n11491), .A(
        n2638), .ZN(n2633) );
  OAI22_X1 U1243 ( .A1(n13525), .A2(n12473), .B1(n13465), .B2(n12467), .ZN(
        n2638) );
  AOI221_X1 U1244 ( .B1(n12485), .B2(n11672), .C1(n12479), .C2(n11492), .A(
        n2619), .ZN(n2614) );
  OAI22_X1 U1245 ( .A1(n13524), .A2(n12473), .B1(n13464), .B2(n12467), .ZN(
        n2619) );
  AOI221_X1 U1246 ( .B1(n12485), .B2(n11673), .C1(n12479), .C2(n11493), .A(
        n2600), .ZN(n2595) );
  OAI22_X1 U1247 ( .A1(n13523), .A2(n12473), .B1(n13463), .B2(n12467), .ZN(
        n2600) );
  AOI221_X1 U1248 ( .B1(n12485), .B2(n11674), .C1(n12479), .C2(n11494), .A(
        n2581), .ZN(n2576) );
  OAI22_X1 U1249 ( .A1(n13522), .A2(n12473), .B1(n13462), .B2(n12467), .ZN(
        n2581) );
  AOI221_X1 U1250 ( .B1(n12485), .B2(n11675), .C1(n12479), .C2(n11495), .A(
        n2562), .ZN(n2557) );
  OAI22_X1 U1251 ( .A1(n13521), .A2(n12473), .B1(n13461), .B2(n12467), .ZN(
        n2562) );
  AOI221_X1 U1252 ( .B1(n12485), .B2(n11676), .C1(n12479), .C2(n11496), .A(
        n2543), .ZN(n2538) );
  OAI22_X1 U1253 ( .A1(n13520), .A2(n12473), .B1(n13460), .B2(n12467), .ZN(
        n2543) );
  AOI221_X1 U1254 ( .B1(n12485), .B2(n11677), .C1(n12479), .C2(n11497), .A(
        n2524), .ZN(n2519) );
  OAI22_X1 U1255 ( .A1(n13519), .A2(n12473), .B1(n13459), .B2(n12467), .ZN(
        n2524) );
  AOI221_X1 U1256 ( .B1(n12486), .B2(n11678), .C1(n12480), .C2(n11498), .A(
        n2505), .ZN(n2500) );
  OAI22_X1 U1257 ( .A1(n13518), .A2(n12474), .B1(n13458), .B2(n12468), .ZN(
        n2505) );
  AOI221_X1 U1258 ( .B1(n12486), .B2(n11679), .C1(n12480), .C2(n11499), .A(
        n2486), .ZN(n2481) );
  OAI22_X1 U1259 ( .A1(n13517), .A2(n12474), .B1(n13457), .B2(n12468), .ZN(
        n2486) );
  AOI221_X1 U1260 ( .B1(n12486), .B2(n11680), .C1(n12480), .C2(n11500), .A(
        n2467), .ZN(n2462) );
  OAI22_X1 U1261 ( .A1(n13516), .A2(n12474), .B1(n13456), .B2(n12468), .ZN(
        n2467) );
  AOI221_X1 U1262 ( .B1(n12486), .B2(n11681), .C1(n12480), .C2(n11501), .A(
        n2448), .ZN(n2443) );
  OAI22_X1 U1263 ( .A1(n14460), .A2(n12474), .B1(n13455), .B2(n12468), .ZN(
        n2448) );
  AOI221_X1 U1264 ( .B1(n12486), .B2(n11682), .C1(n12480), .C2(n11502), .A(
        n2429), .ZN(n2424) );
  OAI22_X1 U1265 ( .A1(n14459), .A2(n12474), .B1(n13454), .B2(n12468), .ZN(
        n2429) );
  AOI221_X1 U1266 ( .B1(n12486), .B2(n11683), .C1(n12480), .C2(n11503), .A(
        n2410), .ZN(n2405) );
  OAI22_X1 U1267 ( .A1(n14458), .A2(n12474), .B1(n13453), .B2(n12468), .ZN(
        n2410) );
  AOI221_X1 U1268 ( .B1(n12486), .B2(n11684), .C1(n12480), .C2(n11504), .A(
        n2391), .ZN(n2386) );
  OAI22_X1 U1269 ( .A1(n14457), .A2(n12474), .B1(n13452), .B2(n12468), .ZN(
        n2391) );
  AOI221_X1 U1270 ( .B1(n12486), .B2(n11685), .C1(n12480), .C2(n11505), .A(
        n2372), .ZN(n2367) );
  OAI22_X1 U1271 ( .A1(n13515), .A2(n12474), .B1(n13451), .B2(n12468), .ZN(
        n2372) );
  AOI221_X1 U1272 ( .B1(n12486), .B2(n11686), .C1(n12480), .C2(n11506), .A(
        n2353), .ZN(n2348) );
  OAI22_X1 U1273 ( .A1(n13514), .A2(n12474), .B1(n13450), .B2(n12468), .ZN(
        n2353) );
  AOI221_X1 U1274 ( .B1(n12486), .B2(n11687), .C1(n12480), .C2(n11507), .A(
        n2334), .ZN(n2329) );
  OAI22_X1 U1275 ( .A1(n13513), .A2(n12474), .B1(n13449), .B2(n12468), .ZN(
        n2334) );
  AOI221_X1 U1276 ( .B1(n12486), .B2(n11688), .C1(n12480), .C2(n11508), .A(
        n2315), .ZN(n2310) );
  OAI22_X1 U1277 ( .A1(n13512), .A2(n12474), .B1(n13448), .B2(n12468), .ZN(
        n2315) );
  AOI221_X1 U1278 ( .B1(n12486), .B2(n11689), .C1(n12480), .C2(n11509), .A(
        n2296), .ZN(n2291) );
  OAI22_X1 U1279 ( .A1(n13511), .A2(n12474), .B1(n13447), .B2(n12468), .ZN(
        n2296) );
  AOI221_X1 U1280 ( .B1(n12487), .B2(n11690), .C1(n12481), .C2(n11510), .A(
        n2277), .ZN(n2272) );
  OAI22_X1 U1281 ( .A1(n13510), .A2(n12475), .B1(n13446), .B2(n12469), .ZN(
        n2277) );
  AOI221_X1 U1282 ( .B1(n12487), .B2(n11691), .C1(n12481), .C2(n11511), .A(
        n2258), .ZN(n2253) );
  OAI22_X1 U1283 ( .A1(n13509), .A2(n12475), .B1(n13445), .B2(n12469), .ZN(
        n2258) );
  AOI221_X1 U1284 ( .B1(n12487), .B2(n11692), .C1(n12481), .C2(n11512), .A(
        n2239), .ZN(n2234) );
  OAI22_X1 U1285 ( .A1(n13508), .A2(n12475), .B1(n13444), .B2(n12469), .ZN(
        n2239) );
  AOI221_X1 U1286 ( .B1(n12487), .B2(n11693), .C1(n12481), .C2(n11513), .A(
        n2220), .ZN(n2215) );
  OAI22_X1 U1287 ( .A1(n13507), .A2(n12475), .B1(n13443), .B2(n12469), .ZN(
        n2220) );
  AOI221_X1 U1288 ( .B1(n12487), .B2(n11694), .C1(n12481), .C2(n11514), .A(
        n2201), .ZN(n2196) );
  OAI22_X1 U1289 ( .A1(n13506), .A2(n12475), .B1(n13442), .B2(n12469), .ZN(
        n2201) );
  AOI221_X1 U1290 ( .B1(n12487), .B2(n11695), .C1(n12481), .C2(n11515), .A(
        n2182), .ZN(n2177) );
  OAI22_X1 U1291 ( .A1(n13505), .A2(n12475), .B1(n13441), .B2(n12469), .ZN(
        n2182) );
  AOI221_X1 U1292 ( .B1(n12487), .B2(n11696), .C1(n12481), .C2(n11516), .A(
        n2163), .ZN(n2158) );
  OAI22_X1 U1293 ( .A1(n13504), .A2(n12475), .B1(n13440), .B2(n12469), .ZN(
        n2163) );
  AOI221_X1 U1294 ( .B1(n12487), .B2(n11697), .C1(n12481), .C2(n11517), .A(
        n2144), .ZN(n2139) );
  OAI22_X1 U1295 ( .A1(n13503), .A2(n12475), .B1(n13439), .B2(n12469), .ZN(
        n2144) );
  AOI221_X1 U1296 ( .B1(n12487), .B2(n11698), .C1(n12481), .C2(n11518), .A(
        n2125), .ZN(n2120) );
  OAI22_X1 U1297 ( .A1(n13502), .A2(n12475), .B1(n13438), .B2(n12469), .ZN(
        n2125) );
  AOI221_X1 U1298 ( .B1(n12487), .B2(n11699), .C1(n12481), .C2(n11519), .A(
        n2106), .ZN(n2101) );
  OAI22_X1 U1299 ( .A1(n13501), .A2(n12475), .B1(n13437), .B2(n12469), .ZN(
        n2106) );
  AOI221_X1 U1300 ( .B1(n12487), .B2(n11700), .C1(n12481), .C2(n11520), .A(
        n2087), .ZN(n2082) );
  OAI22_X1 U1301 ( .A1(n13500), .A2(n12475), .B1(n13436), .B2(n12469), .ZN(
        n2087) );
  AOI221_X1 U1302 ( .B1(n12391), .B2(n13893), .C1(n12385), .C2(n13953), .A(
        n2076), .ZN(n2071) );
  OAI22_X1 U1303 ( .A1(n13735), .A2(n12379), .B1(n13671), .B2(n12373), .ZN(
        n2076) );
  AOI221_X1 U1304 ( .B1(n12487), .B2(n11701), .C1(n12481), .C2(n11521), .A(
        n2068), .ZN(n2063) );
  OAI22_X1 U1305 ( .A1(n13499), .A2(n12475), .B1(n13435), .B2(n12469), .ZN(
        n2068) );
  AOI221_X1 U1306 ( .B1(n12392), .B2(n13819), .C1(n12386), .C2(n13823), .A(
        n2057), .ZN(n2052) );
  OAI22_X1 U1307 ( .A1(n13734), .A2(n12380), .B1(n13670), .B2(n12374), .ZN(
        n2057) );
  AOI221_X1 U1308 ( .B1(n12488), .B2(n13860), .C1(n12482), .C2(n13856), .A(
        n2049), .ZN(n2044) );
  OAI22_X1 U1309 ( .A1(n13498), .A2(n12476), .B1(n13434), .B2(n12470), .ZN(
        n2049) );
  AOI221_X1 U1310 ( .B1(n12392), .B2(n13818), .C1(n12386), .C2(n13822), .A(
        n2038), .ZN(n2033) );
  OAI22_X1 U1311 ( .A1(n13733), .A2(n12380), .B1(n13669), .B2(n12374), .ZN(
        n2038) );
  AOI221_X1 U1312 ( .B1(n12488), .B2(n13859), .C1(n12482), .C2(n13855), .A(
        n2030), .ZN(n2025) );
  OAI22_X1 U1313 ( .A1(n13497), .A2(n12476), .B1(n13433), .B2(n12470), .ZN(
        n2030) );
  AOI221_X1 U1314 ( .B1(n12392), .B2(n13817), .C1(n12386), .C2(n13821), .A(
        n2019), .ZN(n2014) );
  OAI22_X1 U1315 ( .A1(n13732), .A2(n12380), .B1(n13668), .B2(n12374), .ZN(
        n2019) );
  AOI221_X1 U1316 ( .B1(n12488), .B2(n13858), .C1(n12482), .C2(n13854), .A(
        n2011), .ZN(n2006) );
  OAI22_X1 U1317 ( .A1(n13496), .A2(n12476), .B1(n13432), .B2(n12470), .ZN(
        n2011) );
  AOI221_X1 U1318 ( .B1(n12392), .B2(n13816), .C1(n12386), .C2(n13820), .A(
        n1994), .ZN(n1979) );
  OAI22_X1 U1319 ( .A1(n13731), .A2(n12380), .B1(n13667), .B2(n12374), .ZN(
        n1994) );
  AOI221_X1 U1320 ( .B1(n12488), .B2(n13857), .C1(n12482), .C2(n13853), .A(
        n1970), .ZN(n1955) );
  OAI22_X1 U1321 ( .A1(n13495), .A2(n12476), .B1(n13431), .B2(n12470), .ZN(
        n1970) );
  AOI221_X1 U1322 ( .B1(n12363), .B2(n14155), .C1(n12357), .C2(n13831), .A(
        n3210), .ZN(n3199) );
  OAI22_X1 U1323 ( .A1(n13815), .A2(n12351), .B1(n13810), .B2(n12345), .ZN(
        n3210) );
  AOI221_X1 U1324 ( .B1(n12459), .B2(n11702), .C1(n12453), .C2(n11522), .A(
        n3198), .ZN(n3183) );
  OAI22_X1 U1325 ( .A1(n13650), .A2(n12447), .B1(n13603), .B2(n12441), .ZN(
        n3198) );
  AOI221_X1 U1326 ( .B1(n12363), .B2(n14152), .C1(n12357), .C2(n13830), .A(
        n3179), .ZN(n3172) );
  OAI22_X1 U1327 ( .A1(n13814), .A2(n12351), .B1(n13809), .B2(n12345), .ZN(
        n3179) );
  AOI221_X1 U1328 ( .B1(n12459), .B2(n11703), .C1(n12453), .C2(n11523), .A(
        n3171), .ZN(n3164) );
  OAI22_X1 U1329 ( .A1(n13649), .A2(n12447), .B1(n13602), .B2(n12441), .ZN(
        n3171) );
  AOI221_X1 U1330 ( .B1(n12363), .B2(n14151), .C1(n12357), .C2(n13829), .A(
        n3160), .ZN(n3153) );
  OAI22_X1 U1331 ( .A1(n13813), .A2(n12351), .B1(n13808), .B2(n12345), .ZN(
        n3160) );
  AOI221_X1 U1332 ( .B1(n12459), .B2(n11704), .C1(n12453), .C2(n11524), .A(
        n3152), .ZN(n3145) );
  OAI22_X1 U1333 ( .A1(n13648), .A2(n12447), .B1(n13601), .B2(n12441), .ZN(
        n3152) );
  AOI221_X1 U1334 ( .B1(n12363), .B2(n14149), .C1(n12357), .C2(n13828), .A(
        n3141), .ZN(n3134) );
  OAI22_X1 U1335 ( .A1(n13812), .A2(n12351), .B1(n13807), .B2(n12345), .ZN(
        n3141) );
  AOI221_X1 U1336 ( .B1(n12459), .B2(n11705), .C1(n12453), .C2(n11525), .A(
        n3133), .ZN(n3126) );
  OAI22_X1 U1337 ( .A1(n13647), .A2(n12447), .B1(n13600), .B2(n12441), .ZN(
        n3133) );
  AOI221_X1 U1338 ( .B1(n12363), .B2(n14150), .C1(n12357), .C2(n14215), .A(
        n3122), .ZN(n3115) );
  OAI22_X1 U1339 ( .A1(n13811), .A2(n12351), .B1(n13806), .B2(n12345), .ZN(
        n3122) );
  AOI221_X1 U1340 ( .B1(n12459), .B2(n11706), .C1(n12453), .C2(n11526), .A(
        n3114), .ZN(n3107) );
  OAI22_X1 U1341 ( .A1(n14357), .A2(n12447), .B1(n13599), .B2(n12441), .ZN(
        n3114) );
  AOI221_X1 U1342 ( .B1(n12363), .B2(n14148), .C1(n12357), .C2(n14214), .A(
        n3103), .ZN(n3096) );
  OAI22_X1 U1343 ( .A1(n14035), .A2(n12351), .B1(n13805), .B2(n12345), .ZN(
        n3103) );
  AOI221_X1 U1344 ( .B1(n12459), .B2(n11707), .C1(n12453), .C2(n11527), .A(
        n3095), .ZN(n3088) );
  OAI22_X1 U1345 ( .A1(n14356), .A2(n12447), .B1(n13598), .B2(n12441), .ZN(
        n3095) );
  AOI221_X1 U1346 ( .B1(n12363), .B2(n14147), .C1(n12357), .C2(n14213), .A(
        n3084), .ZN(n3077) );
  OAI22_X1 U1347 ( .A1(n14034), .A2(n12351), .B1(n13804), .B2(n12345), .ZN(
        n3084) );
  AOI221_X1 U1348 ( .B1(n12459), .B2(n11708), .C1(n12453), .C2(n11528), .A(
        n3076), .ZN(n3069) );
  OAI22_X1 U1349 ( .A1(n14355), .A2(n12447), .B1(n13597), .B2(n12441), .ZN(
        n3076) );
  AOI221_X1 U1350 ( .B1(n12363), .B2(n14146), .C1(n12357), .C2(n14212), .A(
        n3065), .ZN(n3058) );
  OAI22_X1 U1351 ( .A1(n14033), .A2(n12351), .B1(n13803), .B2(n12345), .ZN(
        n3065) );
  AOI221_X1 U1352 ( .B1(n12459), .B2(n11709), .C1(n12453), .C2(n11529), .A(
        n3057), .ZN(n3050) );
  OAI22_X1 U1353 ( .A1(n14354), .A2(n12447), .B1(n13596), .B2(n12441), .ZN(
        n3057) );
  AOI221_X1 U1354 ( .B1(n12363), .B2(n14145), .C1(n12357), .C2(n14211), .A(
        n3046), .ZN(n3039) );
  OAI22_X1 U1355 ( .A1(n14032), .A2(n12351), .B1(n13802), .B2(n12345), .ZN(
        n3046) );
  AOI221_X1 U1356 ( .B1(n12459), .B2(n11710), .C1(n12453), .C2(n11530), .A(
        n3038), .ZN(n3031) );
  OAI22_X1 U1357 ( .A1(n14353), .A2(n12447), .B1(n13595), .B2(n12441), .ZN(
        n3038) );
  AOI221_X1 U1358 ( .B1(n12363), .B2(n14144), .C1(n12357), .C2(n14210), .A(
        n3027), .ZN(n3020) );
  OAI22_X1 U1359 ( .A1(n14031), .A2(n12351), .B1(n13801), .B2(n12345), .ZN(
        n3027) );
  AOI221_X1 U1360 ( .B1(n12459), .B2(n11711), .C1(n12453), .C2(n11531), .A(
        n3019), .ZN(n3012) );
  OAI22_X1 U1361 ( .A1(n14352), .A2(n12447), .B1(n13594), .B2(n12441), .ZN(
        n3019) );
  AOI221_X1 U1362 ( .B1(n12363), .B2(n14143), .C1(n12357), .C2(n14209), .A(
        n3008), .ZN(n3001) );
  OAI22_X1 U1363 ( .A1(n14030), .A2(n12351), .B1(n13800), .B2(n12345), .ZN(
        n3008) );
  AOI221_X1 U1364 ( .B1(n12459), .B2(n11712), .C1(n12453), .C2(n11532), .A(
        n3000), .ZN(n2993) );
  OAI22_X1 U1365 ( .A1(n14351), .A2(n12447), .B1(n13593), .B2(n12441), .ZN(
        n3000) );
  AOI221_X1 U1366 ( .B1(n12363), .B2(n14142), .C1(n12357), .C2(n14208), .A(
        n2989), .ZN(n2982) );
  OAI22_X1 U1367 ( .A1(n14029), .A2(n12351), .B1(n13799), .B2(n12345), .ZN(
        n2989) );
  AOI221_X1 U1368 ( .B1(n12459), .B2(n11713), .C1(n12453), .C2(n11533), .A(
        n2981), .ZN(n2974) );
  OAI22_X1 U1369 ( .A1(n14350), .A2(n12447), .B1(n13592), .B2(n12441), .ZN(
        n2981) );
  AOI221_X1 U1370 ( .B1(n12364), .B2(n14141), .C1(n12358), .C2(n14207), .A(
        n2970), .ZN(n2963) );
  OAI22_X1 U1371 ( .A1(n14028), .A2(n12352), .B1(n13798), .B2(n12346), .ZN(
        n2970) );
  AOI221_X1 U1372 ( .B1(n12460), .B2(n11714), .C1(n12454), .C2(n11534), .A(
        n2962), .ZN(n2955) );
  OAI22_X1 U1373 ( .A1(n14349), .A2(n12448), .B1(n13591), .B2(n12442), .ZN(
        n2962) );
  AOI221_X1 U1374 ( .B1(n12364), .B2(n14140), .C1(n12358), .C2(n14206), .A(
        n2951), .ZN(n2944) );
  OAI22_X1 U1375 ( .A1(n14027), .A2(n12352), .B1(n13797), .B2(n12346), .ZN(
        n2951) );
  AOI221_X1 U1376 ( .B1(n12460), .B2(n11715), .C1(n12454), .C2(n11535), .A(
        n2943), .ZN(n2936) );
  OAI22_X1 U1377 ( .A1(n14348), .A2(n12448), .B1(n13590), .B2(n12442), .ZN(
        n2943) );
  AOI221_X1 U1378 ( .B1(n12364), .B2(n14139), .C1(n12358), .C2(n14205), .A(
        n2932), .ZN(n2925) );
  OAI22_X1 U1379 ( .A1(n14026), .A2(n12352), .B1(n13796), .B2(n12346), .ZN(
        n2932) );
  AOI221_X1 U1380 ( .B1(n12460), .B2(n11716), .C1(n12454), .C2(n11536), .A(
        n2924), .ZN(n2917) );
  OAI22_X1 U1381 ( .A1(n14347), .A2(n12448), .B1(n13589), .B2(n12442), .ZN(
        n2924) );
  AOI221_X1 U1382 ( .B1(n12364), .B2(n14138), .C1(n12358), .C2(n14204), .A(
        n2913), .ZN(n2906) );
  OAI22_X1 U1383 ( .A1(n14025), .A2(n12352), .B1(n13795), .B2(n12346), .ZN(
        n2913) );
  AOI221_X1 U1384 ( .B1(n12460), .B2(n11717), .C1(n12454), .C2(n11537), .A(
        n2905), .ZN(n2898) );
  OAI22_X1 U1385 ( .A1(n14346), .A2(n12448), .B1(n13588), .B2(n12442), .ZN(
        n2905) );
  AOI221_X1 U1386 ( .B1(n12364), .B2(n14137), .C1(n12358), .C2(n14203), .A(
        n2894), .ZN(n2887) );
  OAI22_X1 U1387 ( .A1(n13952), .A2(n12352), .B1(n13794), .B2(n12346), .ZN(
        n2894) );
  AOI221_X1 U1388 ( .B1(n12460), .B2(n11718), .C1(n12454), .C2(n11538), .A(
        n2886), .ZN(n2879) );
  OAI22_X1 U1389 ( .A1(n13646), .A2(n12448), .B1(n13587), .B2(n12442), .ZN(
        n2886) );
  AOI221_X1 U1390 ( .B1(n12364), .B2(n14136), .C1(n12358), .C2(n14202), .A(
        n2875), .ZN(n2868) );
  OAI22_X1 U1391 ( .A1(n13951), .A2(n12352), .B1(n13793), .B2(n12346), .ZN(
        n2875) );
  AOI221_X1 U1392 ( .B1(n12460), .B2(n11719), .C1(n12454), .C2(n11539), .A(
        n2867), .ZN(n2860) );
  OAI22_X1 U1393 ( .A1(n14345), .A2(n12448), .B1(n13586), .B2(n12442), .ZN(
        n2867) );
  AOI221_X1 U1394 ( .B1(n12364), .B2(n14135), .C1(n12358), .C2(n14201), .A(
        n2856), .ZN(n2849) );
  OAI22_X1 U1395 ( .A1(n13950), .A2(n12352), .B1(n13792), .B2(n12346), .ZN(
        n2856) );
  AOI221_X1 U1396 ( .B1(n12460), .B2(n11720), .C1(n12454), .C2(n11540), .A(
        n2848), .ZN(n2841) );
  OAI22_X1 U1397 ( .A1(n14344), .A2(n12448), .B1(n13585), .B2(n12442), .ZN(
        n2848) );
  AOI221_X1 U1398 ( .B1(n12364), .B2(n14134), .C1(n12358), .C2(n14200), .A(
        n2837), .ZN(n2830) );
  OAI22_X1 U1399 ( .A1(n13949), .A2(n12352), .B1(n13791), .B2(n12346), .ZN(
        n2837) );
  AOI221_X1 U1400 ( .B1(n12460), .B2(n11721), .C1(n12454), .C2(n11541), .A(
        n2829), .ZN(n2822) );
  OAI22_X1 U1401 ( .A1(n14343), .A2(n12448), .B1(n13584), .B2(n12442), .ZN(
        n2829) );
  AOI221_X1 U1402 ( .B1(n12364), .B2(n14133), .C1(n12358), .C2(n14199), .A(
        n2818), .ZN(n2811) );
  OAI22_X1 U1403 ( .A1(n13948), .A2(n12352), .B1(n13790), .B2(n12346), .ZN(
        n2818) );
  AOI221_X1 U1404 ( .B1(n12460), .B2(n11722), .C1(n12454), .C2(n11542), .A(
        n2810), .ZN(n2803) );
  OAI22_X1 U1405 ( .A1(n14342), .A2(n12448), .B1(n13583), .B2(n12442), .ZN(
        n2810) );
  AOI221_X1 U1406 ( .B1(n12364), .B2(n14132), .C1(n12358), .C2(n14198), .A(
        n2799), .ZN(n2792) );
  OAI22_X1 U1407 ( .A1(n13947), .A2(n12352), .B1(n13789), .B2(n12346), .ZN(
        n2799) );
  AOI221_X1 U1408 ( .B1(n12460), .B2(n11723), .C1(n12454), .C2(n11543), .A(
        n2791), .ZN(n2784) );
  OAI22_X1 U1409 ( .A1(n14341), .A2(n12448), .B1(n13582), .B2(n12442), .ZN(
        n2791) );
  AOI221_X1 U1410 ( .B1(n12364), .B2(n14131), .C1(n12358), .C2(n14197), .A(
        n2780), .ZN(n2773) );
  OAI22_X1 U1411 ( .A1(n13946), .A2(n12352), .B1(n13788), .B2(n12346), .ZN(
        n2780) );
  AOI221_X1 U1412 ( .B1(n12460), .B2(n11724), .C1(n12454), .C2(n11544), .A(
        n2772), .ZN(n2765) );
  OAI22_X1 U1413 ( .A1(n13645), .A2(n12448), .B1(n13581), .B2(n12442), .ZN(
        n2772) );
  AOI221_X1 U1414 ( .B1(n12364), .B2(n14130), .C1(n12358), .C2(n14196), .A(
        n2761), .ZN(n2754) );
  OAI22_X1 U1415 ( .A1(n13945), .A2(n12352), .B1(n13787), .B2(n12346), .ZN(
        n2761) );
  AOI221_X1 U1416 ( .B1(n12460), .B2(n11725), .C1(n12454), .C2(n11545), .A(
        n2753), .ZN(n2746) );
  OAI22_X1 U1417 ( .A1(n13644), .A2(n12448), .B1(n13580), .B2(n12442), .ZN(
        n2753) );
  AOI221_X1 U1418 ( .B1(n12365), .B2(n14024), .C1(n12359), .C2(n14195), .A(
        n2742), .ZN(n2735) );
  OAI22_X1 U1419 ( .A1(n13944), .A2(n12353), .B1(n13786), .B2(n12347), .ZN(
        n2742) );
  AOI221_X1 U1420 ( .B1(n12461), .B2(n11726), .C1(n12455), .C2(n11546), .A(
        n2734), .ZN(n2727) );
  OAI22_X1 U1421 ( .A1(n13643), .A2(n12449), .B1(n13579), .B2(n12443), .ZN(
        n2734) );
  AOI221_X1 U1422 ( .B1(n12365), .B2(n14023), .C1(n12359), .C2(n14194), .A(
        n2723), .ZN(n2716) );
  OAI22_X1 U1423 ( .A1(n13943), .A2(n12353), .B1(n13785), .B2(n12347), .ZN(
        n2723) );
  AOI221_X1 U1424 ( .B1(n12461), .B2(n11727), .C1(n12455), .C2(n11547), .A(
        n2715), .ZN(n2708) );
  OAI22_X1 U1425 ( .A1(n13642), .A2(n12449), .B1(n13578), .B2(n12443), .ZN(
        n2715) );
  AOI221_X1 U1426 ( .B1(n12365), .B2(n14022), .C1(n12359), .C2(n14193), .A(
        n2704), .ZN(n2697) );
  OAI22_X1 U1427 ( .A1(n13942), .A2(n12353), .B1(n13784), .B2(n12347), .ZN(
        n2704) );
  AOI221_X1 U1428 ( .B1(n12461), .B2(n11728), .C1(n12455), .C2(n11548), .A(
        n2696), .ZN(n2689) );
  OAI22_X1 U1429 ( .A1(n13641), .A2(n12449), .B1(n13577), .B2(n12443), .ZN(
        n2696) );
  AOI221_X1 U1430 ( .B1(n12365), .B2(n14021), .C1(n12359), .C2(n14192), .A(
        n2685), .ZN(n2678) );
  OAI22_X1 U1431 ( .A1(n13941), .A2(n12353), .B1(n13783), .B2(n12347), .ZN(
        n2685) );
  AOI221_X1 U1432 ( .B1(n12461), .B2(n11729), .C1(n12455), .C2(n11549), .A(
        n2677), .ZN(n2670) );
  OAI22_X1 U1433 ( .A1(n13640), .A2(n12449), .B1(n13576), .B2(n12443), .ZN(
        n2677) );
  AOI221_X1 U1434 ( .B1(n12365), .B2(n14020), .C1(n12359), .C2(n14191), .A(
        n2666), .ZN(n2659) );
  OAI22_X1 U1435 ( .A1(n13940), .A2(n12353), .B1(n13782), .B2(n12347), .ZN(
        n2666) );
  AOI221_X1 U1436 ( .B1(n12461), .B2(n11730), .C1(n12455), .C2(n11550), .A(
        n2658), .ZN(n2651) );
  OAI22_X1 U1437 ( .A1(n13639), .A2(n12449), .B1(n13575), .B2(n12443), .ZN(
        n2658) );
  AOI221_X1 U1438 ( .B1(n12365), .B2(n14019), .C1(n12359), .C2(n14190), .A(
        n2647), .ZN(n2640) );
  OAI22_X1 U1439 ( .A1(n13939), .A2(n12353), .B1(n13781), .B2(n12347), .ZN(
        n2647) );
  AOI221_X1 U1440 ( .B1(n12461), .B2(n11731), .C1(n12455), .C2(n11551), .A(
        n2639), .ZN(n2632) );
  OAI22_X1 U1441 ( .A1(n13638), .A2(n12449), .B1(n13574), .B2(n12443), .ZN(
        n2639) );
  AOI221_X1 U1442 ( .B1(n12365), .B2(n14018), .C1(n12359), .C2(n14189), .A(
        n2628), .ZN(n2621) );
  OAI22_X1 U1443 ( .A1(n13938), .A2(n12353), .B1(n13780), .B2(n12347), .ZN(
        n2628) );
  AOI221_X1 U1444 ( .B1(n12461), .B2(n11732), .C1(n12455), .C2(n11552), .A(
        n2620), .ZN(n2613) );
  OAI22_X1 U1445 ( .A1(n13637), .A2(n12449), .B1(n13573), .B2(n12443), .ZN(
        n2620) );
  AOI221_X1 U1446 ( .B1(n12365), .B2(n14017), .C1(n12359), .C2(n14188), .A(
        n2609), .ZN(n2602) );
  OAI22_X1 U1447 ( .A1(n13937), .A2(n12353), .B1(n13779), .B2(n12347), .ZN(
        n2609) );
  AOI221_X1 U1448 ( .B1(n12461), .B2(n11733), .C1(n12455), .C2(n11553), .A(
        n2601), .ZN(n2594) );
  OAI22_X1 U1449 ( .A1(n13636), .A2(n12449), .B1(n13572), .B2(n12443), .ZN(
        n2601) );
  AOI221_X1 U1450 ( .B1(n12365), .B2(n14016), .C1(n12359), .C2(n14187), .A(
        n2590), .ZN(n2583) );
  OAI22_X1 U1451 ( .A1(n13936), .A2(n12353), .B1(n13778), .B2(n12347), .ZN(
        n2590) );
  AOI221_X1 U1452 ( .B1(n12461), .B2(n11734), .C1(n12455), .C2(n11554), .A(
        n2582), .ZN(n2575) );
  OAI22_X1 U1453 ( .A1(n13635), .A2(n12449), .B1(n13571), .B2(n12443), .ZN(
        n2582) );
  AOI221_X1 U1454 ( .B1(n12365), .B2(n14015), .C1(n12359), .C2(n14186), .A(
        n2571), .ZN(n2564) );
  OAI22_X1 U1455 ( .A1(n13935), .A2(n12353), .B1(n13777), .B2(n12347), .ZN(
        n2571) );
  AOI221_X1 U1456 ( .B1(n12461), .B2(n11735), .C1(n12455), .C2(n11555), .A(
        n2563), .ZN(n2556) );
  OAI22_X1 U1457 ( .A1(n13634), .A2(n12449), .B1(n13570), .B2(n12443), .ZN(
        n2563) );
  AOI221_X1 U1458 ( .B1(n12365), .B2(n14014), .C1(n12359), .C2(n14185), .A(
        n2552), .ZN(n2545) );
  OAI22_X1 U1459 ( .A1(n13934), .A2(n12353), .B1(n13776), .B2(n12347), .ZN(
        n2552) );
  AOI221_X1 U1460 ( .B1(n12461), .B2(n11736), .C1(n12455), .C2(n11556), .A(
        n2544), .ZN(n2537) );
  OAI22_X1 U1461 ( .A1(n13633), .A2(n12449), .B1(n13569), .B2(n12443), .ZN(
        n2544) );
  AOI221_X1 U1462 ( .B1(n12365), .B2(n14013), .C1(n12359), .C2(n14184), .A(
        n2533), .ZN(n2526) );
  OAI22_X1 U1463 ( .A1(n13933), .A2(n12353), .B1(n13775), .B2(n12347), .ZN(
        n2533) );
  AOI221_X1 U1464 ( .B1(n12461), .B2(n11737), .C1(n12455), .C2(n11557), .A(
        n2525), .ZN(n2518) );
  OAI22_X1 U1465 ( .A1(n13632), .A2(n12449), .B1(n13568), .B2(n12443), .ZN(
        n2525) );
  AOI221_X1 U1466 ( .B1(n12366), .B2(n14012), .C1(n12360), .C2(n14183), .A(
        n2514), .ZN(n2507) );
  OAI22_X1 U1467 ( .A1(n13932), .A2(n12354), .B1(n13774), .B2(n12348), .ZN(
        n2514) );
  AOI221_X1 U1468 ( .B1(n12462), .B2(n11738), .C1(n12456), .C2(n11558), .A(
        n2506), .ZN(n2499) );
  OAI22_X1 U1469 ( .A1(n13631), .A2(n12450), .B1(n13567), .B2(n12444), .ZN(
        n2506) );
  AOI221_X1 U1470 ( .B1(n12366), .B2(n14011), .C1(n12360), .C2(n14182), .A(
        n2495), .ZN(n2488) );
  OAI22_X1 U1471 ( .A1(n13931), .A2(n12354), .B1(n13773), .B2(n12348), .ZN(
        n2495) );
  AOI221_X1 U1472 ( .B1(n12462), .B2(n11739), .C1(n12456), .C2(n11559), .A(
        n2487), .ZN(n2480) );
  OAI22_X1 U1473 ( .A1(n13630), .A2(n12450), .B1(n13566), .B2(n12444), .ZN(
        n2487) );
  AOI221_X1 U1474 ( .B1(n12366), .B2(n14010), .C1(n12360), .C2(n14181), .A(
        n2476), .ZN(n2469) );
  OAI22_X1 U1475 ( .A1(n13930), .A2(n12354), .B1(n13772), .B2(n12348), .ZN(
        n2476) );
  AOI221_X1 U1476 ( .B1(n12462), .B2(n11740), .C1(n12456), .C2(n11560), .A(
        n2468), .ZN(n2461) );
  OAI22_X1 U1477 ( .A1(n13629), .A2(n12450), .B1(n13565), .B2(n12444), .ZN(
        n2468) );
  AOI221_X1 U1478 ( .B1(n12366), .B2(n14009), .C1(n12360), .C2(n14180), .A(
        n2457), .ZN(n2450) );
  OAI22_X1 U1479 ( .A1(n13929), .A2(n12354), .B1(n13771), .B2(n12348), .ZN(
        n2457) );
  AOI221_X1 U1480 ( .B1(n12462), .B2(n11741), .C1(n12456), .C2(n11561), .A(
        n2449), .ZN(n2442) );
  OAI22_X1 U1481 ( .A1(n13628), .A2(n12450), .B1(n13564), .B2(n12444), .ZN(
        n2449) );
  AOI221_X1 U1482 ( .B1(n12366), .B2(n14008), .C1(n12360), .C2(n14179), .A(
        n2438), .ZN(n2431) );
  OAI22_X1 U1483 ( .A1(n14106), .A2(n12354), .B1(n13770), .B2(n12348), .ZN(
        n2438) );
  AOI221_X1 U1484 ( .B1(n12462), .B2(n11742), .C1(n12456), .C2(n11562), .A(
        n2430), .ZN(n2423) );
  OAI22_X1 U1485 ( .A1(n13627), .A2(n12450), .B1(n13563), .B2(n12444), .ZN(
        n2430) );
  AOI221_X1 U1486 ( .B1(n12366), .B2(n14007), .C1(n12360), .C2(n14178), .A(
        n2419), .ZN(n2412) );
  OAI22_X1 U1487 ( .A1(n14105), .A2(n12354), .B1(n13769), .B2(n12348), .ZN(
        n2419) );
  AOI221_X1 U1488 ( .B1(n12462), .B2(n11743), .C1(n12456), .C2(n11563), .A(
        n2411), .ZN(n2404) );
  OAI22_X1 U1489 ( .A1(n13626), .A2(n12450), .B1(n13562), .B2(n12444), .ZN(
        n2411) );
  AOI221_X1 U1490 ( .B1(n12366), .B2(n14006), .C1(n12360), .C2(n14177), .A(
        n2400), .ZN(n2393) );
  OAI22_X1 U1491 ( .A1(n14104), .A2(n12354), .B1(n13768), .B2(n12348), .ZN(
        n2400) );
  AOI221_X1 U1492 ( .B1(n12462), .B2(n11744), .C1(n12456), .C2(n11564), .A(
        n2392), .ZN(n2385) );
  OAI22_X1 U1493 ( .A1(n13625), .A2(n12450), .B1(n13561), .B2(n12444), .ZN(
        n2392) );
  AOI221_X1 U1494 ( .B1(n12366), .B2(n14005), .C1(n12360), .C2(n14176), .A(
        n2381), .ZN(n2374) );
  OAI22_X1 U1495 ( .A1(n14103), .A2(n12354), .B1(n13767), .B2(n12348), .ZN(
        n2381) );
  AOI221_X1 U1496 ( .B1(n12462), .B2(n11745), .C1(n12456), .C2(n11565), .A(
        n2373), .ZN(n2366) );
  OAI22_X1 U1497 ( .A1(n13624), .A2(n12450), .B1(n13560), .B2(n12444), .ZN(
        n2373) );
  AOI221_X1 U1498 ( .B1(n12366), .B2(n14004), .C1(n12360), .C2(n14175), .A(
        n2362), .ZN(n2355) );
  OAI22_X1 U1499 ( .A1(n14102), .A2(n12354), .B1(n13766), .B2(n12348), .ZN(
        n2362) );
  AOI221_X1 U1500 ( .B1(n12462), .B2(n11746), .C1(n12456), .C2(n11566), .A(
        n2354), .ZN(n2347) );
  OAI22_X1 U1501 ( .A1(n13623), .A2(n12450), .B1(n13559), .B2(n12444), .ZN(
        n2354) );
  AOI221_X1 U1502 ( .B1(n12366), .B2(n14003), .C1(n12360), .C2(n14174), .A(
        n2343), .ZN(n2336) );
  OAI22_X1 U1503 ( .A1(n14101), .A2(n12354), .B1(n13765), .B2(n12348), .ZN(
        n2343) );
  AOI221_X1 U1504 ( .B1(n12462), .B2(n11747), .C1(n12456), .C2(n11567), .A(
        n2335), .ZN(n2328) );
  OAI22_X1 U1505 ( .A1(n13622), .A2(n12450), .B1(n13558), .B2(n12444), .ZN(
        n2335) );
  AOI221_X1 U1506 ( .B1(n12366), .B2(n14002), .C1(n12360), .C2(n14173), .A(
        n2324), .ZN(n2317) );
  OAI22_X1 U1507 ( .A1(n14100), .A2(n12354), .B1(n13764), .B2(n12348), .ZN(
        n2324) );
  AOI221_X1 U1508 ( .B1(n12462), .B2(n11748), .C1(n12456), .C2(n11568), .A(
        n2316), .ZN(n2309) );
  OAI22_X1 U1509 ( .A1(n13621), .A2(n12450), .B1(n13557), .B2(n12444), .ZN(
        n2316) );
  AOI221_X1 U1510 ( .B1(n12366), .B2(n14001), .C1(n12360), .C2(n14172), .A(
        n2305), .ZN(n2298) );
  OAI22_X1 U1511 ( .A1(n14099), .A2(n12354), .B1(n13763), .B2(n12348), .ZN(
        n2305) );
  AOI221_X1 U1512 ( .B1(n12462), .B2(n11749), .C1(n12456), .C2(n11569), .A(
        n2297), .ZN(n2290) );
  OAI22_X1 U1513 ( .A1(n13620), .A2(n12450), .B1(n13556), .B2(n12444), .ZN(
        n2297) );
  AOI221_X1 U1514 ( .B1(n12367), .B2(n14000), .C1(n12361), .C2(n14171), .A(
        n2286), .ZN(n2279) );
  OAI22_X1 U1515 ( .A1(n14098), .A2(n12355), .B1(n13762), .B2(n12349), .ZN(
        n2286) );
  AOI221_X1 U1516 ( .B1(n12463), .B2(n11750), .C1(n12457), .C2(n11570), .A(
        n2278), .ZN(n2271) );
  OAI22_X1 U1517 ( .A1(n13619), .A2(n12451), .B1(n13555), .B2(n12445), .ZN(
        n2278) );
  AOI221_X1 U1518 ( .B1(n12367), .B2(n13999), .C1(n12361), .C2(n14170), .A(
        n2267), .ZN(n2260) );
  OAI22_X1 U1519 ( .A1(n14097), .A2(n12355), .B1(n13761), .B2(n12349), .ZN(
        n2267) );
  AOI221_X1 U1520 ( .B1(n12463), .B2(n11751), .C1(n12457), .C2(n11571), .A(
        n2259), .ZN(n2252) );
  OAI22_X1 U1521 ( .A1(n13618), .A2(n12451), .B1(n13554), .B2(n12445), .ZN(
        n2259) );
  AOI221_X1 U1522 ( .B1(n12367), .B2(n13998), .C1(n12361), .C2(n14169), .A(
        n2248), .ZN(n2241) );
  OAI22_X1 U1523 ( .A1(n14096), .A2(n12355), .B1(n13760), .B2(n12349), .ZN(
        n2248) );
  AOI221_X1 U1524 ( .B1(n12463), .B2(n11752), .C1(n12457), .C2(n11572), .A(
        n2240), .ZN(n2233) );
  OAI22_X1 U1525 ( .A1(n13617), .A2(n12451), .B1(n13553), .B2(n12445), .ZN(
        n2240) );
  AOI221_X1 U1526 ( .B1(n12367), .B2(n13997), .C1(n12361), .C2(n14168), .A(
        n2229), .ZN(n2222) );
  OAI22_X1 U1527 ( .A1(n14095), .A2(n12355), .B1(n13759), .B2(n12349), .ZN(
        n2229) );
  AOI221_X1 U1528 ( .B1(n12463), .B2(n11753), .C1(n12457), .C2(n11573), .A(
        n2221), .ZN(n2214) );
  OAI22_X1 U1529 ( .A1(n13616), .A2(n12451), .B1(n13552), .B2(n12445), .ZN(
        n2221) );
  AOI221_X1 U1530 ( .B1(n12367), .B2(n13996), .C1(n12361), .C2(n14167), .A(
        n2210), .ZN(n2203) );
  OAI22_X1 U1531 ( .A1(n14094), .A2(n12355), .B1(n13758), .B2(n12349), .ZN(
        n2210) );
  AOI221_X1 U1532 ( .B1(n12463), .B2(n11754), .C1(n12457), .C2(n11574), .A(
        n2202), .ZN(n2195) );
  OAI22_X1 U1533 ( .A1(n13615), .A2(n12451), .B1(n13551), .B2(n12445), .ZN(
        n2202) );
  AOI221_X1 U1534 ( .B1(n12367), .B2(n13995), .C1(n12361), .C2(n14166), .A(
        n2191), .ZN(n2184) );
  OAI22_X1 U1535 ( .A1(n14093), .A2(n12355), .B1(n13757), .B2(n12349), .ZN(
        n2191) );
  AOI221_X1 U1536 ( .B1(n12463), .B2(n11755), .C1(n12457), .C2(n11575), .A(
        n2183), .ZN(n2176) );
  OAI22_X1 U1537 ( .A1(n13614), .A2(n12451), .B1(n13550), .B2(n12445), .ZN(
        n2183) );
  AOI221_X1 U1538 ( .B1(n12367), .B2(n13994), .C1(n12361), .C2(n14165), .A(
        n2172), .ZN(n2165) );
  OAI22_X1 U1539 ( .A1(n14092), .A2(n12355), .B1(n13756), .B2(n12349), .ZN(
        n2172) );
  AOI221_X1 U1540 ( .B1(n12463), .B2(n11756), .C1(n12457), .C2(n11576), .A(
        n2164), .ZN(n2157) );
  OAI22_X1 U1541 ( .A1(n13613), .A2(n12451), .B1(n13549), .B2(n12445), .ZN(
        n2164) );
  AOI221_X1 U1542 ( .B1(n12367), .B2(n13993), .C1(n12361), .C2(n14164), .A(
        n2153), .ZN(n2146) );
  OAI22_X1 U1543 ( .A1(n14091), .A2(n12355), .B1(n13755), .B2(n12349), .ZN(
        n2153) );
  AOI221_X1 U1544 ( .B1(n12463), .B2(n11757), .C1(n12457), .C2(n11577), .A(
        n2145), .ZN(n2138) );
  OAI22_X1 U1545 ( .A1(n13612), .A2(n12451), .B1(n13548), .B2(n12445), .ZN(
        n2145) );
  AOI221_X1 U1546 ( .B1(n12367), .B2(n13992), .C1(n12361), .C2(n14163), .A(
        n2134), .ZN(n2127) );
  OAI22_X1 U1547 ( .A1(n14090), .A2(n12355), .B1(n13754), .B2(n12349), .ZN(
        n2134) );
  AOI221_X1 U1548 ( .B1(n12463), .B2(n11758), .C1(n12457), .C2(n11578), .A(
        n2126), .ZN(n2119) );
  OAI22_X1 U1549 ( .A1(n13611), .A2(n12451), .B1(n13547), .B2(n12445), .ZN(
        n2126) );
  AOI221_X1 U1550 ( .B1(n12367), .B2(n13991), .C1(n12361), .C2(n14162), .A(
        n2115), .ZN(n2108) );
  OAI22_X1 U1551 ( .A1(n14089), .A2(n12355), .B1(n13753), .B2(n12349), .ZN(
        n2115) );
  AOI221_X1 U1552 ( .B1(n12463), .B2(n11759), .C1(n12457), .C2(n11579), .A(
        n2107), .ZN(n2100) );
  OAI22_X1 U1553 ( .A1(n13610), .A2(n12451), .B1(n13546), .B2(n12445), .ZN(
        n2107) );
  AOI221_X1 U1554 ( .B1(n12367), .B2(n13990), .C1(n12361), .C2(n14161), .A(
        n2096), .ZN(n2089) );
  OAI22_X1 U1555 ( .A1(n14088), .A2(n12355), .B1(n13752), .B2(n12349), .ZN(
        n2096) );
  AOI221_X1 U1556 ( .B1(n12463), .B2(n11760), .C1(n12457), .C2(n11580), .A(
        n2088), .ZN(n2081) );
  OAI22_X1 U1557 ( .A1(n13609), .A2(n12451), .B1(n13545), .B2(n12445), .ZN(
        n2088) );
  AOI221_X1 U1558 ( .B1(n12367), .B2(n13989), .C1(n12361), .C2(n14160), .A(
        n2077), .ZN(n2070) );
  OAI22_X1 U1559 ( .A1(n14087), .A2(n12355), .B1(n13751), .B2(n12349), .ZN(
        n2077) );
  AOI221_X1 U1560 ( .B1(n12463), .B2(n11761), .C1(n12457), .C2(n11581), .A(
        n2069), .ZN(n2062) );
  OAI22_X1 U1561 ( .A1(n13608), .A2(n12451), .B1(n13544), .B2(n12445), .ZN(
        n2069) );
  AOI221_X1 U1562 ( .B1(n12368), .B2(n13827), .C1(n12362), .C2(n14159), .A(
        n2058), .ZN(n2051) );
  OAI22_X1 U1563 ( .A1(n14086), .A2(n12356), .B1(n13750), .B2(n12350), .ZN(
        n2058) );
  AOI221_X1 U1564 ( .B1(n12464), .B2(n13864), .C1(n12458), .C2(n13868), .A(
        n2050), .ZN(n2043) );
  OAI22_X1 U1565 ( .A1(n13607), .A2(n12452), .B1(n13543), .B2(n12446), .ZN(
        n2050) );
  AOI221_X1 U1566 ( .B1(n12368), .B2(n13826), .C1(n12362), .C2(n14158), .A(
        n2039), .ZN(n2032) );
  OAI22_X1 U1567 ( .A1(n14085), .A2(n12356), .B1(n13749), .B2(n12350), .ZN(
        n2039) );
  AOI221_X1 U1568 ( .B1(n12464), .B2(n13863), .C1(n12458), .C2(n13867), .A(
        n2031), .ZN(n2024) );
  OAI22_X1 U1569 ( .A1(n13606), .A2(n12452), .B1(n13542), .B2(n12446), .ZN(
        n2031) );
  AOI221_X1 U1570 ( .B1(n12368), .B2(n13825), .C1(n12362), .C2(n14157), .A(
        n2020), .ZN(n2013) );
  OAI22_X1 U1571 ( .A1(n14084), .A2(n12356), .B1(n13748), .B2(n12350), .ZN(
        n2020) );
  AOI221_X1 U1572 ( .B1(n12464), .B2(n13862), .C1(n12458), .C2(n13866), .A(
        n2012), .ZN(n2005) );
  OAI22_X1 U1573 ( .A1(n13605), .A2(n12452), .B1(n13541), .B2(n12446), .ZN(
        n2012) );
  AOI221_X1 U1574 ( .B1(n12368), .B2(n13824), .C1(n12362), .C2(n14156), .A(
        n1999), .ZN(n1978) );
  OAI22_X1 U1575 ( .A1(n14083), .A2(n12356), .B1(n13747), .B2(n12350), .ZN(
        n1999) );
  AOI221_X1 U1576 ( .B1(n12464), .B2(n13861), .C1(n12458), .C2(n13865), .A(
        n1975), .ZN(n1954) );
  OAI22_X1 U1577 ( .A1(n13604), .A2(n12452), .B1(n13540), .B2(n12446), .ZN(
        n1975) );
  NOR3_X1 U1578 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n14461), .ZN(n3204) );
  AOI221_X1 U1579 ( .B1(n12387), .B2(n14079), .C1(n12381), .C2(n14126), .A(
        n3140), .ZN(n3135) );
  OAI22_X1 U1580 ( .A1(n13743), .A2(n12375), .B1(n13727), .B2(n12369), .ZN(
        n3140) );
  AOI221_X1 U1581 ( .B1(n12387), .B2(n14080), .C1(n12381), .C2(n14127), .A(
        n3121), .ZN(n3116) );
  OAI22_X1 U1582 ( .A1(n13892), .A2(n12375), .B1(n13726), .B2(n12369), .ZN(
        n3121) );
  AOI221_X1 U1583 ( .B1(n12387), .B2(n14076), .C1(n12381), .C2(n14123), .A(
        n3064), .ZN(n3059) );
  OAI22_X1 U1584 ( .A1(n13889), .A2(n12375), .B1(n13723), .B2(n12369), .ZN(
        n3064) );
  AOI221_X1 U1585 ( .B1(n12387), .B2(n14075), .C1(n12381), .C2(n14122), .A(
        n3045), .ZN(n3040) );
  OAI22_X1 U1586 ( .A1(n13888), .A2(n12375), .B1(n13722), .B2(n12369), .ZN(
        n3045) );
  AOI221_X1 U1587 ( .B1(n12387), .B2(n14074), .C1(n12381), .C2(n14121), .A(
        n3026), .ZN(n3021) );
  OAI22_X1 U1588 ( .A1(n13887), .A2(n12375), .B1(n13721), .B2(n12369), .ZN(
        n3026) );
  AOI221_X1 U1589 ( .B1(n12387), .B2(n14073), .C1(n12381), .C2(n14120), .A(
        n3007), .ZN(n3002) );
  OAI22_X1 U1590 ( .A1(n13886), .A2(n12375), .B1(n13720), .B2(n12369), .ZN(
        n3007) );
  AOI221_X1 U1591 ( .B1(n12387), .B2(n14072), .C1(n12381), .C2(n14119), .A(
        n2988), .ZN(n2983) );
  OAI22_X1 U1592 ( .A1(n13885), .A2(n12375), .B1(n13719), .B2(n12369), .ZN(
        n2988) );
  AOI221_X1 U1593 ( .B1(n12388), .B2(n14071), .C1(n12382), .C2(n14118), .A(
        n2969), .ZN(n2964) );
  OAI22_X1 U1594 ( .A1(n13884), .A2(n12376), .B1(n13718), .B2(n12370), .ZN(
        n2969) );
  AOI221_X1 U1595 ( .B1(n12388), .B2(n14070), .C1(n12382), .C2(n14117), .A(
        n2950), .ZN(n2945) );
  OAI22_X1 U1596 ( .A1(n13883), .A2(n12376), .B1(n13717), .B2(n12370), .ZN(
        n2950) );
  AOI221_X1 U1597 ( .B1(n12388), .B2(n14069), .C1(n12382), .C2(n14116), .A(
        n2931), .ZN(n2926) );
  OAI22_X1 U1598 ( .A1(n13882), .A2(n12376), .B1(n13716), .B2(n12370), .ZN(
        n2931) );
  AOI221_X1 U1599 ( .B1(n12388), .B2(n14068), .C1(n12382), .C2(n14115), .A(
        n2912), .ZN(n2907) );
  OAI22_X1 U1600 ( .A1(n13881), .A2(n12376), .B1(n13715), .B2(n12370), .ZN(
        n2912) );
  AOI221_X1 U1601 ( .B1(n12388), .B2(n14067), .C1(n12382), .C2(n14114), .A(
        n2893), .ZN(n2888) );
  OAI22_X1 U1602 ( .A1(n13880), .A2(n12376), .B1(n13714), .B2(n12370), .ZN(
        n2893) );
  AOI221_X1 U1603 ( .B1(n12388), .B2(n14066), .C1(n12382), .C2(n14113), .A(
        n2874), .ZN(n2869) );
  OAI22_X1 U1604 ( .A1(n13879), .A2(n12376), .B1(n13713), .B2(n12370), .ZN(
        n2874) );
  AOI221_X1 U1605 ( .B1(n12388), .B2(n14065), .C1(n12382), .C2(n14112), .A(
        n2855), .ZN(n2850) );
  OAI22_X1 U1606 ( .A1(n13878), .A2(n12376), .B1(n13712), .B2(n12370), .ZN(
        n2855) );
  AOI221_X1 U1607 ( .B1(n12388), .B2(n14064), .C1(n12382), .C2(n14111), .A(
        n2836), .ZN(n2831) );
  OAI22_X1 U1608 ( .A1(n13877), .A2(n12376), .B1(n13711), .B2(n12370), .ZN(
        n2836) );
  AOI221_X1 U1609 ( .B1(n12388), .B2(n14063), .C1(n12382), .C2(n14110), .A(
        n2817), .ZN(n2812) );
  OAI22_X1 U1610 ( .A1(n13876), .A2(n12376), .B1(n13710), .B2(n12370), .ZN(
        n2817) );
  AOI221_X1 U1611 ( .B1(n12388), .B2(n14062), .C1(n12382), .C2(n14109), .A(
        n2798), .ZN(n2793) );
  OAI22_X1 U1612 ( .A1(n13875), .A2(n12376), .B1(n13709), .B2(n12370), .ZN(
        n2798) );
  AOI221_X1 U1613 ( .B1(n12388), .B2(n14061), .C1(n12382), .C2(n14108), .A(
        n2779), .ZN(n2774) );
  OAI22_X1 U1614 ( .A1(n13874), .A2(n12376), .B1(n13708), .B2(n12370), .ZN(
        n2779) );
  AOI221_X1 U1615 ( .B1(n12388), .B2(n14060), .C1(n12382), .C2(n14107), .A(
        n2760), .ZN(n2755) );
  OAI22_X1 U1616 ( .A1(n13873), .A2(n12376), .B1(n13707), .B2(n12370), .ZN(
        n2760) );
  AOI221_X1 U1617 ( .B1(n12389), .B2(n13928), .C1(n12383), .C2(n13988), .A(
        n2741), .ZN(n2736) );
  OAI22_X1 U1618 ( .A1(n13872), .A2(n12377), .B1(n13706), .B2(n12371), .ZN(
        n2741) );
  AOI221_X1 U1619 ( .B1(n12389), .B2(n13927), .C1(n12383), .C2(n13987), .A(
        n2722), .ZN(n2717) );
  OAI22_X1 U1620 ( .A1(n13871), .A2(n12377), .B1(n13705), .B2(n12371), .ZN(
        n2722) );
  AOI221_X1 U1621 ( .B1(n12389), .B2(n13926), .C1(n12383), .C2(n13986), .A(
        n2703), .ZN(n2698) );
  OAI22_X1 U1622 ( .A1(n13870), .A2(n12377), .B1(n13704), .B2(n12371), .ZN(
        n2703) );
  AOI221_X1 U1623 ( .B1(n12389), .B2(n13925), .C1(n12383), .C2(n13985), .A(
        n2684), .ZN(n2679) );
  OAI22_X1 U1624 ( .A1(n13869), .A2(n12377), .B1(n13703), .B2(n12371), .ZN(
        n2684) );
  AOI221_X1 U1625 ( .B1(n12389), .B2(n13924), .C1(n12383), .C2(n13984), .A(
        n2665), .ZN(n2660) );
  OAI22_X1 U1626 ( .A1(n14059), .A2(n12377), .B1(n13702), .B2(n12371), .ZN(
        n2665) );
  AOI221_X1 U1627 ( .B1(n12389), .B2(n13923), .C1(n12383), .C2(n13983), .A(
        n2646), .ZN(n2641) );
  OAI22_X1 U1628 ( .A1(n14058), .A2(n12377), .B1(n13701), .B2(n12371), .ZN(
        n2646) );
  AOI221_X1 U1629 ( .B1(n12389), .B2(n13922), .C1(n12383), .C2(n13982), .A(
        n2627), .ZN(n2622) );
  OAI22_X1 U1630 ( .A1(n14057), .A2(n12377), .B1(n13700), .B2(n12371), .ZN(
        n2627) );
  AOI221_X1 U1631 ( .B1(n12389), .B2(n13921), .C1(n12383), .C2(n13981), .A(
        n2608), .ZN(n2603) );
  OAI22_X1 U1632 ( .A1(n14056), .A2(n12377), .B1(n13699), .B2(n12371), .ZN(
        n2608) );
  AOI221_X1 U1633 ( .B1(n12389), .B2(n13920), .C1(n12383), .C2(n13980), .A(
        n2589), .ZN(n2584) );
  OAI22_X1 U1634 ( .A1(n14055), .A2(n12377), .B1(n13698), .B2(n12371), .ZN(
        n2589) );
  AOI221_X1 U1635 ( .B1(n12389), .B2(n13919), .C1(n12383), .C2(n13979), .A(
        n2570), .ZN(n2565) );
  OAI22_X1 U1636 ( .A1(n14054), .A2(n12377), .B1(n13697), .B2(n12371), .ZN(
        n2570) );
  AOI221_X1 U1637 ( .B1(n12389), .B2(n13918), .C1(n12383), .C2(n13978), .A(
        n2551), .ZN(n2546) );
  OAI22_X1 U1638 ( .A1(n14053), .A2(n12377), .B1(n13696), .B2(n12371), .ZN(
        n2551) );
  AOI221_X1 U1639 ( .B1(n12389), .B2(n13917), .C1(n12383), .C2(n13977), .A(
        n2532), .ZN(n2527) );
  OAI22_X1 U1640 ( .A1(n14052), .A2(n12377), .B1(n13695), .B2(n12371), .ZN(
        n2532) );
  AOI221_X1 U1641 ( .B1(n12390), .B2(n13916), .C1(n12384), .C2(n13976), .A(
        n2513), .ZN(n2508) );
  OAI22_X1 U1642 ( .A1(n14051), .A2(n12378), .B1(n13694), .B2(n12372), .ZN(
        n2513) );
  AOI221_X1 U1643 ( .B1(n12390), .B2(n13915), .C1(n12384), .C2(n13975), .A(
        n2494), .ZN(n2489) );
  OAI22_X1 U1644 ( .A1(n14050), .A2(n12378), .B1(n13693), .B2(n12372), .ZN(
        n2494) );
  AOI221_X1 U1645 ( .B1(n12390), .B2(n13914), .C1(n12384), .C2(n13974), .A(
        n2475), .ZN(n2470) );
  OAI22_X1 U1646 ( .A1(n14049), .A2(n12378), .B1(n13692), .B2(n12372), .ZN(
        n2475) );
  AOI221_X1 U1647 ( .B1(n12390), .B2(n13913), .C1(n12384), .C2(n13973), .A(
        n2456), .ZN(n2451) );
  OAI22_X1 U1648 ( .A1(n14048), .A2(n12378), .B1(n13691), .B2(n12372), .ZN(
        n2456) );
  AOI221_X1 U1649 ( .B1(n12390), .B2(n13912), .C1(n12384), .C2(n13972), .A(
        n2437), .ZN(n2432) );
  OAI22_X1 U1650 ( .A1(n14047), .A2(n12378), .B1(n13690), .B2(n12372), .ZN(
        n2437) );
  AOI221_X1 U1651 ( .B1(n12390), .B2(n13911), .C1(n12384), .C2(n13971), .A(
        n2418), .ZN(n2413) );
  OAI22_X1 U1652 ( .A1(n14046), .A2(n12378), .B1(n13689), .B2(n12372), .ZN(
        n2418) );
  AOI221_X1 U1653 ( .B1(n12390), .B2(n13910), .C1(n12384), .C2(n13970), .A(
        n2399), .ZN(n2394) );
  OAI22_X1 U1654 ( .A1(n14045), .A2(n12378), .B1(n13688), .B2(n12372), .ZN(
        n2399) );
  AOI221_X1 U1655 ( .B1(n12390), .B2(n13909), .C1(n12384), .C2(n13969), .A(
        n2380), .ZN(n2375) );
  OAI22_X1 U1656 ( .A1(n14044), .A2(n12378), .B1(n13687), .B2(n12372), .ZN(
        n2380) );
  AOI221_X1 U1657 ( .B1(n12390), .B2(n13908), .C1(n12384), .C2(n13968), .A(
        n2361), .ZN(n2356) );
  OAI22_X1 U1658 ( .A1(n14043), .A2(n12378), .B1(n13686), .B2(n12372), .ZN(
        n2361) );
  AOI221_X1 U1659 ( .B1(n12390), .B2(n13907), .C1(n12384), .C2(n13967), .A(
        n2342), .ZN(n2337) );
  OAI22_X1 U1660 ( .A1(n14042), .A2(n12378), .B1(n13685), .B2(n12372), .ZN(
        n2342) );
  AOI221_X1 U1661 ( .B1(n12390), .B2(n13906), .C1(n12384), .C2(n13966), .A(
        n2323), .ZN(n2318) );
  OAI22_X1 U1662 ( .A1(n14041), .A2(n12378), .B1(n13684), .B2(n12372), .ZN(
        n2323) );
  AOI221_X1 U1663 ( .B1(n12390), .B2(n13905), .C1(n12384), .C2(n13965), .A(
        n2304), .ZN(n2299) );
  OAI22_X1 U1664 ( .A1(n14040), .A2(n12378), .B1(n13683), .B2(n12372), .ZN(
        n2304) );
  AOI221_X1 U1665 ( .B1(n12391), .B2(n13904), .C1(n12385), .C2(n13964), .A(
        n2285), .ZN(n2280) );
  OAI22_X1 U1666 ( .A1(n14039), .A2(n12379), .B1(n13682), .B2(n12373), .ZN(
        n2285) );
  AOI221_X1 U1667 ( .B1(n12391), .B2(n13903), .C1(n12385), .C2(n13963), .A(
        n2266), .ZN(n2261) );
  OAI22_X1 U1668 ( .A1(n14038), .A2(n12379), .B1(n13681), .B2(n12373), .ZN(
        n2266) );
  AOI221_X1 U1669 ( .B1(n12391), .B2(n13902), .C1(n12385), .C2(n13962), .A(
        n2247), .ZN(n2242) );
  OAI22_X1 U1670 ( .A1(n14037), .A2(n12379), .B1(n13680), .B2(n12373), .ZN(
        n2247) );
  AOI221_X1 U1671 ( .B1(n12391), .B2(n13901), .C1(n12385), .C2(n13961), .A(
        n2228), .ZN(n2223) );
  OAI22_X1 U1672 ( .A1(n14036), .A2(n12379), .B1(n13679), .B2(n12373), .ZN(
        n2228) );
  AOI221_X1 U1673 ( .B1(n12391), .B2(n13900), .C1(n12385), .C2(n13960), .A(
        n2209), .ZN(n2204) );
  OAI22_X1 U1674 ( .A1(n13742), .A2(n12379), .B1(n13678), .B2(n12373), .ZN(
        n2209) );
  AOI221_X1 U1675 ( .B1(n12391), .B2(n13899), .C1(n12385), .C2(n13959), .A(
        n2190), .ZN(n2185) );
  OAI22_X1 U1676 ( .A1(n13741), .A2(n12379), .B1(n13677), .B2(n12373), .ZN(
        n2190) );
  AOI221_X1 U1677 ( .B1(n12391), .B2(n13898), .C1(n12385), .C2(n13958), .A(
        n2171), .ZN(n2166) );
  OAI22_X1 U1678 ( .A1(n13740), .A2(n12379), .B1(n13676), .B2(n12373), .ZN(
        n2171) );
  AOI221_X1 U1679 ( .B1(n12391), .B2(n13897), .C1(n12385), .C2(n13957), .A(
        n2152), .ZN(n2147) );
  OAI22_X1 U1680 ( .A1(n13739), .A2(n12379), .B1(n13675), .B2(n12373), .ZN(
        n2152) );
  AOI221_X1 U1681 ( .B1(n12391), .B2(n13896), .C1(n12385), .C2(n13956), .A(
        n2133), .ZN(n2128) );
  OAI22_X1 U1682 ( .A1(n13738), .A2(n12379), .B1(n13674), .B2(n12373), .ZN(
        n2133) );
  AOI221_X1 U1683 ( .B1(n12391), .B2(n13895), .C1(n12385), .C2(n13955), .A(
        n2114), .ZN(n2109) );
  OAI22_X1 U1684 ( .A1(n13737), .A2(n12379), .B1(n13673), .B2(n12373), .ZN(
        n2114) );
  AOI221_X1 U1685 ( .B1(n12391), .B2(n13894), .C1(n12385), .C2(n13954), .A(
        n2095), .ZN(n2090) );
  OAI22_X1 U1686 ( .A1(n13736), .A2(n12379), .B1(n13672), .B2(n12373), .ZN(
        n2095) );
  OAI22_X1 U1687 ( .A1(n13107), .A2(n13173), .B1(n13093), .B2(n14408), .ZN(
        n6719) );
  OAI22_X1 U1688 ( .A1(n13107), .A2(n13176), .B1(n13094), .B2(n14407), .ZN(
        n6720) );
  OAI22_X1 U1689 ( .A1(n13107), .A2(n13179), .B1(n13091), .B2(n14406), .ZN(
        n6721) );
  OAI22_X1 U1690 ( .A1(n13106), .A2(n13182), .B1(n13093), .B2(n14405), .ZN(
        n6722) );
  OAI22_X1 U1691 ( .A1(n13106), .A2(n13185), .B1(n13094), .B2(n14404), .ZN(
        n6723) );
  OAI22_X1 U1692 ( .A1(n13106), .A2(n13188), .B1(n13090), .B2(n14403), .ZN(
        n6724) );
  OAI22_X1 U1693 ( .A1(n13106), .A2(n13191), .B1(n1914), .B2(n14402), .ZN(
        n6725) );
  OAI22_X1 U1694 ( .A1(n13106), .A2(n13194), .B1(n1914), .B2(n14401), .ZN(
        n6726) );
  OAI22_X1 U1695 ( .A1(n13105), .A2(n13197), .B1(n1914), .B2(n14400), .ZN(
        n6727) );
  OAI22_X1 U1696 ( .A1(n13105), .A2(n13200), .B1(n1914), .B2(n14399), .ZN(
        n6728) );
  OAI22_X1 U1697 ( .A1(n13105), .A2(n13203), .B1(n1914), .B2(n14398), .ZN(
        n6729) );
  OAI22_X1 U1698 ( .A1(n13105), .A2(n13206), .B1(n13091), .B2(n14397), .ZN(
        n6730) );
  OAI22_X1 U1699 ( .A1(n13105), .A2(n13209), .B1(n13091), .B2(n14396), .ZN(
        n6731) );
  OAI22_X1 U1700 ( .A1(n13104), .A2(n13212), .B1(n13091), .B2(n14395), .ZN(
        n6732) );
  OAI22_X1 U1701 ( .A1(n13104), .A2(n13215), .B1(n13091), .B2(n14394), .ZN(
        n6733) );
  OAI22_X1 U1702 ( .A1(n13104), .A2(n13218), .B1(n13091), .B2(n14393), .ZN(
        n6734) );
  OAI22_X1 U1703 ( .A1(n13104), .A2(n13221), .B1(n13091), .B2(n14392), .ZN(
        n6735) );
  OAI22_X1 U1704 ( .A1(n13104), .A2(n13224), .B1(n13091), .B2(n14391), .ZN(
        n6736) );
  OAI22_X1 U1705 ( .A1(n13103), .A2(n13227), .B1(n13091), .B2(n14390), .ZN(
        n6737) );
  OAI22_X1 U1706 ( .A1(n13103), .A2(n13230), .B1(n13091), .B2(n14389), .ZN(
        n6738) );
  OAI22_X1 U1707 ( .A1(n13103), .A2(n13233), .B1(n13091), .B2(n14388), .ZN(
        n6739) );
  OAI22_X1 U1708 ( .A1(n13103), .A2(n13236), .B1(n13091), .B2(n14387), .ZN(
        n6740) );
  OAI22_X1 U1709 ( .A1(n13103), .A2(n13239), .B1(n13091), .B2(n14386), .ZN(
        n6741) );
  OAI22_X1 U1710 ( .A1(n13087), .A2(n13173), .B1(n13073), .B2(n14385), .ZN(
        n6655) );
  OAI22_X1 U1711 ( .A1(n13087), .A2(n13176), .B1(n13074), .B2(n14384), .ZN(
        n6656) );
  OAI22_X1 U1712 ( .A1(n13087), .A2(n13179), .B1(n13071), .B2(n14383), .ZN(
        n6657) );
  OAI22_X1 U1713 ( .A1(n13086), .A2(n13182), .B1(n13073), .B2(n14382), .ZN(
        n6658) );
  OAI22_X1 U1714 ( .A1(n13086), .A2(n13185), .B1(n13074), .B2(n14381), .ZN(
        n6659) );
  OAI22_X1 U1715 ( .A1(n13086), .A2(n13188), .B1(n13070), .B2(n14380), .ZN(
        n6660) );
  OAI22_X1 U1716 ( .A1(n13086), .A2(n13191), .B1(n1916), .B2(n14379), .ZN(
        n6661) );
  OAI22_X1 U1717 ( .A1(n13086), .A2(n13194), .B1(n1916), .B2(n14378), .ZN(
        n6662) );
  OAI22_X1 U1718 ( .A1(n13085), .A2(n13197), .B1(n1916), .B2(n14377), .ZN(
        n6663) );
  OAI22_X1 U1719 ( .A1(n13085), .A2(n13200), .B1(n1916), .B2(n14376), .ZN(
        n6664) );
  OAI22_X1 U1720 ( .A1(n13085), .A2(n13203), .B1(n1916), .B2(n14375), .ZN(
        n6665) );
  OAI22_X1 U1721 ( .A1(n13085), .A2(n13206), .B1(n13071), .B2(n14374), .ZN(
        n6666) );
  OAI22_X1 U1722 ( .A1(n13085), .A2(n13209), .B1(n13071), .B2(n14373), .ZN(
        n6667) );
  OAI22_X1 U1723 ( .A1(n13084), .A2(n13212), .B1(n13071), .B2(n14372), .ZN(
        n6668) );
  OAI22_X1 U1724 ( .A1(n13084), .A2(n13215), .B1(n13071), .B2(n14371), .ZN(
        n6669) );
  OAI22_X1 U1725 ( .A1(n13084), .A2(n13218), .B1(n13071), .B2(n14370), .ZN(
        n6670) );
  OAI22_X1 U1726 ( .A1(n13084), .A2(n13221), .B1(n13071), .B2(n14369), .ZN(
        n6671) );
  OAI22_X1 U1727 ( .A1(n13084), .A2(n13224), .B1(n13071), .B2(n14368), .ZN(
        n6672) );
  OAI22_X1 U1728 ( .A1(n13083), .A2(n13227), .B1(n13071), .B2(n14367), .ZN(
        n6673) );
  OAI22_X1 U1729 ( .A1(n13083), .A2(n13230), .B1(n13071), .B2(n14366), .ZN(
        n6674) );
  OAI22_X1 U1730 ( .A1(n13083), .A2(n13233), .B1(n13071), .B2(n14365), .ZN(
        n6675) );
  OAI22_X1 U1731 ( .A1(n13083), .A2(n13236), .B1(n13071), .B2(n14364), .ZN(
        n6676) );
  OAI22_X1 U1732 ( .A1(n13083), .A2(n13239), .B1(n13071), .B2(n14363), .ZN(
        n6677) );
  OAI22_X1 U1733 ( .A1(n13107), .A2(n13170), .B1(n1914), .B2(n14362), .ZN(
        n6718) );
  OAI22_X1 U1734 ( .A1(n13087), .A2(n13170), .B1(n1916), .B2(n14361), .ZN(
        n6654) );
  OAI22_X1 U1735 ( .A1(n12966), .A2(n13182), .B1(n12951), .B2(n14360), .ZN(
        n6274) );
  OAI22_X1 U1736 ( .A1(n12966), .A2(n13185), .B1(n12951), .B2(n14359), .ZN(
        n6275) );
  OAI22_X1 U1737 ( .A1(n12966), .A2(n13188), .B1(n12951), .B2(n14358), .ZN(
        n6276) );
  OAI22_X1 U1738 ( .A1(n12886), .A2(n13183), .B1(n12871), .B2(n14357), .ZN(
        n6018) );
  OAI22_X1 U1739 ( .A1(n12886), .A2(n13186), .B1(n12871), .B2(n14356), .ZN(
        n6019) );
  OAI22_X1 U1740 ( .A1(n12886), .A2(n13189), .B1(n12871), .B2(n14355), .ZN(
        n6020) );
  OAI22_X1 U1741 ( .A1(n12886), .A2(n13192), .B1(n12871), .B2(n14354), .ZN(
        n6021) );
  OAI22_X1 U1742 ( .A1(n12886), .A2(n13195), .B1(n12871), .B2(n14353), .ZN(
        n6022) );
  OAI22_X1 U1743 ( .A1(n12885), .A2(n13198), .B1(n12871), .B2(n14352), .ZN(
        n6023) );
  OAI22_X1 U1744 ( .A1(n12885), .A2(n13201), .B1(n12871), .B2(n14351), .ZN(
        n6024) );
  OAI22_X1 U1745 ( .A1(n12885), .A2(n13204), .B1(n12871), .B2(n14350), .ZN(
        n6025) );
  OAI22_X1 U1746 ( .A1(n12885), .A2(n13207), .B1(n12873), .B2(n14349), .ZN(
        n6026) );
  OAI22_X1 U1747 ( .A1(n12885), .A2(n13210), .B1(n12874), .B2(n14348), .ZN(
        n6027) );
  OAI22_X1 U1748 ( .A1(n12884), .A2(n13213), .B1(n12871), .B2(n14347), .ZN(
        n6028) );
  OAI22_X1 U1749 ( .A1(n12884), .A2(n13216), .B1(n12873), .B2(n14346), .ZN(
        n6029) );
  OAI22_X1 U1750 ( .A1(n12884), .A2(n13222), .B1(n12874), .B2(n14345), .ZN(
        n6031) );
  OAI22_X1 U1751 ( .A1(n12884), .A2(n13225), .B1(n12870), .B2(n14344), .ZN(
        n6032) );
  OAI22_X1 U1752 ( .A1(n12883), .A2(n13228), .B1(n1931), .B2(n14343), .ZN(
        n6033) );
  OAI22_X1 U1753 ( .A1(n12883), .A2(n13231), .B1(n1931), .B2(n14342), .ZN(
        n6034) );
  OAI22_X1 U1754 ( .A1(n12883), .A2(n13234), .B1(n1931), .B2(n14341), .ZN(
        n6035) );
  OAI22_X1 U1755 ( .A1(n12966), .A2(n13191), .B1(n12951), .B2(n14340), .ZN(
        n6277) );
  OAI22_X1 U1756 ( .A1(n12966), .A2(n13194), .B1(n12951), .B2(n14339), .ZN(
        n6278) );
  OAI22_X1 U1757 ( .A1(n12965), .A2(n13197), .B1(n12951), .B2(n14338), .ZN(
        n6279) );
  OAI22_X1 U1758 ( .A1(n12965), .A2(n13200), .B1(n12951), .B2(n14337), .ZN(
        n6280) );
  OAI22_X1 U1759 ( .A1(n12965), .A2(n13203), .B1(n12951), .B2(n14336), .ZN(
        n6281) );
  OAI22_X1 U1760 ( .A1(n12965), .A2(n13206), .B1(n12953), .B2(n14335), .ZN(
        n6282) );
  OAI22_X1 U1761 ( .A1(n12965), .A2(n13209), .B1(n12954), .B2(n14334), .ZN(
        n6283) );
  OAI22_X1 U1762 ( .A1(n12964), .A2(n13212), .B1(n12951), .B2(n14333), .ZN(
        n6284) );
  OAI22_X1 U1763 ( .A1(n12964), .A2(n13215), .B1(n12953), .B2(n14332), .ZN(
        n6285) );
  OAI22_X1 U1764 ( .A1(n12964), .A2(n13221), .B1(n12954), .B2(n14331), .ZN(
        n6287) );
  OAI22_X1 U1765 ( .A1(n12964), .A2(n13224), .B1(n12950), .B2(n14330), .ZN(
        n6288) );
  OAI22_X1 U1766 ( .A1(n12963), .A2(n13227), .B1(n1927), .B2(n14329), .ZN(
        n6289) );
  OAI22_X1 U1767 ( .A1(n13376), .A2(n13173), .B1(n13362), .B2(n14328), .ZN(
        n6975) );
  OAI22_X1 U1768 ( .A1(n13376), .A2(n13176), .B1(n13363), .B2(n14327), .ZN(
        n6976) );
  OAI22_X1 U1769 ( .A1(n13376), .A2(n13179), .B1(n13360), .B2(n14326), .ZN(
        n6977) );
  OAI22_X1 U1770 ( .A1(n13375), .A2(n13182), .B1(n13362), .B2(n14325), .ZN(
        n6978) );
  OAI22_X1 U1771 ( .A1(n13375), .A2(n13185), .B1(n13363), .B2(n14324), .ZN(
        n6979) );
  OAI22_X1 U1772 ( .A1(n13375), .A2(n13194), .B1(n13359), .B2(n14323), .ZN(
        n6982) );
  OAI22_X1 U1773 ( .A1(n13375), .A2(n13188), .B1(n1842), .B2(n14311), .ZN(
        n6980) );
  OAI22_X1 U1774 ( .A1(n13375), .A2(n13191), .B1(n1842), .B2(n14310), .ZN(
        n6981) );
  OAI22_X1 U1775 ( .A1(n13374), .A2(n13197), .B1(n1842), .B2(n14309), .ZN(
        n6983) );
  OAI22_X1 U1776 ( .A1(n13374), .A2(n13200), .B1(n1842), .B2(n14308), .ZN(
        n6984) );
  OAI22_X1 U1777 ( .A1(n13374), .A2(n13203), .B1(n1842), .B2(n14307), .ZN(
        n6985) );
  OAI22_X1 U1778 ( .A1(n13374), .A2(n13206), .B1(n13360), .B2(n14306), .ZN(
        n6986) );
  OAI22_X1 U1779 ( .A1(n13374), .A2(n13209), .B1(n13360), .B2(n14305), .ZN(
        n6987) );
  OAI22_X1 U1780 ( .A1(n13373), .A2(n13212), .B1(n13360), .B2(n14304), .ZN(
        n6988) );
  OAI22_X1 U1781 ( .A1(n13373), .A2(n13215), .B1(n13360), .B2(n14303), .ZN(
        n6989) );
  OAI22_X1 U1782 ( .A1(n13373), .A2(n13218), .B1(n13360), .B2(n14302), .ZN(
        n6990) );
  OAI22_X1 U1783 ( .A1(n13373), .A2(n13221), .B1(n13360), .B2(n14301), .ZN(
        n6991) );
  OAI22_X1 U1784 ( .A1(n13373), .A2(n13224), .B1(n13360), .B2(n14300), .ZN(
        n6992) );
  OAI22_X1 U1785 ( .A1(n13372), .A2(n13227), .B1(n13360), .B2(n14299), .ZN(
        n6993) );
  OAI22_X1 U1786 ( .A1(n13372), .A2(n13230), .B1(n13360), .B2(n14298), .ZN(
        n6994) );
  OAI22_X1 U1787 ( .A1(n13372), .A2(n13233), .B1(n13360), .B2(n14297), .ZN(
        n6995) );
  OAI22_X1 U1788 ( .A1(n13372), .A2(n13236), .B1(n13360), .B2(n14296), .ZN(
        n6996) );
  OAI22_X1 U1789 ( .A1(n13372), .A2(n13239), .B1(n13360), .B2(n14295), .ZN(
        n6997) );
  OAI22_X1 U1790 ( .A1(n13376), .A2(n13170), .B1(n1842), .B2(n14216), .ZN(
        n6974) );
  OAI22_X1 U1791 ( .A1(n12611), .A2(n13187), .B1(n12597), .B2(n14035), .ZN(
        n5123) );
  OAI22_X1 U1792 ( .A1(n12611), .A2(n13190), .B1(n12598), .B2(n14034), .ZN(
        n5124) );
  OAI22_X1 U1793 ( .A1(n12611), .A2(n13193), .B1(n12599), .B2(n14033), .ZN(
        n5125) );
  OAI22_X1 U1794 ( .A1(n12611), .A2(n13196), .B1(n12597), .B2(n14032), .ZN(
        n5126) );
  OAI22_X1 U1795 ( .A1(n12610), .A2(n13199), .B1(n12598), .B2(n14031), .ZN(
        n5127) );
  OAI22_X1 U1796 ( .A1(n12610), .A2(n13202), .B1(n12596), .B2(n14030), .ZN(
        n5128) );
  OAI22_X1 U1797 ( .A1(n12610), .A2(n13205), .B1(n1947), .B2(n14029), .ZN(
        n5129) );
  OAI22_X1 U1798 ( .A1(n12610), .A2(n13208), .B1(n12599), .B2(n14028), .ZN(
        n5130) );
  OAI22_X1 U1799 ( .A1(n12610), .A2(n13211), .B1(n12596), .B2(n14027), .ZN(
        n5131) );
  OAI22_X1 U1800 ( .A1(n12609), .A2(n13214), .B1(n12596), .B2(n14026), .ZN(
        n5132) );
  OAI22_X1 U1801 ( .A1(n12609), .A2(n13217), .B1(n1947), .B2(n14025), .ZN(
        n5133) );
  OAI22_X1 U1802 ( .A1(n12609), .A2(n13220), .B1(n1947), .B2(n13952), .ZN(
        n5134) );
  OAI22_X1 U1803 ( .A1(n12609), .A2(n13223), .B1(n1947), .B2(n13951), .ZN(
        n5135) );
  OAI22_X1 U1804 ( .A1(n12609), .A2(n13226), .B1(n1947), .B2(n13950), .ZN(
        n5136) );
  OAI22_X1 U1805 ( .A1(n12608), .A2(n13229), .B1(n1947), .B2(n13949), .ZN(
        n5137) );
  OAI22_X1 U1806 ( .A1(n12608), .A2(n13232), .B1(n12596), .B2(n13948), .ZN(
        n5138) );
  OAI22_X1 U1807 ( .A1(n12608), .A2(n13235), .B1(n12596), .B2(n13947), .ZN(
        n5139) );
  OAI22_X1 U1808 ( .A1(n12608), .A2(n13238), .B1(n12596), .B2(n13946), .ZN(
        n5140) );
  OAI22_X1 U1809 ( .A1(n12608), .A2(n13241), .B1(n12596), .B2(n13945), .ZN(
        n5141) );
  OAI22_X1 U1810 ( .A1(n12687), .A2(n13184), .B1(n12673), .B2(n13892), .ZN(
        n5378) );
  OAI22_X1 U1811 ( .A1(n12687), .A2(n13187), .B1(n12675), .B2(n13891), .ZN(
        n5379) );
  OAI22_X1 U1812 ( .A1(n12687), .A2(n13190), .B1(n12674), .B2(n13890), .ZN(
        n5380) );
  OAI22_X1 U1813 ( .A1(n12687), .A2(n13193), .B1(n12673), .B2(n13889), .ZN(
        n5381) );
  OAI22_X1 U1814 ( .A1(n12687), .A2(n13196), .B1(n12675), .B2(n13888), .ZN(
        n5382) );
  OAI22_X1 U1815 ( .A1(n12686), .A2(n13199), .B1(n12672), .B2(n13887), .ZN(
        n5383) );
  OAI22_X1 U1816 ( .A1(n12686), .A2(n13202), .B1(n1943), .B2(n13886), .ZN(
        n5384) );
  OAI22_X1 U1817 ( .A1(n12686), .A2(n13205), .B1(n1943), .B2(n13885), .ZN(
        n5385) );
  OAI22_X1 U1818 ( .A1(n12686), .A2(n13208), .B1(n12674), .B2(n13884), .ZN(
        n5386) );
  OAI22_X1 U1819 ( .A1(n12686), .A2(n13211), .B1(n12672), .B2(n13883), .ZN(
        n5387) );
  OAI22_X1 U1820 ( .A1(n12685), .A2(n13214), .B1(n12672), .B2(n13882), .ZN(
        n5388) );
  OAI22_X1 U1821 ( .A1(n12685), .A2(n13217), .B1(n1943), .B2(n13881), .ZN(
        n5389) );
  OAI22_X1 U1822 ( .A1(n12685), .A2(n13220), .B1(n1943), .B2(n13880), .ZN(
        n5390) );
  OAI22_X1 U1823 ( .A1(n12685), .A2(n13223), .B1(n1943), .B2(n13879), .ZN(
        n5391) );
  OAI22_X1 U1824 ( .A1(n12685), .A2(n13226), .B1(n1943), .B2(n13878), .ZN(
        n5392) );
  OAI22_X1 U1825 ( .A1(n12684), .A2(n13229), .B1(n1943), .B2(n13877), .ZN(
        n5393) );
  OAI22_X1 U1826 ( .A1(n12684), .A2(n13232), .B1(n12672), .B2(n13876), .ZN(
        n5394) );
  OAI22_X1 U1827 ( .A1(n12684), .A2(n13235), .B1(n12672), .B2(n13875), .ZN(
        n5395) );
  OAI22_X1 U1828 ( .A1(n12684), .A2(n13238), .B1(n12672), .B2(n13874), .ZN(
        n5396) );
  OAI22_X1 U1829 ( .A1(n12684), .A2(n13241), .B1(n12672), .B2(n13873), .ZN(
        n5397) );
  OAI22_X1 U1830 ( .A1(n12612), .A2(n13172), .B1(n1947), .B2(n13815), .ZN(
        n5118) );
  OAI22_X1 U1831 ( .A1(n12612), .A2(n13175), .B1(n1947), .B2(n13814), .ZN(
        n5119) );
  OAI22_X1 U1832 ( .A1(n12612), .A2(n13178), .B1(n1947), .B2(n13813), .ZN(
        n5120) );
  OAI22_X1 U1833 ( .A1(n12612), .A2(n13181), .B1(n1947), .B2(n13812), .ZN(
        n5121) );
  OAI22_X1 U1834 ( .A1(n12611), .A2(n13184), .B1(n1947), .B2(n13811), .ZN(
        n5122) );
  OAI22_X1 U1835 ( .A1(n12631), .A2(n13172), .B1(n12616), .B2(n13810), .ZN(
        n5182) );
  OAI22_X1 U1836 ( .A1(n12631), .A2(n13175), .B1(n12615), .B2(n13809), .ZN(
        n5183) );
  OAI22_X1 U1837 ( .A1(n12631), .A2(n13178), .B1(n12615), .B2(n13808), .ZN(
        n5184) );
  OAI22_X1 U1838 ( .A1(n12631), .A2(n13181), .B1(n1946), .B2(n13807), .ZN(
        n5185) );
  OAI22_X1 U1839 ( .A1(n12630), .A2(n13184), .B1(n1946), .B2(n13806), .ZN(
        n5186) );
  OAI22_X1 U1840 ( .A1(n12630), .A2(n13187), .B1(n1946), .B2(n13805), .ZN(
        n5187) );
  OAI22_X1 U1841 ( .A1(n12630), .A2(n13190), .B1(n1946), .B2(n13804), .ZN(
        n5188) );
  OAI22_X1 U1842 ( .A1(n12630), .A2(n13193), .B1(n1946), .B2(n13803), .ZN(
        n5189) );
  OAI22_X1 U1843 ( .A1(n12630), .A2(n13196), .B1(n12615), .B2(n13802), .ZN(
        n5190) );
  OAI22_X1 U1844 ( .A1(n12629), .A2(n13199), .B1(n12615), .B2(n13801), .ZN(
        n5191) );
  OAI22_X1 U1845 ( .A1(n12629), .A2(n13202), .B1(n12615), .B2(n13800), .ZN(
        n5192) );
  OAI22_X1 U1846 ( .A1(n12629), .A2(n13205), .B1(n12615), .B2(n13799), .ZN(
        n5193) );
  OAI22_X1 U1847 ( .A1(n12629), .A2(n13208), .B1(n12617), .B2(n13798), .ZN(
        n5194) );
  OAI22_X1 U1848 ( .A1(n12629), .A2(n13211), .B1(n12618), .B2(n13797), .ZN(
        n5195) );
  OAI22_X1 U1849 ( .A1(n12628), .A2(n13214), .B1(n12616), .B2(n13796), .ZN(
        n5196) );
  OAI22_X1 U1850 ( .A1(n12628), .A2(n13217), .B1(n12617), .B2(n13795), .ZN(
        n5197) );
  OAI22_X1 U1851 ( .A1(n12628), .A2(n13220), .B1(n12618), .B2(n13794), .ZN(
        n5198) );
  OAI22_X1 U1852 ( .A1(n12628), .A2(n13223), .B1(n12615), .B2(n13793), .ZN(
        n5199) );
  OAI22_X1 U1853 ( .A1(n12628), .A2(n13226), .B1(n1946), .B2(n13792), .ZN(
        n5200) );
  OAI22_X1 U1854 ( .A1(n12627), .A2(n13229), .B1(n1946), .B2(n13791), .ZN(
        n5201) );
  OAI22_X1 U1855 ( .A1(n12627), .A2(n13232), .B1(n1946), .B2(n13790), .ZN(
        n5202) );
  OAI22_X1 U1856 ( .A1(n12627), .A2(n13235), .B1(n1946), .B2(n13789), .ZN(
        n5203) );
  OAI22_X1 U1857 ( .A1(n12627), .A2(n13238), .B1(n1946), .B2(n13788), .ZN(
        n5204) );
  OAI22_X1 U1858 ( .A1(n12627), .A2(n13241), .B1(n1946), .B2(n13787), .ZN(
        n5205) );
  OAI22_X1 U1859 ( .A1(n12688), .A2(n13172), .B1(n1943), .B2(n13746), .ZN(
        n5374) );
  OAI22_X1 U1860 ( .A1(n12688), .A2(n13175), .B1(n1943), .B2(n13745), .ZN(
        n5375) );
  OAI22_X1 U1861 ( .A1(n12688), .A2(n13178), .B1(n1943), .B2(n13744), .ZN(
        n5376) );
  OAI22_X1 U1862 ( .A1(n12688), .A2(n13181), .B1(n1943), .B2(n13743), .ZN(
        n5377) );
  OAI22_X1 U1863 ( .A1(n12707), .A2(n13172), .B1(n12692), .B2(n13730), .ZN(
        n5438) );
  OAI22_X1 U1864 ( .A1(n12707), .A2(n13175), .B1(n12691), .B2(n13729), .ZN(
        n5439) );
  OAI22_X1 U1865 ( .A1(n12707), .A2(n13178), .B1(n12691), .B2(n13728), .ZN(
        n5440) );
  OAI22_X1 U1866 ( .A1(n12707), .A2(n13181), .B1(n1941), .B2(n13727), .ZN(
        n5441) );
  OAI22_X1 U1867 ( .A1(n12706), .A2(n13184), .B1(n1941), .B2(n13726), .ZN(
        n5442) );
  OAI22_X1 U1868 ( .A1(n12706), .A2(n13187), .B1(n1941), .B2(n13725), .ZN(
        n5443) );
  OAI22_X1 U1869 ( .A1(n12706), .A2(n13190), .B1(n1941), .B2(n13724), .ZN(
        n5444) );
  OAI22_X1 U1870 ( .A1(n12706), .A2(n13193), .B1(n1941), .B2(n13723), .ZN(
        n5445) );
  OAI22_X1 U1871 ( .A1(n12706), .A2(n13196), .B1(n12691), .B2(n13722), .ZN(
        n5446) );
  OAI22_X1 U1872 ( .A1(n12705), .A2(n13199), .B1(n12691), .B2(n13721), .ZN(
        n5447) );
  OAI22_X1 U1873 ( .A1(n12705), .A2(n13202), .B1(n12691), .B2(n13720), .ZN(
        n5448) );
  OAI22_X1 U1874 ( .A1(n12705), .A2(n13205), .B1(n12691), .B2(n13719), .ZN(
        n5449) );
  OAI22_X1 U1875 ( .A1(n12705), .A2(n13208), .B1(n12693), .B2(n13718), .ZN(
        n5450) );
  OAI22_X1 U1876 ( .A1(n12705), .A2(n13211), .B1(n12694), .B2(n13717), .ZN(
        n5451) );
  OAI22_X1 U1877 ( .A1(n12704), .A2(n13214), .B1(n12692), .B2(n13716), .ZN(
        n5452) );
  OAI22_X1 U1878 ( .A1(n12704), .A2(n13217), .B1(n12693), .B2(n13715), .ZN(
        n5453) );
  OAI22_X1 U1879 ( .A1(n12704), .A2(n13220), .B1(n12694), .B2(n13714), .ZN(
        n5454) );
  OAI22_X1 U1880 ( .A1(n12704), .A2(n13223), .B1(n12691), .B2(n13713), .ZN(
        n5455) );
  OAI22_X1 U1881 ( .A1(n12704), .A2(n13226), .B1(n1941), .B2(n13712), .ZN(
        n5456) );
  OAI22_X1 U1882 ( .A1(n12703), .A2(n13229), .B1(n1941), .B2(n13711), .ZN(
        n5457) );
  OAI22_X1 U1883 ( .A1(n12703), .A2(n13232), .B1(n1941), .B2(n13710), .ZN(
        n5458) );
  OAI22_X1 U1884 ( .A1(n12703), .A2(n13235), .B1(n1941), .B2(n13709), .ZN(
        n5459) );
  OAI22_X1 U1885 ( .A1(n12703), .A2(n13238), .B1(n1941), .B2(n13708), .ZN(
        n5460) );
  OAI22_X1 U1886 ( .A1(n12703), .A2(n13241), .B1(n1941), .B2(n13707), .ZN(
        n5461) );
  OAI22_X1 U1887 ( .A1(n12887), .A2(n13171), .B1(n12871), .B2(n13650), .ZN(
        n6014) );
  OAI22_X1 U1888 ( .A1(n12887), .A2(n13174), .B1(n12871), .B2(n13649), .ZN(
        n6015) );
  OAI22_X1 U1889 ( .A1(n12887), .A2(n13177), .B1(n12871), .B2(n13648), .ZN(
        n6016) );
  OAI22_X1 U1890 ( .A1(n12887), .A2(n13180), .B1(n12871), .B2(n13647), .ZN(
        n6017) );
  OAI22_X1 U1891 ( .A1(n12884), .A2(n13219), .B1(n1931), .B2(n13646), .ZN(
        n6030) );
  OAI22_X1 U1892 ( .A1(n12883), .A2(n13237), .B1(n1931), .B2(n13645), .ZN(
        n6036) );
  OAI22_X1 U1893 ( .A1(n12883), .A2(n13240), .B1(n1931), .B2(n13644), .ZN(
        n6037) );
  OAI22_X1 U1894 ( .A1(n12907), .A2(n13171), .B1(n12891), .B2(n13603), .ZN(
        n6078) );
  OAI22_X1 U1895 ( .A1(n12907), .A2(n13174), .B1(n12891), .B2(n13602), .ZN(
        n6079) );
  OAI22_X1 U1896 ( .A1(n12907), .A2(n13177), .B1(n12891), .B2(n13601), .ZN(
        n6080) );
  OAI22_X1 U1897 ( .A1(n12907), .A2(n13180), .B1(n12891), .B2(n13600), .ZN(
        n6081) );
  OAI22_X1 U1898 ( .A1(n12906), .A2(n13183), .B1(n12891), .B2(n13599), .ZN(
        n6082) );
  OAI22_X1 U1899 ( .A1(n12906), .A2(n13186), .B1(n12891), .B2(n13598), .ZN(
        n6083) );
  OAI22_X1 U1900 ( .A1(n12906), .A2(n13189), .B1(n12891), .B2(n13597), .ZN(
        n6084) );
  OAI22_X1 U1901 ( .A1(n12906), .A2(n13192), .B1(n12891), .B2(n13596), .ZN(
        n6085) );
  OAI22_X1 U1902 ( .A1(n12906), .A2(n13195), .B1(n12891), .B2(n13595), .ZN(
        n6086) );
  OAI22_X1 U1903 ( .A1(n12905), .A2(n13198), .B1(n12891), .B2(n13594), .ZN(
        n6087) );
  OAI22_X1 U1904 ( .A1(n12905), .A2(n13201), .B1(n12891), .B2(n13593), .ZN(
        n6088) );
  OAI22_X1 U1905 ( .A1(n12905), .A2(n13204), .B1(n12891), .B2(n13592), .ZN(
        n6089) );
  OAI22_X1 U1906 ( .A1(n12905), .A2(n13207), .B1(n12893), .B2(n13591), .ZN(
        n6090) );
  OAI22_X1 U1907 ( .A1(n12905), .A2(n13210), .B1(n12894), .B2(n13590), .ZN(
        n6091) );
  OAI22_X1 U1908 ( .A1(n12904), .A2(n13213), .B1(n12891), .B2(n13589), .ZN(
        n6092) );
  OAI22_X1 U1909 ( .A1(n12904), .A2(n13216), .B1(n12893), .B2(n13588), .ZN(
        n6093) );
  OAI22_X1 U1910 ( .A1(n12904), .A2(n13219), .B1(n12894), .B2(n13587), .ZN(
        n6094) );
  OAI22_X1 U1911 ( .A1(n12904), .A2(n13222), .B1(n12890), .B2(n13586), .ZN(
        n6095) );
  OAI22_X1 U1912 ( .A1(n12904), .A2(n13225), .B1(n1930), .B2(n13585), .ZN(
        n6096) );
  OAI22_X1 U1913 ( .A1(n12903), .A2(n13228), .B1(n1930), .B2(n13584), .ZN(
        n6097) );
  OAI22_X1 U1914 ( .A1(n12903), .A2(n13231), .B1(n1930), .B2(n13583), .ZN(
        n6098) );
  OAI22_X1 U1915 ( .A1(n12903), .A2(n13234), .B1(n1930), .B2(n13582), .ZN(
        n6099) );
  OAI22_X1 U1916 ( .A1(n12903), .A2(n13237), .B1(n1930), .B2(n13581), .ZN(
        n6100) );
  OAI22_X1 U1917 ( .A1(n12903), .A2(n13240), .B1(n1930), .B2(n13580), .ZN(
        n6101) );
  OAI22_X1 U1918 ( .A1(n12967), .A2(n13170), .B1(n12951), .B2(n13539), .ZN(
        n6270) );
  OAI22_X1 U1919 ( .A1(n12967), .A2(n13173), .B1(n12951), .B2(n13538), .ZN(
        n6271) );
  OAI22_X1 U1920 ( .A1(n12967), .A2(n13176), .B1(n12951), .B2(n13537), .ZN(
        n6272) );
  OAI22_X1 U1921 ( .A1(n12967), .A2(n13179), .B1(n12951), .B2(n13536), .ZN(
        n6273) );
  OAI22_X1 U1922 ( .A1(n12964), .A2(n13218), .B1(n1927), .B2(n13535), .ZN(
        n6286) );
  OAI22_X1 U1923 ( .A1(n12963), .A2(n13230), .B1(n1927), .B2(n13534), .ZN(
        n6290) );
  OAI22_X1 U1924 ( .A1(n12963), .A2(n13233), .B1(n1927), .B2(n13533), .ZN(
        n6291) );
  OAI22_X1 U1925 ( .A1(n12963), .A2(n13236), .B1(n1927), .B2(n13532), .ZN(
        n6292) );
  OAI22_X1 U1926 ( .A1(n12963), .A2(n13239), .B1(n1927), .B2(n13531), .ZN(
        n6293) );
  OAI22_X1 U1927 ( .A1(n12987), .A2(n13170), .B1(n12971), .B2(n13494), .ZN(
        n6334) );
  OAI22_X1 U1928 ( .A1(n12987), .A2(n13173), .B1(n12971), .B2(n13493), .ZN(
        n6335) );
  OAI22_X1 U1929 ( .A1(n12987), .A2(n13176), .B1(n12971), .B2(n13492), .ZN(
        n6336) );
  OAI22_X1 U1930 ( .A1(n12987), .A2(n13179), .B1(n12971), .B2(n13491), .ZN(
        n6337) );
  OAI22_X1 U1931 ( .A1(n12986), .A2(n13182), .B1(n12971), .B2(n13490), .ZN(
        n6338) );
  OAI22_X1 U1932 ( .A1(n12986), .A2(n13185), .B1(n12971), .B2(n13489), .ZN(
        n6339) );
  OAI22_X1 U1933 ( .A1(n12986), .A2(n13188), .B1(n12971), .B2(n13488), .ZN(
        n6340) );
  OAI22_X1 U1934 ( .A1(n12986), .A2(n13191), .B1(n12971), .B2(n13487), .ZN(
        n6341) );
  OAI22_X1 U1935 ( .A1(n12986), .A2(n13194), .B1(n12971), .B2(n13486), .ZN(
        n6342) );
  OAI22_X1 U1936 ( .A1(n12985), .A2(n13197), .B1(n12971), .B2(n13485), .ZN(
        n6343) );
  OAI22_X1 U1937 ( .A1(n12985), .A2(n13200), .B1(n12971), .B2(n13484), .ZN(
        n6344) );
  OAI22_X1 U1938 ( .A1(n12985), .A2(n13203), .B1(n12971), .B2(n13483), .ZN(
        n6345) );
  OAI22_X1 U1939 ( .A1(n12985), .A2(n13206), .B1(n12973), .B2(n13482), .ZN(
        n6346) );
  OAI22_X1 U1940 ( .A1(n12985), .A2(n13209), .B1(n12974), .B2(n13481), .ZN(
        n6347) );
  OAI22_X1 U1941 ( .A1(n12984), .A2(n13212), .B1(n12971), .B2(n13480), .ZN(
        n6348) );
  OAI22_X1 U1942 ( .A1(n12984), .A2(n13215), .B1(n12973), .B2(n13479), .ZN(
        n6349) );
  OAI22_X1 U1943 ( .A1(n12984), .A2(n13218), .B1(n12974), .B2(n13478), .ZN(
        n6350) );
  OAI22_X1 U1944 ( .A1(n12984), .A2(n13221), .B1(n12970), .B2(n13477), .ZN(
        n6351) );
  OAI22_X1 U1945 ( .A1(n12984), .A2(n13224), .B1(n1926), .B2(n13476), .ZN(
        n6352) );
  OAI22_X1 U1946 ( .A1(n12983), .A2(n13227), .B1(n1926), .B2(n13475), .ZN(
        n6353) );
  OAI22_X1 U1947 ( .A1(n12983), .A2(n13230), .B1(n1926), .B2(n13474), .ZN(
        n6354) );
  OAI22_X1 U1948 ( .A1(n12983), .A2(n13233), .B1(n1926), .B2(n13473), .ZN(
        n6355) );
  OAI22_X1 U1949 ( .A1(n12983), .A2(n13236), .B1(n1926), .B2(n13472), .ZN(
        n6356) );
  OAI22_X1 U1950 ( .A1(n12983), .A2(n13239), .B1(n1926), .B2(n13471), .ZN(
        n6357) );
  OAI22_X1 U1951 ( .A1(n13167), .A2(n13170), .B1(n13151), .B2(n13430), .ZN(
        n6910) );
  OAI22_X1 U1952 ( .A1(n13167), .A2(n13173), .B1(n13151), .B2(n13429), .ZN(
        n6911) );
  OAI22_X1 U1953 ( .A1(n13167), .A2(n13176), .B1(n13151), .B2(n13428), .ZN(
        n6912) );
  OAI22_X1 U1954 ( .A1(n13167), .A2(n13179), .B1(n13151), .B2(n13427), .ZN(
        n6913) );
  OAI22_X1 U1955 ( .A1(n13166), .A2(n13182), .B1(n13151), .B2(n13426), .ZN(
        n6914) );
  OAI22_X1 U1956 ( .A1(n13166), .A2(n13185), .B1(n13151), .B2(n13425), .ZN(
        n6915) );
  OAI22_X1 U1957 ( .A1(n13166), .A2(n13188), .B1(n13151), .B2(n13424), .ZN(
        n6916) );
  OAI22_X1 U1958 ( .A1(n13166), .A2(n13191), .B1(n13151), .B2(n13423), .ZN(
        n6917) );
  OAI22_X1 U1959 ( .A1(n13166), .A2(n13194), .B1(n13151), .B2(n13422), .ZN(
        n6918) );
  OAI22_X1 U1960 ( .A1(n13165), .A2(n13197), .B1(n13151), .B2(n13421), .ZN(
        n6919) );
  OAI22_X1 U1961 ( .A1(n13165), .A2(n13200), .B1(n13151), .B2(n13420), .ZN(
        n6920) );
  OAI22_X1 U1962 ( .A1(n13165), .A2(n13203), .B1(n13151), .B2(n13419), .ZN(
        n6921) );
  OAI22_X1 U1963 ( .A1(n13165), .A2(n13206), .B1(n13153), .B2(n13418), .ZN(
        n6922) );
  OAI22_X1 U1964 ( .A1(n13165), .A2(n13209), .B1(n13152), .B2(n13417), .ZN(
        n6923) );
  OAI22_X1 U1965 ( .A1(n13164), .A2(n13212), .B1(n13151), .B2(n13416), .ZN(
        n6924) );
  OAI22_X1 U1966 ( .A1(n13164), .A2(n13215), .B1(n13153), .B2(n13415), .ZN(
        n6925) );
  OAI22_X1 U1967 ( .A1(n13164), .A2(n13218), .B1(n13152), .B2(n13414), .ZN(
        n6926) );
  OAI22_X1 U1968 ( .A1(n13164), .A2(n13221), .B1(n13150), .B2(n13413), .ZN(
        n6927) );
  OAI22_X1 U1969 ( .A1(n13164), .A2(n13224), .B1(n1908), .B2(n13412), .ZN(
        n6928) );
  OAI22_X1 U1970 ( .A1(n13163), .A2(n13227), .B1(n1908), .B2(n13411), .ZN(
        n6929) );
  OAI22_X1 U1971 ( .A1(n13163), .A2(n13230), .B1(n1908), .B2(n13410), .ZN(
        n6930) );
  OAI22_X1 U1972 ( .A1(n13163), .A2(n13233), .B1(n1908), .B2(n13409), .ZN(
        n6931) );
  OAI22_X1 U1973 ( .A1(n13163), .A2(n13236), .B1(n1908), .B2(n13408), .ZN(
        n6932) );
  OAI22_X1 U1974 ( .A1(n13163), .A2(n13239), .B1(n1908), .B2(n13407), .ZN(
        n6933) );
  OAI22_X1 U1975 ( .A1(n12959), .A2(n13287), .B1(n12953), .B2(n14460), .ZN(
        n6309) );
  OAI22_X1 U1976 ( .A1(n12959), .A2(n13290), .B1(n12953), .B2(n14459), .ZN(
        n6310) );
  OAI22_X1 U1977 ( .A1(n12959), .A2(n13293), .B1(n12953), .B2(n14458), .ZN(
        n6311) );
  OAI22_X1 U1978 ( .A1(n12959), .A2(n13296), .B1(n12953), .B2(n14457), .ZN(
        n6312) );
  OAI22_X1 U1979 ( .A1(n13370), .A2(n13260), .B1(n13361), .B2(n14456), .ZN(
        n7004) );
  OAI22_X1 U1980 ( .A1(n13370), .A2(n13263), .B1(n13361), .B2(n14455), .ZN(
        n7005) );
  OAI22_X1 U1981 ( .A1(n13370), .A2(n13266), .B1(n13361), .B2(n14454), .ZN(
        n7006) );
  OAI22_X1 U1982 ( .A1(n13370), .A2(n13269), .B1(n13361), .B2(n14453), .ZN(
        n7007) );
  OAI22_X1 U1983 ( .A1(n13369), .A2(n13272), .B1(n13361), .B2(n14452), .ZN(
        n7008) );
  OAI22_X1 U1984 ( .A1(n13369), .A2(n13275), .B1(n13361), .B2(n14451), .ZN(
        n7009) );
  OAI22_X1 U1985 ( .A1(n13369), .A2(n13278), .B1(n13362), .B2(n14450), .ZN(
        n7010) );
  OAI22_X1 U1986 ( .A1(n13369), .A2(n13281), .B1(n13362), .B2(n14449), .ZN(
        n7011) );
  OAI22_X1 U1987 ( .A1(n13369), .A2(n13284), .B1(n13362), .B2(n14448), .ZN(
        n7012) );
  OAI22_X1 U1988 ( .A1(n13368), .A2(n13287), .B1(n13362), .B2(n14447), .ZN(
        n7013) );
  OAI22_X1 U1989 ( .A1(n13368), .A2(n13290), .B1(n13362), .B2(n14446), .ZN(
        n7014) );
  OAI22_X1 U1990 ( .A1(n13368), .A2(n13293), .B1(n13362), .B2(n14445), .ZN(
        n7015) );
  OAI22_X1 U1991 ( .A1(n13368), .A2(n13296), .B1(n13362), .B2(n14444), .ZN(
        n7016) );
  OAI22_X1 U1992 ( .A1(n13368), .A2(n13299), .B1(n13362), .B2(n14443), .ZN(
        n7017) );
  OAI22_X1 U1993 ( .A1(n13367), .A2(n13302), .B1(n13362), .B2(n14442), .ZN(
        n7018) );
  OAI22_X1 U1994 ( .A1(n13367), .A2(n13305), .B1(n13362), .B2(n14441), .ZN(
        n7019) );
  OAI22_X1 U1995 ( .A1(n13365), .A2(n13335), .B1(n13363), .B2(n14440), .ZN(
        n7029) );
  OAI22_X1 U1996 ( .A1(n13365), .A2(n13338), .B1(n13363), .B2(n14439), .ZN(
        n7030) );
  OAI22_X1 U1997 ( .A1(n13365), .A2(n13341), .B1(n13363), .B2(n14438), .ZN(
        n7031) );
  OAI22_X1 U1998 ( .A1(n13365), .A2(n13344), .B1(n13363), .B2(n14437), .ZN(
        n7032) );
  OAI22_X1 U1999 ( .A1(n13364), .A2(n13347), .B1(n13363), .B2(n14436), .ZN(
        n7033) );
  OAI22_X1 U2000 ( .A1(n13159), .A2(n13290), .B1(n13153), .B2(n14432), .ZN(
        n6950) );
  OAI22_X1 U2001 ( .A1(n13159), .A2(n13293), .B1(n13153), .B2(n14431), .ZN(
        n6951) );
  OAI22_X1 U2002 ( .A1(n13159), .A2(n13296), .B1(n13153), .B2(n14430), .ZN(
        n6952) );
  OAI22_X1 U2003 ( .A1(n13159), .A2(n13299), .B1(n13153), .B2(n14429), .ZN(
        n6953) );
  OAI22_X1 U2004 ( .A1(n13158), .A2(n13302), .B1(n13153), .B2(n14428), .ZN(
        n6954) );
  OAI22_X1 U2005 ( .A1(n13158), .A2(n13305), .B1(n13153), .B2(n14427), .ZN(
        n6955) );
  OAI22_X1 U2006 ( .A1(n13158), .A2(n13308), .B1(n13153), .B2(n14426), .ZN(
        n6956) );
  OAI22_X1 U2007 ( .A1(n13158), .A2(n13311), .B1(n13153), .B2(n14425), .ZN(
        n6957) );
  OAI22_X1 U2008 ( .A1(n13158), .A2(n13314), .B1(n13154), .B2(n14424), .ZN(
        n6958) );
  OAI22_X1 U2009 ( .A1(n13157), .A2(n13317), .B1(n13154), .B2(n14423), .ZN(
        n6959) );
  OAI22_X1 U2010 ( .A1(n13157), .A2(n13320), .B1(n13154), .B2(n14422), .ZN(
        n6960) );
  OAI22_X1 U2011 ( .A1(n13157), .A2(n13323), .B1(n13154), .B2(n14421), .ZN(
        n6961) );
  OAI22_X1 U2012 ( .A1(n13157), .A2(n13326), .B1(n13154), .B2(n14420), .ZN(
        n6962) );
  OAI22_X1 U2013 ( .A1(n13157), .A2(n13329), .B1(n13154), .B2(n14419), .ZN(
        n6963) );
  OAI22_X1 U2014 ( .A1(n13156), .A2(n13332), .B1(n13154), .B2(n14418), .ZN(
        n6964) );
  OAI22_X1 U2015 ( .A1(n13156), .A2(n13335), .B1(n13154), .B2(n14417), .ZN(
        n6965) );
  OAI22_X1 U2016 ( .A1(n13156), .A2(n13338), .B1(n13154), .B2(n14416), .ZN(
        n6966) );
  OAI22_X1 U2017 ( .A1(n13156), .A2(n13341), .B1(n13154), .B2(n14415), .ZN(
        n6967) );
  OAI22_X1 U2018 ( .A1(n13156), .A2(n13344), .B1(n13154), .B2(n14414), .ZN(
        n6968) );
  OAI22_X1 U2019 ( .A1(n13155), .A2(n13347), .B1(n13154), .B2(n14413), .ZN(
        n6969) );
  OAI22_X1 U2020 ( .A1(n13161), .A2(n13257), .B1(n13152), .B2(n14322), .ZN(
        n6939) );
  OAI22_X1 U2021 ( .A1(n13161), .A2(n13260), .B1(n13152), .B2(n14321), .ZN(
        n6940) );
  OAI22_X1 U2022 ( .A1(n13161), .A2(n13263), .B1(n13152), .B2(n14320), .ZN(
        n6941) );
  OAI22_X1 U2023 ( .A1(n13161), .A2(n13266), .B1(n13152), .B2(n14319), .ZN(
        n6942) );
  OAI22_X1 U2024 ( .A1(n13161), .A2(n13269), .B1(n13152), .B2(n14318), .ZN(
        n6943) );
  OAI22_X1 U2025 ( .A1(n13160), .A2(n13272), .B1(n13152), .B2(n14317), .ZN(
        n6944) );
  OAI22_X1 U2026 ( .A1(n13160), .A2(n13275), .B1(n13152), .B2(n14316), .ZN(
        n6945) );
  OAI22_X1 U2027 ( .A1(n13160), .A2(n13278), .B1(n13153), .B2(n14315), .ZN(
        n6946) );
  OAI22_X1 U2028 ( .A1(n13160), .A2(n13281), .B1(n13153), .B2(n14314), .ZN(
        n6947) );
  OAI22_X1 U2029 ( .A1(n13160), .A2(n13284), .B1(n13153), .B2(n14313), .ZN(
        n6948) );
  OAI22_X1 U2030 ( .A1(n13159), .A2(n13287), .B1(n13153), .B2(n14312), .ZN(
        n6949) );
  OAI22_X1 U2031 ( .A1(n13371), .A2(n13242), .B1(n13361), .B2(n14294), .ZN(
        n6998) );
  OAI22_X1 U2032 ( .A1(n13371), .A2(n13245), .B1(n13361), .B2(n14293), .ZN(
        n6999) );
  OAI22_X1 U2033 ( .A1(n13371), .A2(n13248), .B1(n13361), .B2(n14292), .ZN(
        n7000) );
  OAI22_X1 U2034 ( .A1(n13371), .A2(n13251), .B1(n13361), .B2(n14291), .ZN(
        n7001) );
  OAI22_X1 U2035 ( .A1(n13371), .A2(n13254), .B1(n13361), .B2(n14290), .ZN(
        n7002) );
  OAI22_X1 U2036 ( .A1(n13370), .A2(n13257), .B1(n13361), .B2(n14289), .ZN(
        n7003) );
  OAI22_X1 U2037 ( .A1(n13102), .A2(n13242), .B1(n13092), .B2(n14288), .ZN(
        n6742) );
  OAI22_X1 U2038 ( .A1(n13102), .A2(n13245), .B1(n13092), .B2(n14287), .ZN(
        n6743) );
  OAI22_X1 U2039 ( .A1(n13102), .A2(n13248), .B1(n13092), .B2(n14286), .ZN(
        n6744) );
  OAI22_X1 U2040 ( .A1(n13102), .A2(n13251), .B1(n13092), .B2(n14285), .ZN(
        n6745) );
  OAI22_X1 U2041 ( .A1(n13102), .A2(n13254), .B1(n13092), .B2(n14284), .ZN(
        n6746) );
  OAI22_X1 U2042 ( .A1(n13101), .A2(n13257), .B1(n13092), .B2(n14283), .ZN(
        n6747) );
  OAI22_X1 U2043 ( .A1(n13101), .A2(n13260), .B1(n13092), .B2(n14282), .ZN(
        n6748) );
  OAI22_X1 U2044 ( .A1(n13101), .A2(n13263), .B1(n13092), .B2(n14281), .ZN(
        n6749) );
  OAI22_X1 U2045 ( .A1(n13101), .A2(n13266), .B1(n13092), .B2(n14280), .ZN(
        n6750) );
  OAI22_X1 U2046 ( .A1(n13101), .A2(n13269), .B1(n13092), .B2(n14279), .ZN(
        n6751) );
  OAI22_X1 U2047 ( .A1(n13100), .A2(n13272), .B1(n13092), .B2(n14278), .ZN(
        n6752) );
  OAI22_X1 U2048 ( .A1(n13100), .A2(n13275), .B1(n13092), .B2(n14277), .ZN(
        n6753) );
  OAI22_X1 U2049 ( .A1(n13100), .A2(n13278), .B1(n13093), .B2(n14276), .ZN(
        n6754) );
  OAI22_X1 U2050 ( .A1(n13100), .A2(n13281), .B1(n13093), .B2(n14275), .ZN(
        n6755) );
  OAI22_X1 U2051 ( .A1(n13100), .A2(n13284), .B1(n13093), .B2(n14274), .ZN(
        n6756) );
  OAI22_X1 U2052 ( .A1(n13099), .A2(n13287), .B1(n13093), .B2(n14273), .ZN(
        n6757) );
  OAI22_X1 U2053 ( .A1(n13099), .A2(n13290), .B1(n13093), .B2(n14272), .ZN(
        n6758) );
  OAI22_X1 U2054 ( .A1(n13099), .A2(n13293), .B1(n13093), .B2(n14271), .ZN(
        n6759) );
  OAI22_X1 U2055 ( .A1(n13099), .A2(n13296), .B1(n13093), .B2(n14270), .ZN(
        n6760) );
  OAI22_X1 U2056 ( .A1(n13099), .A2(n13299), .B1(n13093), .B2(n14269), .ZN(
        n6761) );
  OAI22_X1 U2057 ( .A1(n13098), .A2(n13302), .B1(n13093), .B2(n14268), .ZN(
        n6762) );
  OAI22_X1 U2058 ( .A1(n13098), .A2(n13305), .B1(n13093), .B2(n14267), .ZN(
        n6763) );
  OAI22_X1 U2059 ( .A1(n13098), .A2(n13308), .B1(n13093), .B2(n14266), .ZN(
        n6764) );
  OAI22_X1 U2060 ( .A1(n13098), .A2(n13311), .B1(n13093), .B2(n14265), .ZN(
        n6765) );
  OAI22_X1 U2061 ( .A1(n13098), .A2(n13314), .B1(n13094), .B2(n14264), .ZN(
        n6766) );
  OAI22_X1 U2062 ( .A1(n13097), .A2(n13317), .B1(n13094), .B2(n14263), .ZN(
        n6767) );
  OAI22_X1 U2063 ( .A1(n13097), .A2(n13320), .B1(n13094), .B2(n14262), .ZN(
        n6768) );
  OAI22_X1 U2064 ( .A1(n13097), .A2(n13323), .B1(n13094), .B2(n14261), .ZN(
        n6769) );
  OAI22_X1 U2065 ( .A1(n13097), .A2(n13326), .B1(n13094), .B2(n14260), .ZN(
        n6770) );
  OAI22_X1 U2066 ( .A1(n13097), .A2(n13329), .B1(n13094), .B2(n14259), .ZN(
        n6771) );
  OAI22_X1 U2067 ( .A1(n13096), .A2(n13332), .B1(n13094), .B2(n14258), .ZN(
        n6772) );
  OAI22_X1 U2068 ( .A1(n13096), .A2(n13335), .B1(n13094), .B2(n14257), .ZN(
        n6773) );
  OAI22_X1 U2069 ( .A1(n13096), .A2(n13338), .B1(n13094), .B2(n14256), .ZN(
        n6774) );
  OAI22_X1 U2070 ( .A1(n13096), .A2(n13341), .B1(n13094), .B2(n14255), .ZN(
        n6775) );
  OAI22_X1 U2071 ( .A1(n13096), .A2(n13344), .B1(n13094), .B2(n14254), .ZN(
        n6776) );
  OAI22_X1 U2072 ( .A1(n13095), .A2(n13347), .B1(n13094), .B2(n14253), .ZN(
        n6777) );
  OAI22_X1 U2073 ( .A1(n13082), .A2(n13242), .B1(n13072), .B2(n14252), .ZN(
        n6678) );
  OAI22_X1 U2074 ( .A1(n13082), .A2(n13245), .B1(n13072), .B2(n14251), .ZN(
        n6679) );
  OAI22_X1 U2075 ( .A1(n13082), .A2(n13248), .B1(n13072), .B2(n14250), .ZN(
        n6680) );
  OAI22_X1 U2076 ( .A1(n13082), .A2(n13251), .B1(n13072), .B2(n14249), .ZN(
        n6681) );
  OAI22_X1 U2077 ( .A1(n13082), .A2(n13254), .B1(n13072), .B2(n14248), .ZN(
        n6682) );
  OAI22_X1 U2078 ( .A1(n13081), .A2(n13257), .B1(n13072), .B2(n14247), .ZN(
        n6683) );
  OAI22_X1 U2079 ( .A1(n13081), .A2(n13260), .B1(n13072), .B2(n14246), .ZN(
        n6684) );
  OAI22_X1 U2080 ( .A1(n13081), .A2(n13263), .B1(n13072), .B2(n14245), .ZN(
        n6685) );
  OAI22_X1 U2081 ( .A1(n13081), .A2(n13266), .B1(n13072), .B2(n14244), .ZN(
        n6686) );
  OAI22_X1 U2082 ( .A1(n13081), .A2(n13269), .B1(n13072), .B2(n14243), .ZN(
        n6687) );
  OAI22_X1 U2083 ( .A1(n13080), .A2(n13272), .B1(n13072), .B2(n14242), .ZN(
        n6688) );
  OAI22_X1 U2084 ( .A1(n13080), .A2(n13275), .B1(n13072), .B2(n14241), .ZN(
        n6689) );
  OAI22_X1 U2085 ( .A1(n13080), .A2(n13278), .B1(n13073), .B2(n14240), .ZN(
        n6690) );
  OAI22_X1 U2086 ( .A1(n13080), .A2(n13281), .B1(n13073), .B2(n14239), .ZN(
        n6691) );
  OAI22_X1 U2087 ( .A1(n13080), .A2(n13284), .B1(n13073), .B2(n14238), .ZN(
        n6692) );
  OAI22_X1 U2088 ( .A1(n13079), .A2(n13287), .B1(n13073), .B2(n14237), .ZN(
        n6693) );
  OAI22_X1 U2089 ( .A1(n13079), .A2(n13290), .B1(n13073), .B2(n14236), .ZN(
        n6694) );
  OAI22_X1 U2090 ( .A1(n13079), .A2(n13293), .B1(n13073), .B2(n14235), .ZN(
        n6695) );
  OAI22_X1 U2091 ( .A1(n13079), .A2(n13296), .B1(n13073), .B2(n14234), .ZN(
        n6696) );
  OAI22_X1 U2092 ( .A1(n13079), .A2(n13299), .B1(n13073), .B2(n14233), .ZN(
        n6697) );
  OAI22_X1 U2093 ( .A1(n13078), .A2(n13302), .B1(n13073), .B2(n14232), .ZN(
        n6698) );
  OAI22_X1 U2094 ( .A1(n13078), .A2(n13305), .B1(n13073), .B2(n14231), .ZN(
        n6699) );
  OAI22_X1 U2095 ( .A1(n13078), .A2(n13308), .B1(n13073), .B2(n14230), .ZN(
        n6700) );
  OAI22_X1 U2096 ( .A1(n13078), .A2(n13311), .B1(n13073), .B2(n14229), .ZN(
        n6701) );
  OAI22_X1 U2097 ( .A1(n13078), .A2(n13314), .B1(n13074), .B2(n14228), .ZN(
        n6702) );
  OAI22_X1 U2098 ( .A1(n13077), .A2(n13317), .B1(n13074), .B2(n14227), .ZN(
        n6703) );
  OAI22_X1 U2099 ( .A1(n13077), .A2(n13320), .B1(n13074), .B2(n14226), .ZN(
        n6704) );
  OAI22_X1 U2100 ( .A1(n13077), .A2(n13323), .B1(n13074), .B2(n14225), .ZN(
        n6705) );
  OAI22_X1 U2101 ( .A1(n13077), .A2(n13326), .B1(n13074), .B2(n14224), .ZN(
        n6706) );
  OAI22_X1 U2102 ( .A1(n13077), .A2(n13329), .B1(n13074), .B2(n14223), .ZN(
        n6707) );
  OAI22_X1 U2103 ( .A1(n13076), .A2(n13332), .B1(n13074), .B2(n14222), .ZN(
        n6708) );
  OAI22_X1 U2104 ( .A1(n13076), .A2(n13335), .B1(n13074), .B2(n14221), .ZN(
        n6709) );
  OAI22_X1 U2105 ( .A1(n13076), .A2(n13338), .B1(n13074), .B2(n14220), .ZN(
        n6710) );
  OAI22_X1 U2106 ( .A1(n13076), .A2(n13341), .B1(n13074), .B2(n14219), .ZN(
        n6711) );
  OAI22_X1 U2107 ( .A1(n13076), .A2(n13344), .B1(n13074), .B2(n14218), .ZN(
        n6712) );
  OAI22_X1 U2108 ( .A1(n13075), .A2(n13347), .B1(n13074), .B2(n14217), .ZN(
        n6713) );
  OAI22_X1 U2109 ( .A1(n12604), .A2(n13292), .B1(n12598), .B2(n14106), .ZN(
        n5158) );
  OAI22_X1 U2110 ( .A1(n12604), .A2(n13295), .B1(n12598), .B2(n14105), .ZN(
        n5159) );
  OAI22_X1 U2111 ( .A1(n12604), .A2(n13298), .B1(n12598), .B2(n14104), .ZN(
        n5160) );
  OAI22_X1 U2112 ( .A1(n12604), .A2(n13301), .B1(n12598), .B2(n14103), .ZN(
        n5161) );
  OAI22_X1 U2113 ( .A1(n12603), .A2(n13304), .B1(n12598), .B2(n14102), .ZN(
        n5162) );
  OAI22_X1 U2114 ( .A1(n12603), .A2(n13307), .B1(n12598), .B2(n14101), .ZN(
        n5163) );
  OAI22_X1 U2115 ( .A1(n12603), .A2(n13310), .B1(n12598), .B2(n14100), .ZN(
        n5164) );
  OAI22_X1 U2116 ( .A1(n12603), .A2(n13313), .B1(n12598), .B2(n14099), .ZN(
        n5165) );
  OAI22_X1 U2117 ( .A1(n12603), .A2(n13316), .B1(n12599), .B2(n14098), .ZN(
        n5166) );
  OAI22_X1 U2118 ( .A1(n12602), .A2(n13319), .B1(n12599), .B2(n14097), .ZN(
        n5167) );
  OAI22_X1 U2119 ( .A1(n12602), .A2(n13322), .B1(n12599), .B2(n14096), .ZN(
        n5168) );
  OAI22_X1 U2120 ( .A1(n12602), .A2(n13325), .B1(n12599), .B2(n14095), .ZN(
        n5169) );
  OAI22_X1 U2121 ( .A1(n12602), .A2(n13328), .B1(n12599), .B2(n14094), .ZN(
        n5170) );
  OAI22_X1 U2122 ( .A1(n12602), .A2(n13331), .B1(n12599), .B2(n14093), .ZN(
        n5171) );
  OAI22_X1 U2123 ( .A1(n12601), .A2(n13334), .B1(n12599), .B2(n14092), .ZN(
        n5172) );
  OAI22_X1 U2124 ( .A1(n12601), .A2(n13337), .B1(n12599), .B2(n14091), .ZN(
        n5173) );
  OAI22_X1 U2125 ( .A1(n12601), .A2(n13340), .B1(n12599), .B2(n14090), .ZN(
        n5174) );
  OAI22_X1 U2126 ( .A1(n12601), .A2(n13343), .B1(n12599), .B2(n14089), .ZN(
        n5175) );
  OAI22_X1 U2127 ( .A1(n12601), .A2(n13346), .B1(n12599), .B2(n14088), .ZN(
        n5176) );
  OAI22_X1 U2128 ( .A1(n12600), .A2(n13349), .B1(n12599), .B2(n14087), .ZN(
        n5177) );
  OAI22_X1 U2129 ( .A1(n12683), .A2(n13256), .B1(n12673), .B2(n14059), .ZN(
        n5402) );
  OAI22_X1 U2130 ( .A1(n12682), .A2(n13259), .B1(n12673), .B2(n14058), .ZN(
        n5403) );
  OAI22_X1 U2131 ( .A1(n12682), .A2(n13262), .B1(n12673), .B2(n14057), .ZN(
        n5404) );
  OAI22_X1 U2132 ( .A1(n12682), .A2(n13265), .B1(n12673), .B2(n14056), .ZN(
        n5405) );
  OAI22_X1 U2133 ( .A1(n12682), .A2(n13268), .B1(n12673), .B2(n14055), .ZN(
        n5406) );
  OAI22_X1 U2134 ( .A1(n12682), .A2(n13271), .B1(n12673), .B2(n14054), .ZN(
        n5407) );
  OAI22_X1 U2135 ( .A1(n12681), .A2(n13274), .B1(n12673), .B2(n14053), .ZN(
        n5408) );
  OAI22_X1 U2136 ( .A1(n12681), .A2(n13277), .B1(n12673), .B2(n14052), .ZN(
        n5409) );
  OAI22_X1 U2137 ( .A1(n12681), .A2(n13280), .B1(n12674), .B2(n14051), .ZN(
        n5410) );
  OAI22_X1 U2138 ( .A1(n12681), .A2(n13283), .B1(n12674), .B2(n14050), .ZN(
        n5411) );
  OAI22_X1 U2139 ( .A1(n12681), .A2(n13286), .B1(n12674), .B2(n14049), .ZN(
        n5412) );
  OAI22_X1 U2140 ( .A1(n12680), .A2(n13289), .B1(n12674), .B2(n14048), .ZN(
        n5413) );
  OAI22_X1 U2141 ( .A1(n12680), .A2(n13292), .B1(n12674), .B2(n14047), .ZN(
        n5414) );
  OAI22_X1 U2142 ( .A1(n12680), .A2(n13295), .B1(n12674), .B2(n14046), .ZN(
        n5415) );
  OAI22_X1 U2143 ( .A1(n12680), .A2(n13298), .B1(n12674), .B2(n14045), .ZN(
        n5416) );
  OAI22_X1 U2144 ( .A1(n12680), .A2(n13301), .B1(n12674), .B2(n14044), .ZN(
        n5417) );
  OAI22_X1 U2145 ( .A1(n12679), .A2(n13304), .B1(n12674), .B2(n14043), .ZN(
        n5418) );
  OAI22_X1 U2146 ( .A1(n12679), .A2(n13307), .B1(n12674), .B2(n14042), .ZN(
        n5419) );
  OAI22_X1 U2147 ( .A1(n12679), .A2(n13310), .B1(n12674), .B2(n14041), .ZN(
        n5420) );
  OAI22_X1 U2148 ( .A1(n12679), .A2(n13313), .B1(n12674), .B2(n14040), .ZN(
        n5421) );
  OAI22_X1 U2149 ( .A1(n12679), .A2(n13316), .B1(n12675), .B2(n14039), .ZN(
        n5422) );
  OAI22_X1 U2150 ( .A1(n12678), .A2(n13319), .B1(n12675), .B2(n14038), .ZN(
        n5423) );
  OAI22_X1 U2151 ( .A1(n12678), .A2(n13322), .B1(n12675), .B2(n14037), .ZN(
        n5424) );
  OAI22_X1 U2152 ( .A1(n12678), .A2(n13325), .B1(n12675), .B2(n14036), .ZN(
        n5425) );
  OAI22_X1 U2153 ( .A1(n12607), .A2(n13244), .B1(n12597), .B2(n13944), .ZN(
        n5142) );
  OAI22_X1 U2154 ( .A1(n12607), .A2(n13247), .B1(n12597), .B2(n13943), .ZN(
        n5143) );
  OAI22_X1 U2155 ( .A1(n12607), .A2(n13250), .B1(n12597), .B2(n13942), .ZN(
        n5144) );
  OAI22_X1 U2156 ( .A1(n12607), .A2(n13253), .B1(n12597), .B2(n13941), .ZN(
        n5145) );
  OAI22_X1 U2157 ( .A1(n12607), .A2(n13256), .B1(n12597), .B2(n13940), .ZN(
        n5146) );
  OAI22_X1 U2158 ( .A1(n12606), .A2(n13259), .B1(n12597), .B2(n13939), .ZN(
        n5147) );
  OAI22_X1 U2159 ( .A1(n12606), .A2(n13262), .B1(n12597), .B2(n13938), .ZN(
        n5148) );
  OAI22_X1 U2160 ( .A1(n12606), .A2(n13265), .B1(n12597), .B2(n13937), .ZN(
        n5149) );
  OAI22_X1 U2161 ( .A1(n12606), .A2(n13268), .B1(n12597), .B2(n13936), .ZN(
        n5150) );
  OAI22_X1 U2162 ( .A1(n12606), .A2(n13271), .B1(n12597), .B2(n13935), .ZN(
        n5151) );
  OAI22_X1 U2163 ( .A1(n12605), .A2(n13274), .B1(n12597), .B2(n13934), .ZN(
        n5152) );
  OAI22_X1 U2164 ( .A1(n12605), .A2(n13277), .B1(n12597), .B2(n13933), .ZN(
        n5153) );
  OAI22_X1 U2165 ( .A1(n12605), .A2(n13280), .B1(n12598), .B2(n13932), .ZN(
        n5154) );
  OAI22_X1 U2166 ( .A1(n12605), .A2(n13283), .B1(n12598), .B2(n13931), .ZN(
        n5155) );
  OAI22_X1 U2167 ( .A1(n12605), .A2(n13286), .B1(n12598), .B2(n13930), .ZN(
        n5156) );
  OAI22_X1 U2168 ( .A1(n12604), .A2(n13289), .B1(n12598), .B2(n13929), .ZN(
        n5157) );
  OAI22_X1 U2169 ( .A1(n12683), .A2(n13244), .B1(n12673), .B2(n13872), .ZN(
        n5398) );
  OAI22_X1 U2170 ( .A1(n12683), .A2(n13247), .B1(n12673), .B2(n13871), .ZN(
        n5399) );
  OAI22_X1 U2171 ( .A1(n12683), .A2(n13250), .B1(n12673), .B2(n13870), .ZN(
        n5400) );
  OAI22_X1 U2172 ( .A1(n12683), .A2(n13253), .B1(n12673), .B2(n13869), .ZN(
        n5401) );
  OAI22_X1 U2173 ( .A1(n12626), .A2(n13244), .B1(n12616), .B2(n13786), .ZN(
        n5206) );
  OAI22_X1 U2174 ( .A1(n12626), .A2(n13247), .B1(n12616), .B2(n13785), .ZN(
        n5207) );
  OAI22_X1 U2175 ( .A1(n12626), .A2(n13250), .B1(n12616), .B2(n13784), .ZN(
        n5208) );
  OAI22_X1 U2176 ( .A1(n12626), .A2(n13253), .B1(n12616), .B2(n13783), .ZN(
        n5209) );
  OAI22_X1 U2177 ( .A1(n12626), .A2(n13256), .B1(n12616), .B2(n13782), .ZN(
        n5210) );
  OAI22_X1 U2178 ( .A1(n12625), .A2(n13259), .B1(n12616), .B2(n13781), .ZN(
        n5211) );
  OAI22_X1 U2179 ( .A1(n12625), .A2(n13262), .B1(n12616), .B2(n13780), .ZN(
        n5212) );
  OAI22_X1 U2180 ( .A1(n12625), .A2(n13265), .B1(n12616), .B2(n13779), .ZN(
        n5213) );
  OAI22_X1 U2181 ( .A1(n12625), .A2(n13268), .B1(n12616), .B2(n13778), .ZN(
        n5214) );
  OAI22_X1 U2182 ( .A1(n12625), .A2(n13271), .B1(n12616), .B2(n13777), .ZN(
        n5215) );
  OAI22_X1 U2183 ( .A1(n12624), .A2(n13274), .B1(n12616), .B2(n13776), .ZN(
        n5216) );
  OAI22_X1 U2184 ( .A1(n12624), .A2(n13277), .B1(n12616), .B2(n13775), .ZN(
        n5217) );
  OAI22_X1 U2185 ( .A1(n12624), .A2(n13280), .B1(n12617), .B2(n13774), .ZN(
        n5218) );
  OAI22_X1 U2186 ( .A1(n12624), .A2(n13283), .B1(n12617), .B2(n13773), .ZN(
        n5219) );
  OAI22_X1 U2187 ( .A1(n12624), .A2(n13286), .B1(n12617), .B2(n13772), .ZN(
        n5220) );
  OAI22_X1 U2188 ( .A1(n12623), .A2(n13289), .B1(n12617), .B2(n13771), .ZN(
        n5221) );
  OAI22_X1 U2189 ( .A1(n12623), .A2(n13292), .B1(n12617), .B2(n13770), .ZN(
        n5222) );
  OAI22_X1 U2190 ( .A1(n12623), .A2(n13295), .B1(n12617), .B2(n13769), .ZN(
        n5223) );
  OAI22_X1 U2191 ( .A1(n12623), .A2(n13298), .B1(n12617), .B2(n13768), .ZN(
        n5224) );
  OAI22_X1 U2192 ( .A1(n12623), .A2(n13301), .B1(n12617), .B2(n13767), .ZN(
        n5225) );
  OAI22_X1 U2193 ( .A1(n12622), .A2(n13304), .B1(n12617), .B2(n13766), .ZN(
        n5226) );
  OAI22_X1 U2194 ( .A1(n12622), .A2(n13307), .B1(n12617), .B2(n13765), .ZN(
        n5227) );
  OAI22_X1 U2195 ( .A1(n12622), .A2(n13310), .B1(n12617), .B2(n13764), .ZN(
        n5228) );
  OAI22_X1 U2196 ( .A1(n12622), .A2(n13313), .B1(n12617), .B2(n13763), .ZN(
        n5229) );
  OAI22_X1 U2197 ( .A1(n12622), .A2(n13316), .B1(n12618), .B2(n13762), .ZN(
        n5230) );
  OAI22_X1 U2198 ( .A1(n12621), .A2(n13319), .B1(n12618), .B2(n13761), .ZN(
        n5231) );
  OAI22_X1 U2199 ( .A1(n12621), .A2(n13322), .B1(n12618), .B2(n13760), .ZN(
        n5232) );
  OAI22_X1 U2200 ( .A1(n12621), .A2(n13325), .B1(n12618), .B2(n13759), .ZN(
        n5233) );
  OAI22_X1 U2201 ( .A1(n12621), .A2(n13328), .B1(n12618), .B2(n13758), .ZN(
        n5234) );
  OAI22_X1 U2202 ( .A1(n12621), .A2(n13331), .B1(n12618), .B2(n13757), .ZN(
        n5235) );
  OAI22_X1 U2203 ( .A1(n12620), .A2(n13334), .B1(n12618), .B2(n13756), .ZN(
        n5236) );
  OAI22_X1 U2204 ( .A1(n12620), .A2(n13337), .B1(n12618), .B2(n13755), .ZN(
        n5237) );
  OAI22_X1 U2205 ( .A1(n12620), .A2(n13340), .B1(n12618), .B2(n13754), .ZN(
        n5238) );
  OAI22_X1 U2206 ( .A1(n12620), .A2(n13343), .B1(n12618), .B2(n13753), .ZN(
        n5239) );
  OAI22_X1 U2207 ( .A1(n12620), .A2(n13346), .B1(n12618), .B2(n13752), .ZN(
        n5240) );
  OAI22_X1 U2208 ( .A1(n12619), .A2(n13349), .B1(n12618), .B2(n13751), .ZN(
        n5241) );
  OAI22_X1 U2209 ( .A1(n12678), .A2(n13328), .B1(n12675), .B2(n13742), .ZN(
        n5426) );
  OAI22_X1 U2210 ( .A1(n12678), .A2(n13331), .B1(n12675), .B2(n13741), .ZN(
        n5427) );
  OAI22_X1 U2211 ( .A1(n12677), .A2(n13334), .B1(n12675), .B2(n13740), .ZN(
        n5428) );
  OAI22_X1 U2212 ( .A1(n12677), .A2(n13337), .B1(n12675), .B2(n13739), .ZN(
        n5429) );
  OAI22_X1 U2213 ( .A1(n12677), .A2(n13340), .B1(n12675), .B2(n13738), .ZN(
        n5430) );
  OAI22_X1 U2214 ( .A1(n12677), .A2(n13343), .B1(n12675), .B2(n13737), .ZN(
        n5431) );
  OAI22_X1 U2215 ( .A1(n12677), .A2(n13346), .B1(n12675), .B2(n13736), .ZN(
        n5432) );
  OAI22_X1 U2216 ( .A1(n12676), .A2(n13349), .B1(n12675), .B2(n13735), .ZN(
        n5433) );
  OAI22_X1 U2217 ( .A1(n12702), .A2(n13244), .B1(n12692), .B2(n13706), .ZN(
        n5462) );
  OAI22_X1 U2218 ( .A1(n12702), .A2(n13247), .B1(n12692), .B2(n13705), .ZN(
        n5463) );
  OAI22_X1 U2219 ( .A1(n12702), .A2(n13250), .B1(n12692), .B2(n13704), .ZN(
        n5464) );
  OAI22_X1 U2220 ( .A1(n12702), .A2(n13253), .B1(n12692), .B2(n13703), .ZN(
        n5465) );
  OAI22_X1 U2221 ( .A1(n12702), .A2(n13256), .B1(n12692), .B2(n13702), .ZN(
        n5466) );
  OAI22_X1 U2222 ( .A1(n12701), .A2(n13259), .B1(n12692), .B2(n13701), .ZN(
        n5467) );
  OAI22_X1 U2223 ( .A1(n12701), .A2(n13262), .B1(n12692), .B2(n13700), .ZN(
        n5468) );
  OAI22_X1 U2224 ( .A1(n12701), .A2(n13265), .B1(n12692), .B2(n13699), .ZN(
        n5469) );
  OAI22_X1 U2225 ( .A1(n12701), .A2(n13268), .B1(n12692), .B2(n13698), .ZN(
        n5470) );
  OAI22_X1 U2226 ( .A1(n12701), .A2(n13271), .B1(n12692), .B2(n13697), .ZN(
        n5471) );
  OAI22_X1 U2227 ( .A1(n12700), .A2(n13274), .B1(n12692), .B2(n13696), .ZN(
        n5472) );
  OAI22_X1 U2228 ( .A1(n12700), .A2(n13277), .B1(n12692), .B2(n13695), .ZN(
        n5473) );
  OAI22_X1 U2229 ( .A1(n12700), .A2(n13280), .B1(n12693), .B2(n13694), .ZN(
        n5474) );
  OAI22_X1 U2230 ( .A1(n12700), .A2(n13283), .B1(n12693), .B2(n13693), .ZN(
        n5475) );
  OAI22_X1 U2231 ( .A1(n12700), .A2(n13286), .B1(n12693), .B2(n13692), .ZN(
        n5476) );
  OAI22_X1 U2232 ( .A1(n12699), .A2(n13289), .B1(n12693), .B2(n13691), .ZN(
        n5477) );
  OAI22_X1 U2233 ( .A1(n12699), .A2(n13292), .B1(n12693), .B2(n13690), .ZN(
        n5478) );
  OAI22_X1 U2234 ( .A1(n12699), .A2(n13295), .B1(n12693), .B2(n13689), .ZN(
        n5479) );
  OAI22_X1 U2235 ( .A1(n12699), .A2(n13298), .B1(n12693), .B2(n13688), .ZN(
        n5480) );
  OAI22_X1 U2236 ( .A1(n12699), .A2(n13301), .B1(n12693), .B2(n13687), .ZN(
        n5481) );
  OAI22_X1 U2237 ( .A1(n12698), .A2(n13304), .B1(n12693), .B2(n13686), .ZN(
        n5482) );
  OAI22_X1 U2238 ( .A1(n12698), .A2(n13307), .B1(n12693), .B2(n13685), .ZN(
        n5483) );
  OAI22_X1 U2239 ( .A1(n12698), .A2(n13310), .B1(n12693), .B2(n13684), .ZN(
        n5484) );
  OAI22_X1 U2240 ( .A1(n12698), .A2(n13313), .B1(n12693), .B2(n13683), .ZN(
        n5485) );
  OAI22_X1 U2241 ( .A1(n12698), .A2(n13316), .B1(n12694), .B2(n13682), .ZN(
        n5486) );
  OAI22_X1 U2242 ( .A1(n12697), .A2(n13319), .B1(n12694), .B2(n13681), .ZN(
        n5487) );
  OAI22_X1 U2243 ( .A1(n12697), .A2(n13322), .B1(n12694), .B2(n13680), .ZN(
        n5488) );
  OAI22_X1 U2244 ( .A1(n12697), .A2(n13325), .B1(n12694), .B2(n13679), .ZN(
        n5489) );
  OAI22_X1 U2245 ( .A1(n12697), .A2(n13328), .B1(n12694), .B2(n13678), .ZN(
        n5490) );
  OAI22_X1 U2246 ( .A1(n12697), .A2(n13331), .B1(n12694), .B2(n13677), .ZN(
        n5491) );
  OAI22_X1 U2247 ( .A1(n12696), .A2(n13334), .B1(n12694), .B2(n13676), .ZN(
        n5492) );
  OAI22_X1 U2248 ( .A1(n12696), .A2(n13337), .B1(n12694), .B2(n13675), .ZN(
        n5493) );
  OAI22_X1 U2249 ( .A1(n12696), .A2(n13340), .B1(n12694), .B2(n13674), .ZN(
        n5494) );
  OAI22_X1 U2250 ( .A1(n12696), .A2(n13343), .B1(n12694), .B2(n13673), .ZN(
        n5495) );
  OAI22_X1 U2251 ( .A1(n12696), .A2(n13346), .B1(n12694), .B2(n13672), .ZN(
        n5496) );
  OAI22_X1 U2252 ( .A1(n12695), .A2(n13349), .B1(n12694), .B2(n13671), .ZN(
        n5497) );
  OAI22_X1 U2253 ( .A1(n12882), .A2(n13243), .B1(n12872), .B2(n13643), .ZN(
        n6038) );
  OAI22_X1 U2254 ( .A1(n12882), .A2(n13246), .B1(n12872), .B2(n13642), .ZN(
        n6039) );
  OAI22_X1 U2255 ( .A1(n12882), .A2(n13249), .B1(n12872), .B2(n13641), .ZN(
        n6040) );
  OAI22_X1 U2256 ( .A1(n12882), .A2(n13252), .B1(n12872), .B2(n13640), .ZN(
        n6041) );
  OAI22_X1 U2257 ( .A1(n12882), .A2(n13255), .B1(n12872), .B2(n13639), .ZN(
        n6042) );
  OAI22_X1 U2258 ( .A1(n12881), .A2(n13258), .B1(n12872), .B2(n13638), .ZN(
        n6043) );
  OAI22_X1 U2259 ( .A1(n12881), .A2(n13261), .B1(n12872), .B2(n13637), .ZN(
        n6044) );
  OAI22_X1 U2260 ( .A1(n12881), .A2(n13264), .B1(n12872), .B2(n13636), .ZN(
        n6045) );
  OAI22_X1 U2261 ( .A1(n12881), .A2(n13267), .B1(n12872), .B2(n13635), .ZN(
        n6046) );
  OAI22_X1 U2262 ( .A1(n12881), .A2(n13270), .B1(n12872), .B2(n13634), .ZN(
        n6047) );
  OAI22_X1 U2263 ( .A1(n12880), .A2(n13273), .B1(n12872), .B2(n13633), .ZN(
        n6048) );
  OAI22_X1 U2264 ( .A1(n12880), .A2(n13276), .B1(n12872), .B2(n13632), .ZN(
        n6049) );
  OAI22_X1 U2265 ( .A1(n12880), .A2(n13279), .B1(n12873), .B2(n13631), .ZN(
        n6050) );
  OAI22_X1 U2266 ( .A1(n12880), .A2(n13282), .B1(n12873), .B2(n13630), .ZN(
        n6051) );
  OAI22_X1 U2267 ( .A1(n12880), .A2(n13285), .B1(n12873), .B2(n13629), .ZN(
        n6052) );
  OAI22_X1 U2268 ( .A1(n12879), .A2(n13288), .B1(n12873), .B2(n13628), .ZN(
        n6053) );
  OAI22_X1 U2269 ( .A1(n12879), .A2(n13291), .B1(n12873), .B2(n13627), .ZN(
        n6054) );
  OAI22_X1 U2270 ( .A1(n12879), .A2(n13294), .B1(n12873), .B2(n13626), .ZN(
        n6055) );
  OAI22_X1 U2271 ( .A1(n12879), .A2(n13297), .B1(n12873), .B2(n13625), .ZN(
        n6056) );
  OAI22_X1 U2272 ( .A1(n12879), .A2(n13300), .B1(n12873), .B2(n13624), .ZN(
        n6057) );
  OAI22_X1 U2273 ( .A1(n12878), .A2(n13303), .B1(n12873), .B2(n13623), .ZN(
        n6058) );
  OAI22_X1 U2274 ( .A1(n12878), .A2(n13306), .B1(n12873), .B2(n13622), .ZN(
        n6059) );
  OAI22_X1 U2275 ( .A1(n12878), .A2(n13309), .B1(n12873), .B2(n13621), .ZN(
        n6060) );
  OAI22_X1 U2276 ( .A1(n12878), .A2(n13312), .B1(n12873), .B2(n13620), .ZN(
        n6061) );
  OAI22_X1 U2277 ( .A1(n12878), .A2(n13315), .B1(n12874), .B2(n13619), .ZN(
        n6062) );
  OAI22_X1 U2278 ( .A1(n12877), .A2(n13318), .B1(n12874), .B2(n13618), .ZN(
        n6063) );
  OAI22_X1 U2279 ( .A1(n12877), .A2(n13321), .B1(n12874), .B2(n13617), .ZN(
        n6064) );
  OAI22_X1 U2280 ( .A1(n12877), .A2(n13324), .B1(n12874), .B2(n13616), .ZN(
        n6065) );
  OAI22_X1 U2281 ( .A1(n12877), .A2(n13327), .B1(n12874), .B2(n13615), .ZN(
        n6066) );
  OAI22_X1 U2282 ( .A1(n12877), .A2(n13330), .B1(n12874), .B2(n13614), .ZN(
        n6067) );
  OAI22_X1 U2283 ( .A1(n12876), .A2(n13333), .B1(n12874), .B2(n13613), .ZN(
        n6068) );
  OAI22_X1 U2284 ( .A1(n12876), .A2(n13336), .B1(n12874), .B2(n13612), .ZN(
        n6069) );
  OAI22_X1 U2285 ( .A1(n12876), .A2(n13339), .B1(n12874), .B2(n13611), .ZN(
        n6070) );
  OAI22_X1 U2286 ( .A1(n12876), .A2(n13342), .B1(n12874), .B2(n13610), .ZN(
        n6071) );
  OAI22_X1 U2287 ( .A1(n12876), .A2(n13345), .B1(n12874), .B2(n13609), .ZN(
        n6072) );
  OAI22_X1 U2288 ( .A1(n12875), .A2(n13348), .B1(n12874), .B2(n13608), .ZN(
        n6073) );
  OAI22_X1 U2289 ( .A1(n12902), .A2(n13243), .B1(n12892), .B2(n13579), .ZN(
        n6102) );
  OAI22_X1 U2290 ( .A1(n12902), .A2(n13246), .B1(n12892), .B2(n13578), .ZN(
        n6103) );
  OAI22_X1 U2291 ( .A1(n12902), .A2(n13249), .B1(n12892), .B2(n13577), .ZN(
        n6104) );
  OAI22_X1 U2292 ( .A1(n12902), .A2(n13252), .B1(n12892), .B2(n13576), .ZN(
        n6105) );
  OAI22_X1 U2293 ( .A1(n12902), .A2(n13255), .B1(n12892), .B2(n13575), .ZN(
        n6106) );
  OAI22_X1 U2294 ( .A1(n12901), .A2(n13258), .B1(n12892), .B2(n13574), .ZN(
        n6107) );
  OAI22_X1 U2295 ( .A1(n12901), .A2(n13261), .B1(n12892), .B2(n13573), .ZN(
        n6108) );
  OAI22_X1 U2296 ( .A1(n12901), .A2(n13264), .B1(n12892), .B2(n13572), .ZN(
        n6109) );
  OAI22_X1 U2297 ( .A1(n12901), .A2(n13267), .B1(n12892), .B2(n13571), .ZN(
        n6110) );
  OAI22_X1 U2298 ( .A1(n12901), .A2(n13270), .B1(n12892), .B2(n13570), .ZN(
        n6111) );
  OAI22_X1 U2299 ( .A1(n12900), .A2(n13273), .B1(n12892), .B2(n13569), .ZN(
        n6112) );
  OAI22_X1 U2300 ( .A1(n12900), .A2(n13276), .B1(n12892), .B2(n13568), .ZN(
        n6113) );
  OAI22_X1 U2301 ( .A1(n12900), .A2(n13279), .B1(n12893), .B2(n13567), .ZN(
        n6114) );
  OAI22_X1 U2302 ( .A1(n12900), .A2(n13282), .B1(n12893), .B2(n13566), .ZN(
        n6115) );
  OAI22_X1 U2303 ( .A1(n12900), .A2(n13285), .B1(n12893), .B2(n13565), .ZN(
        n6116) );
  OAI22_X1 U2304 ( .A1(n12899), .A2(n13288), .B1(n12893), .B2(n13564), .ZN(
        n6117) );
  OAI22_X1 U2305 ( .A1(n12899), .A2(n13291), .B1(n12893), .B2(n13563), .ZN(
        n6118) );
  OAI22_X1 U2306 ( .A1(n12899), .A2(n13294), .B1(n12893), .B2(n13562), .ZN(
        n6119) );
  OAI22_X1 U2307 ( .A1(n12899), .A2(n13297), .B1(n12893), .B2(n13561), .ZN(
        n6120) );
  OAI22_X1 U2308 ( .A1(n12899), .A2(n13300), .B1(n12893), .B2(n13560), .ZN(
        n6121) );
  OAI22_X1 U2309 ( .A1(n12898), .A2(n13303), .B1(n12893), .B2(n13559), .ZN(
        n6122) );
  OAI22_X1 U2310 ( .A1(n12898), .A2(n13306), .B1(n12893), .B2(n13558), .ZN(
        n6123) );
  OAI22_X1 U2311 ( .A1(n12898), .A2(n13309), .B1(n12893), .B2(n13557), .ZN(
        n6124) );
  OAI22_X1 U2312 ( .A1(n12898), .A2(n13312), .B1(n12893), .B2(n13556), .ZN(
        n6125) );
  OAI22_X1 U2313 ( .A1(n12898), .A2(n13315), .B1(n12894), .B2(n13555), .ZN(
        n6126) );
  OAI22_X1 U2314 ( .A1(n12897), .A2(n13318), .B1(n12894), .B2(n13554), .ZN(
        n6127) );
  OAI22_X1 U2315 ( .A1(n12897), .A2(n13321), .B1(n12894), .B2(n13553), .ZN(
        n6128) );
  OAI22_X1 U2316 ( .A1(n12897), .A2(n13324), .B1(n12894), .B2(n13552), .ZN(
        n6129) );
  OAI22_X1 U2317 ( .A1(n12897), .A2(n13327), .B1(n12894), .B2(n13551), .ZN(
        n6130) );
  OAI22_X1 U2318 ( .A1(n12897), .A2(n13330), .B1(n12894), .B2(n13550), .ZN(
        n6131) );
  OAI22_X1 U2319 ( .A1(n12896), .A2(n13333), .B1(n12894), .B2(n13549), .ZN(
        n6132) );
  OAI22_X1 U2320 ( .A1(n12896), .A2(n13336), .B1(n12894), .B2(n13548), .ZN(
        n6133) );
  OAI22_X1 U2321 ( .A1(n12896), .A2(n13339), .B1(n12894), .B2(n13547), .ZN(
        n6134) );
  OAI22_X1 U2322 ( .A1(n12896), .A2(n13342), .B1(n12894), .B2(n13546), .ZN(
        n6135) );
  OAI22_X1 U2323 ( .A1(n12896), .A2(n13345), .B1(n12894), .B2(n13545), .ZN(
        n6136) );
  OAI22_X1 U2324 ( .A1(n12895), .A2(n13348), .B1(n12894), .B2(n13544), .ZN(
        n6137) );
  OAI22_X1 U2325 ( .A1(n12962), .A2(n13242), .B1(n12952), .B2(n13530), .ZN(
        n6294) );
  OAI22_X1 U2326 ( .A1(n12962), .A2(n13245), .B1(n12952), .B2(n13529), .ZN(
        n6295) );
  OAI22_X1 U2327 ( .A1(n12962), .A2(n13248), .B1(n12952), .B2(n13528), .ZN(
        n6296) );
  OAI22_X1 U2328 ( .A1(n12962), .A2(n13251), .B1(n12952), .B2(n13527), .ZN(
        n6297) );
  OAI22_X1 U2329 ( .A1(n12962), .A2(n13254), .B1(n12952), .B2(n13526), .ZN(
        n6298) );
  OAI22_X1 U2330 ( .A1(n12961), .A2(n13257), .B1(n12952), .B2(n13525), .ZN(
        n6299) );
  OAI22_X1 U2331 ( .A1(n12961), .A2(n13260), .B1(n12952), .B2(n13524), .ZN(
        n6300) );
  OAI22_X1 U2332 ( .A1(n12961), .A2(n13263), .B1(n12952), .B2(n13523), .ZN(
        n6301) );
  OAI22_X1 U2333 ( .A1(n12961), .A2(n13266), .B1(n12952), .B2(n13522), .ZN(
        n6302) );
  OAI22_X1 U2334 ( .A1(n12961), .A2(n13269), .B1(n12952), .B2(n13521), .ZN(
        n6303) );
  OAI22_X1 U2335 ( .A1(n12960), .A2(n13272), .B1(n12952), .B2(n13520), .ZN(
        n6304) );
  OAI22_X1 U2336 ( .A1(n12960), .A2(n13275), .B1(n12952), .B2(n13519), .ZN(
        n6305) );
  OAI22_X1 U2337 ( .A1(n12960), .A2(n13278), .B1(n12953), .B2(n13518), .ZN(
        n6306) );
  OAI22_X1 U2338 ( .A1(n12960), .A2(n13281), .B1(n12953), .B2(n13517), .ZN(
        n6307) );
  OAI22_X1 U2339 ( .A1(n12960), .A2(n13284), .B1(n12953), .B2(n13516), .ZN(
        n6308) );
  OAI22_X1 U2340 ( .A1(n12959), .A2(n13299), .B1(n12953), .B2(n13515), .ZN(
        n6313) );
  OAI22_X1 U2341 ( .A1(n12958), .A2(n13302), .B1(n12953), .B2(n13514), .ZN(
        n6314) );
  OAI22_X1 U2342 ( .A1(n12958), .A2(n13305), .B1(n12953), .B2(n13513), .ZN(
        n6315) );
  OAI22_X1 U2343 ( .A1(n12958), .A2(n13308), .B1(n12953), .B2(n13512), .ZN(
        n6316) );
  OAI22_X1 U2344 ( .A1(n12958), .A2(n13311), .B1(n12953), .B2(n13511), .ZN(
        n6317) );
  OAI22_X1 U2345 ( .A1(n12958), .A2(n13314), .B1(n12954), .B2(n13510), .ZN(
        n6318) );
  OAI22_X1 U2346 ( .A1(n12957), .A2(n13317), .B1(n12954), .B2(n13509), .ZN(
        n6319) );
  OAI22_X1 U2347 ( .A1(n12957), .A2(n13320), .B1(n12954), .B2(n13508), .ZN(
        n6320) );
  OAI22_X1 U2348 ( .A1(n12957), .A2(n13323), .B1(n12954), .B2(n13507), .ZN(
        n6321) );
  OAI22_X1 U2349 ( .A1(n12957), .A2(n13326), .B1(n12954), .B2(n13506), .ZN(
        n6322) );
  OAI22_X1 U2350 ( .A1(n12957), .A2(n13329), .B1(n12954), .B2(n13505), .ZN(
        n6323) );
  OAI22_X1 U2351 ( .A1(n12956), .A2(n13332), .B1(n12954), .B2(n13504), .ZN(
        n6324) );
  OAI22_X1 U2352 ( .A1(n12956), .A2(n13335), .B1(n12954), .B2(n13503), .ZN(
        n6325) );
  OAI22_X1 U2353 ( .A1(n12956), .A2(n13338), .B1(n12954), .B2(n13502), .ZN(
        n6326) );
  OAI22_X1 U2354 ( .A1(n12956), .A2(n13341), .B1(n12954), .B2(n13501), .ZN(
        n6327) );
  OAI22_X1 U2355 ( .A1(n12956), .A2(n13344), .B1(n12954), .B2(n13500), .ZN(
        n6328) );
  OAI22_X1 U2356 ( .A1(n12955), .A2(n13347), .B1(n12954), .B2(n13499), .ZN(
        n6329) );
  OAI22_X1 U2357 ( .A1(n12982), .A2(n13242), .B1(n12972), .B2(n13470), .ZN(
        n6358) );
  OAI22_X1 U2358 ( .A1(n12982), .A2(n13245), .B1(n12972), .B2(n13469), .ZN(
        n6359) );
  OAI22_X1 U2359 ( .A1(n12982), .A2(n13248), .B1(n12972), .B2(n13468), .ZN(
        n6360) );
  OAI22_X1 U2360 ( .A1(n12982), .A2(n13251), .B1(n12972), .B2(n13467), .ZN(
        n6361) );
  OAI22_X1 U2361 ( .A1(n12982), .A2(n13254), .B1(n12972), .B2(n13466), .ZN(
        n6362) );
  OAI22_X1 U2362 ( .A1(n12981), .A2(n13257), .B1(n12972), .B2(n13465), .ZN(
        n6363) );
  OAI22_X1 U2363 ( .A1(n12981), .A2(n13260), .B1(n12972), .B2(n13464), .ZN(
        n6364) );
  OAI22_X1 U2364 ( .A1(n12981), .A2(n13263), .B1(n12972), .B2(n13463), .ZN(
        n6365) );
  OAI22_X1 U2365 ( .A1(n12981), .A2(n13266), .B1(n12972), .B2(n13462), .ZN(
        n6366) );
  OAI22_X1 U2366 ( .A1(n12981), .A2(n13269), .B1(n12972), .B2(n13461), .ZN(
        n6367) );
  OAI22_X1 U2367 ( .A1(n12980), .A2(n13272), .B1(n12972), .B2(n13460), .ZN(
        n6368) );
  OAI22_X1 U2368 ( .A1(n12980), .A2(n13275), .B1(n12972), .B2(n13459), .ZN(
        n6369) );
  OAI22_X1 U2369 ( .A1(n12980), .A2(n13278), .B1(n12973), .B2(n13458), .ZN(
        n6370) );
  OAI22_X1 U2370 ( .A1(n12980), .A2(n13281), .B1(n12973), .B2(n13457), .ZN(
        n6371) );
  OAI22_X1 U2371 ( .A1(n12980), .A2(n13284), .B1(n12973), .B2(n13456), .ZN(
        n6372) );
  OAI22_X1 U2372 ( .A1(n12979), .A2(n13287), .B1(n12973), .B2(n13455), .ZN(
        n6373) );
  OAI22_X1 U2373 ( .A1(n12979), .A2(n13290), .B1(n12973), .B2(n13454), .ZN(
        n6374) );
  OAI22_X1 U2374 ( .A1(n12979), .A2(n13293), .B1(n12973), .B2(n13453), .ZN(
        n6375) );
  OAI22_X1 U2375 ( .A1(n12979), .A2(n13296), .B1(n12973), .B2(n13452), .ZN(
        n6376) );
  OAI22_X1 U2376 ( .A1(n12979), .A2(n13299), .B1(n12973), .B2(n13451), .ZN(
        n6377) );
  OAI22_X1 U2377 ( .A1(n12978), .A2(n13302), .B1(n12973), .B2(n13450), .ZN(
        n6378) );
  OAI22_X1 U2378 ( .A1(n12978), .A2(n13305), .B1(n12973), .B2(n13449), .ZN(
        n6379) );
  OAI22_X1 U2379 ( .A1(n12978), .A2(n13308), .B1(n12973), .B2(n13448), .ZN(
        n6380) );
  OAI22_X1 U2380 ( .A1(n12978), .A2(n13311), .B1(n12973), .B2(n13447), .ZN(
        n6381) );
  OAI22_X1 U2381 ( .A1(n12978), .A2(n13314), .B1(n12974), .B2(n13446), .ZN(
        n6382) );
  OAI22_X1 U2382 ( .A1(n12977), .A2(n13317), .B1(n12974), .B2(n13445), .ZN(
        n6383) );
  OAI22_X1 U2383 ( .A1(n12977), .A2(n13320), .B1(n12974), .B2(n13444), .ZN(
        n6384) );
  OAI22_X1 U2384 ( .A1(n12977), .A2(n13323), .B1(n12974), .B2(n13443), .ZN(
        n6385) );
  OAI22_X1 U2385 ( .A1(n12977), .A2(n13326), .B1(n12974), .B2(n13442), .ZN(
        n6386) );
  OAI22_X1 U2386 ( .A1(n12977), .A2(n13329), .B1(n12974), .B2(n13441), .ZN(
        n6387) );
  OAI22_X1 U2387 ( .A1(n12976), .A2(n13332), .B1(n12974), .B2(n13440), .ZN(
        n6388) );
  OAI22_X1 U2388 ( .A1(n12976), .A2(n13335), .B1(n12974), .B2(n13439), .ZN(
        n6389) );
  OAI22_X1 U2389 ( .A1(n12976), .A2(n13338), .B1(n12974), .B2(n13438), .ZN(
        n6390) );
  OAI22_X1 U2390 ( .A1(n12976), .A2(n13341), .B1(n12974), .B2(n13437), .ZN(
        n6391) );
  OAI22_X1 U2391 ( .A1(n12976), .A2(n13344), .B1(n12974), .B2(n13436), .ZN(
        n6392) );
  OAI22_X1 U2392 ( .A1(n12975), .A2(n13347), .B1(n12974), .B2(n13435), .ZN(
        n6393) );
  OAI22_X1 U2393 ( .A1(n13162), .A2(n13242), .B1(n13152), .B2(n13406), .ZN(
        n6934) );
  OAI22_X1 U2394 ( .A1(n13162), .A2(n13245), .B1(n13152), .B2(n13405), .ZN(
        n6935) );
  OAI22_X1 U2395 ( .A1(n13162), .A2(n13248), .B1(n13152), .B2(n13404), .ZN(
        n6936) );
  OAI22_X1 U2396 ( .A1(n13162), .A2(n13251), .B1(n13152), .B2(n13403), .ZN(
        n6937) );
  OAI22_X1 U2397 ( .A1(n13162), .A2(n13254), .B1(n13152), .B2(n13402), .ZN(
        n6938) );
  OAI22_X1 U2398 ( .A1(n13367), .A2(n13308), .B1(n13362), .B2(n13401), .ZN(
        n7020) );
  OAI22_X1 U2399 ( .A1(n13367), .A2(n13311), .B1(n13362), .B2(n13400), .ZN(
        n7021) );
  OAI22_X1 U2400 ( .A1(n13367), .A2(n13314), .B1(n13363), .B2(n13399), .ZN(
        n7022) );
  OAI22_X1 U2401 ( .A1(n13366), .A2(n13317), .B1(n13363), .B2(n13398), .ZN(
        n7023) );
  OAI22_X1 U2402 ( .A1(n13366), .A2(n13320), .B1(n13363), .B2(n13397), .ZN(
        n7024) );
  OAI22_X1 U2403 ( .A1(n13366), .A2(n13323), .B1(n13363), .B2(n13396), .ZN(
        n7025) );
  OAI22_X1 U2404 ( .A1(n13366), .A2(n13326), .B1(n13363), .B2(n13395), .ZN(
        n7026) );
  OAI22_X1 U2405 ( .A1(n13366), .A2(n13329), .B1(n13363), .B2(n13394), .ZN(
        n7027) );
  OAI22_X1 U2406 ( .A1(n13365), .A2(n13332), .B1(n13363), .B2(n13393), .ZN(
        n7028) );
  OAI22_X1 U2407 ( .A1(n13364), .A2(n13350), .B1(n13361), .B2(n14435), .ZN(
        n7034) );
  OAI22_X1 U2408 ( .A1(n13364), .A2(n13353), .B1(n13362), .B2(n14434), .ZN(
        n7035) );
  OAI22_X1 U2409 ( .A1(n13364), .A2(n13356), .B1(n13363), .B2(n14433), .ZN(
        n7036) );
  OAI22_X1 U2410 ( .A1(n13155), .A2(n13350), .B1(n13154), .B2(n14412), .ZN(
        n6970) );
  OAI22_X1 U2411 ( .A1(n13155), .A2(n13353), .B1(n13153), .B2(n14411), .ZN(
        n6971) );
  OAI22_X1 U2412 ( .A1(n13155), .A2(n13356), .B1(n13152), .B2(n14410), .ZN(
        n6972) );
  OAI22_X1 U2413 ( .A1(n13155), .A2(n13379), .B1(n13154), .B2(n14409), .ZN(
        n6973) );
  OAI22_X1 U2414 ( .A1(n12600), .A2(n13352), .B1(n12599), .B2(n14086), .ZN(
        n5178) );
  OAI22_X1 U2415 ( .A1(n12600), .A2(n13355), .B1(n12597), .B2(n14085), .ZN(
        n5179) );
  OAI22_X1 U2416 ( .A1(n12600), .A2(n13358), .B1(n12598), .B2(n14084), .ZN(
        n5180) );
  OAI22_X1 U2417 ( .A1(n12600), .A2(n13381), .B1(n12599), .B2(n14083), .ZN(
        n5181) );
  OAI22_X1 U2418 ( .A1(n13095), .A2(n13350), .B1(n13092), .B2(n13847), .ZN(
        n6778) );
  OAI22_X1 U2419 ( .A1(n13095), .A2(n13353), .B1(n13093), .B2(n13846), .ZN(
        n6779) );
  OAI22_X1 U2420 ( .A1(n13095), .A2(n13356), .B1(n13094), .B2(n13845), .ZN(
        n6780) );
  OAI22_X1 U2421 ( .A1(n13095), .A2(n13379), .B1(n13092), .B2(n13844), .ZN(
        n6781) );
  OAI22_X1 U2422 ( .A1(n13075), .A2(n13350), .B1(n13072), .B2(n13843), .ZN(
        n6714) );
  OAI22_X1 U2423 ( .A1(n13075), .A2(n13353), .B1(n13073), .B2(n13842), .ZN(
        n6715) );
  OAI22_X1 U2424 ( .A1(n13075), .A2(n13356), .B1(n13074), .B2(n13841), .ZN(
        n6716) );
  OAI22_X1 U2425 ( .A1(n13075), .A2(n13379), .B1(n13072), .B2(n13840), .ZN(
        n6717) );
  OAI22_X1 U2426 ( .A1(n12619), .A2(n13352), .B1(n12616), .B2(n13750), .ZN(
        n5242) );
  OAI22_X1 U2427 ( .A1(n12619), .A2(n13355), .B1(n12617), .B2(n13749), .ZN(
        n5243) );
  OAI22_X1 U2428 ( .A1(n12619), .A2(n13358), .B1(n12618), .B2(n13748), .ZN(
        n5244) );
  OAI22_X1 U2429 ( .A1(n12619), .A2(n13381), .B1(n12616), .B2(n13747), .ZN(
        n5245) );
  OAI22_X1 U2430 ( .A1(n12676), .A2(n13352), .B1(n12674), .B2(n13734), .ZN(
        n5434) );
  OAI22_X1 U2431 ( .A1(n12676), .A2(n13355), .B1(n12673), .B2(n13733), .ZN(
        n5435) );
  OAI22_X1 U2432 ( .A1(n12676), .A2(n13358), .B1(n12675), .B2(n13732), .ZN(
        n5436) );
  OAI22_X1 U2433 ( .A1(n12676), .A2(n13381), .B1(n12674), .B2(n13731), .ZN(
        n5437) );
  OAI22_X1 U2434 ( .A1(n12695), .A2(n13352), .B1(n12692), .B2(n13670), .ZN(
        n5498) );
  OAI22_X1 U2435 ( .A1(n12695), .A2(n13355), .B1(n12693), .B2(n13669), .ZN(
        n5499) );
  OAI22_X1 U2436 ( .A1(n12695), .A2(n13358), .B1(n12694), .B2(n13668), .ZN(
        n5500) );
  OAI22_X1 U2437 ( .A1(n12695), .A2(n13381), .B1(n12692), .B2(n13667), .ZN(
        n5501) );
  OAI22_X1 U2438 ( .A1(n12875), .A2(n13351), .B1(n12872), .B2(n13607), .ZN(
        n6074) );
  OAI22_X1 U2439 ( .A1(n12875), .A2(n13354), .B1(n12873), .B2(n13606), .ZN(
        n6075) );
  OAI22_X1 U2440 ( .A1(n12875), .A2(n13357), .B1(n12874), .B2(n13605), .ZN(
        n6076) );
  OAI22_X1 U2441 ( .A1(n12875), .A2(n13380), .B1(n12872), .B2(n13604), .ZN(
        n6077) );
  OAI22_X1 U2442 ( .A1(n12895), .A2(n13351), .B1(n12892), .B2(n13543), .ZN(
        n6138) );
  OAI22_X1 U2443 ( .A1(n12895), .A2(n13354), .B1(n12893), .B2(n13542), .ZN(
        n6139) );
  OAI22_X1 U2444 ( .A1(n12895), .A2(n13357), .B1(n12894), .B2(n13541), .ZN(
        n6140) );
  OAI22_X1 U2445 ( .A1(n12895), .A2(n13380), .B1(n12892), .B2(n13540), .ZN(
        n6141) );
  OAI22_X1 U2446 ( .A1(n12955), .A2(n13350), .B1(n12952), .B2(n13498), .ZN(
        n6330) );
  OAI22_X1 U2447 ( .A1(n12955), .A2(n13353), .B1(n12953), .B2(n13497), .ZN(
        n6331) );
  OAI22_X1 U2448 ( .A1(n12955), .A2(n13356), .B1(n12954), .B2(n13496), .ZN(
        n6332) );
  OAI22_X1 U2449 ( .A1(n12955), .A2(n13379), .B1(n12952), .B2(n13495), .ZN(
        n6333) );
  OAI22_X1 U2450 ( .A1(n12975), .A2(n13350), .B1(n12972), .B2(n13434), .ZN(
        n6394) );
  OAI22_X1 U2451 ( .A1(n12975), .A2(n13353), .B1(n12973), .B2(n13433), .ZN(
        n6395) );
  OAI22_X1 U2452 ( .A1(n12975), .A2(n13356), .B1(n12974), .B2(n13432), .ZN(
        n6396) );
  OAI22_X1 U2453 ( .A1(n12975), .A2(n13379), .B1(n12972), .B2(n13431), .ZN(
        n6397) );
  OAI22_X1 U2454 ( .A1(n13364), .A2(n13379), .B1(n13361), .B2(n13392), .ZN(
        n7037) );
  INV_X1 U2455 ( .A(ADD_RD1[3]), .ZN(n14462) );
  INV_X1 U2456 ( .A(ADD_RD1[4]), .ZN(n14461) );
  INV_X1 U2457 ( .A(ADD_RD1[0]), .ZN(n14465) );
  INV_X1 U2458 ( .A(ADD_RD1[1]), .ZN(n14464) );
  INV_X1 U2459 ( .A(ADD_RD1[2]), .ZN(n14463) );
  INV_X1 U2460 ( .A(ADD_WR[2]), .ZN(n13384) );
  INV_X1 U2461 ( .A(ADD_WR[0]), .ZN(n13386) );
  INV_X1 U2462 ( .A(ADD_WR[1]), .ZN(n13385) );
  INV_X1 U2463 ( .A(ADD_WR[3]), .ZN(n13383) );
  NOR2_X1 U2464 ( .A1(n13389), .A2(n13390), .ZN(n4455) );
  NOR3_X1 U2465 ( .A1(n13391), .A2(n13387), .A3(n13388), .ZN(n4470) );
  AOI221_X1 U2466 ( .B1(n12302), .B2(n11586), .C1(n12296), .C2(n11406), .A(
        n4453), .ZN(n4446) );
  OAI22_X1 U2467 ( .A1(n14362), .A2(n12290), .B1(n14361), .B2(n12284), .ZN(
        n4453) );
  AOI221_X1 U2468 ( .B1(n12302), .B2(n11587), .C1(n12296), .C2(n11407), .A(
        n4411), .ZN(n4408) );
  OAI22_X1 U2469 ( .A1(n14407), .A2(n12290), .B1(n14384), .B2(n12284), .ZN(
        n4411) );
  AOI221_X1 U2470 ( .B1(n12302), .B2(n11588), .C1(n12296), .C2(n11408), .A(
        n4392), .ZN(n4389) );
  OAI22_X1 U2471 ( .A1(n14406), .A2(n12290), .B1(n14383), .B2(n12284), .ZN(
        n4392) );
  AOI221_X1 U2472 ( .B1(n12302), .B2(n11589), .C1(n12296), .C2(n11409), .A(
        n4373), .ZN(n4370) );
  OAI22_X1 U2473 ( .A1(n14405), .A2(n12290), .B1(n14382), .B2(n12284), .ZN(
        n4373) );
  AOI221_X1 U2474 ( .B1(n12302), .B2(n11590), .C1(n12296), .C2(n11410), .A(
        n4316), .ZN(n4313) );
  OAI22_X1 U2475 ( .A1(n14402), .A2(n12290), .B1(n14379), .B2(n12284), .ZN(
        n4316) );
  AOI221_X1 U2476 ( .B1(n12302), .B2(n11591), .C1(n12296), .C2(n11411), .A(
        n4297), .ZN(n4294) );
  OAI22_X1 U2477 ( .A1(n14401), .A2(n12290), .B1(n14378), .B2(n12284), .ZN(
        n4297) );
  AOI221_X1 U2478 ( .B1(n12302), .B2(n11592), .C1(n12296), .C2(n11412), .A(
        n4278), .ZN(n4275) );
  OAI22_X1 U2479 ( .A1(n14400), .A2(n12290), .B1(n14377), .B2(n12284), .ZN(
        n4278) );
  AOI221_X1 U2480 ( .B1(n12302), .B2(n11593), .C1(n12296), .C2(n11413), .A(
        n4259), .ZN(n4256) );
  OAI22_X1 U2481 ( .A1(n14399), .A2(n12290), .B1(n14376), .B2(n12284), .ZN(
        n4259) );
  AOI221_X1 U2482 ( .B1(n12302), .B2(n11594), .C1(n12296), .C2(n11414), .A(
        n4240), .ZN(n4237) );
  OAI22_X1 U2483 ( .A1(n14398), .A2(n12290), .B1(n14375), .B2(n12284), .ZN(
        n4240) );
  AOI221_X1 U2484 ( .B1(n12303), .B2(n11595), .C1(n12297), .C2(n11415), .A(
        n4221), .ZN(n4218) );
  OAI22_X1 U2485 ( .A1(n14397), .A2(n12291), .B1(n14374), .B2(n12285), .ZN(
        n4221) );
  AOI221_X1 U2486 ( .B1(n12303), .B2(n11596), .C1(n12297), .C2(n11416), .A(
        n4202), .ZN(n4199) );
  OAI22_X1 U2487 ( .A1(n14396), .A2(n12291), .B1(n14373), .B2(n12285), .ZN(
        n4202) );
  AOI221_X1 U2488 ( .B1(n12303), .B2(n11597), .C1(n12297), .C2(n11417), .A(
        n4183), .ZN(n4180) );
  OAI22_X1 U2489 ( .A1(n14395), .A2(n12291), .B1(n14372), .B2(n12285), .ZN(
        n4183) );
  AOI221_X1 U2490 ( .B1(n12303), .B2(n11598), .C1(n12297), .C2(n11418), .A(
        n4164), .ZN(n4161) );
  OAI22_X1 U2491 ( .A1(n14394), .A2(n12291), .B1(n14371), .B2(n12285), .ZN(
        n4164) );
  AOI221_X1 U2492 ( .B1(n12303), .B2(n11599), .C1(n12297), .C2(n11419), .A(
        n4145), .ZN(n4142) );
  OAI22_X1 U2493 ( .A1(n14393), .A2(n12291), .B1(n14370), .B2(n12285), .ZN(
        n4145) );
  AOI221_X1 U2494 ( .B1(n12303), .B2(n11600), .C1(n12297), .C2(n11420), .A(
        n4126), .ZN(n4123) );
  OAI22_X1 U2495 ( .A1(n14392), .A2(n12291), .B1(n14369), .B2(n12285), .ZN(
        n4126) );
  AOI221_X1 U2496 ( .B1(n12303), .B2(n11601), .C1(n12297), .C2(n11421), .A(
        n4107), .ZN(n4104) );
  OAI22_X1 U2497 ( .A1(n14391), .A2(n12291), .B1(n14368), .B2(n12285), .ZN(
        n4107) );
  AOI221_X1 U2498 ( .B1(n12303), .B2(n11602), .C1(n12297), .C2(n11422), .A(
        n4088), .ZN(n4085) );
  OAI22_X1 U2499 ( .A1(n14390), .A2(n12291), .B1(n14367), .B2(n12285), .ZN(
        n4088) );
  AOI221_X1 U2500 ( .B1(n12303), .B2(n11603), .C1(n12297), .C2(n11423), .A(
        n4069), .ZN(n4066) );
  OAI22_X1 U2501 ( .A1(n14389), .A2(n12291), .B1(n14366), .B2(n12285), .ZN(
        n4069) );
  AOI221_X1 U2502 ( .B1(n12303), .B2(n11604), .C1(n12297), .C2(n11424), .A(
        n4050), .ZN(n4047) );
  OAI22_X1 U2503 ( .A1(n14388), .A2(n12291), .B1(n14365), .B2(n12285), .ZN(
        n4050) );
  AOI221_X1 U2504 ( .B1(n12303), .B2(n11605), .C1(n12297), .C2(n11425), .A(
        n4031), .ZN(n4028) );
  OAI22_X1 U2505 ( .A1(n14387), .A2(n12291), .B1(n14364), .B2(n12285), .ZN(
        n4031) );
  AOI221_X1 U2506 ( .B1(n12303), .B2(n11606), .C1(n12297), .C2(n11426), .A(
        n4012), .ZN(n4009) );
  OAI22_X1 U2507 ( .A1(n14386), .A2(n12291), .B1(n14363), .B2(n12285), .ZN(
        n4012) );
  AOI221_X1 U2508 ( .B1(n12304), .B2(n11607), .C1(n12298), .C2(n11427), .A(
        n3993), .ZN(n3990) );
  OAI22_X1 U2509 ( .A1(n14288), .A2(n12292), .B1(n14252), .B2(n12286), .ZN(
        n3993) );
  AOI221_X1 U2510 ( .B1(n12304), .B2(n11608), .C1(n12298), .C2(n11428), .A(
        n3974), .ZN(n3971) );
  OAI22_X1 U2511 ( .A1(n14287), .A2(n12292), .B1(n14251), .B2(n12286), .ZN(
        n3974) );
  AOI221_X1 U2512 ( .B1(n12304), .B2(n11609), .C1(n12298), .C2(n11429), .A(
        n3955), .ZN(n3952) );
  OAI22_X1 U2513 ( .A1(n14286), .A2(n12292), .B1(n14250), .B2(n12286), .ZN(
        n3955) );
  AOI221_X1 U2514 ( .B1(n12304), .B2(n11610), .C1(n12298), .C2(n11430), .A(
        n3936), .ZN(n3933) );
  OAI22_X1 U2515 ( .A1(n14285), .A2(n12292), .B1(n14249), .B2(n12286), .ZN(
        n3936) );
  AOI221_X1 U2516 ( .B1(n12304), .B2(n11611), .C1(n12298), .C2(n11431), .A(
        n3917), .ZN(n3914) );
  OAI22_X1 U2517 ( .A1(n14284), .A2(n12292), .B1(n14248), .B2(n12286), .ZN(
        n3917) );
  AOI221_X1 U2518 ( .B1(n12304), .B2(n11612), .C1(n12298), .C2(n11432), .A(
        n3898), .ZN(n3895) );
  OAI22_X1 U2519 ( .A1(n14283), .A2(n12292), .B1(n14247), .B2(n12286), .ZN(
        n3898) );
  AOI221_X1 U2520 ( .B1(n12304), .B2(n11613), .C1(n12298), .C2(n11433), .A(
        n3879), .ZN(n3876) );
  OAI22_X1 U2521 ( .A1(n14282), .A2(n12292), .B1(n14246), .B2(n12286), .ZN(
        n3879) );
  AOI221_X1 U2522 ( .B1(n12304), .B2(n11614), .C1(n12298), .C2(n11434), .A(
        n3860), .ZN(n3857) );
  OAI22_X1 U2523 ( .A1(n14281), .A2(n12292), .B1(n14245), .B2(n12286), .ZN(
        n3860) );
  AOI221_X1 U2524 ( .B1(n12304), .B2(n11615), .C1(n12298), .C2(n11435), .A(
        n3841), .ZN(n3838) );
  OAI22_X1 U2525 ( .A1(n14280), .A2(n12292), .B1(n14244), .B2(n12286), .ZN(
        n3841) );
  AOI221_X1 U2526 ( .B1(n12304), .B2(n11616), .C1(n12298), .C2(n11436), .A(
        n3822), .ZN(n3819) );
  OAI22_X1 U2527 ( .A1(n14279), .A2(n12292), .B1(n14243), .B2(n12286), .ZN(
        n3822) );
  AOI221_X1 U2528 ( .B1(n12304), .B2(n11617), .C1(n12298), .C2(n11437), .A(
        n3803), .ZN(n3800) );
  OAI22_X1 U2529 ( .A1(n14278), .A2(n12292), .B1(n14242), .B2(n12286), .ZN(
        n3803) );
  AOI221_X1 U2530 ( .B1(n12304), .B2(n11618), .C1(n12298), .C2(n11438), .A(
        n3784), .ZN(n3781) );
  OAI22_X1 U2531 ( .A1(n14277), .A2(n12292), .B1(n14241), .B2(n12286), .ZN(
        n3784) );
  AOI221_X1 U2532 ( .B1(n12305), .B2(n11619), .C1(n12299), .C2(n11439), .A(
        n3765), .ZN(n3762) );
  OAI22_X1 U2533 ( .A1(n14276), .A2(n12293), .B1(n14240), .B2(n12287), .ZN(
        n3765) );
  AOI221_X1 U2534 ( .B1(n12305), .B2(n11620), .C1(n12299), .C2(n11440), .A(
        n3746), .ZN(n3743) );
  OAI22_X1 U2535 ( .A1(n14275), .A2(n12293), .B1(n14239), .B2(n12287), .ZN(
        n3746) );
  AOI221_X1 U2536 ( .B1(n12305), .B2(n11621), .C1(n12299), .C2(n11441), .A(
        n3727), .ZN(n3724) );
  OAI22_X1 U2537 ( .A1(n14274), .A2(n12293), .B1(n14238), .B2(n12287), .ZN(
        n3727) );
  AOI221_X1 U2538 ( .B1(n12305), .B2(n11622), .C1(n12299), .C2(n11442), .A(
        n3708), .ZN(n3705) );
  OAI22_X1 U2539 ( .A1(n14273), .A2(n12293), .B1(n14237), .B2(n12287), .ZN(
        n3708) );
  AOI221_X1 U2540 ( .B1(n12305), .B2(n11623), .C1(n12299), .C2(n11443), .A(
        n3689), .ZN(n3686) );
  OAI22_X1 U2541 ( .A1(n14272), .A2(n12293), .B1(n14236), .B2(n12287), .ZN(
        n3689) );
  AOI221_X1 U2542 ( .B1(n12305), .B2(n11624), .C1(n12299), .C2(n11444), .A(
        n3670), .ZN(n3667) );
  OAI22_X1 U2543 ( .A1(n14271), .A2(n12293), .B1(n14235), .B2(n12287), .ZN(
        n3670) );
  AOI221_X1 U2544 ( .B1(n12305), .B2(n11625), .C1(n12299), .C2(n11445), .A(
        n3651), .ZN(n3648) );
  OAI22_X1 U2545 ( .A1(n14270), .A2(n12293), .B1(n14234), .B2(n12287), .ZN(
        n3651) );
  AOI221_X1 U2546 ( .B1(n12305), .B2(n11626), .C1(n12299), .C2(n11446), .A(
        n3632), .ZN(n3629) );
  OAI22_X1 U2547 ( .A1(n14269), .A2(n12293), .B1(n14233), .B2(n12287), .ZN(
        n3632) );
  AOI221_X1 U2548 ( .B1(n12305), .B2(n11627), .C1(n12299), .C2(n11447), .A(
        n3613), .ZN(n3610) );
  OAI22_X1 U2549 ( .A1(n14268), .A2(n12293), .B1(n14232), .B2(n12287), .ZN(
        n3613) );
  AOI221_X1 U2550 ( .B1(n12305), .B2(n11628), .C1(n12299), .C2(n11448), .A(
        n3594), .ZN(n3591) );
  OAI22_X1 U2551 ( .A1(n14267), .A2(n12293), .B1(n14231), .B2(n12287), .ZN(
        n3594) );
  AOI221_X1 U2552 ( .B1(n12305), .B2(n11629), .C1(n12299), .C2(n11449), .A(
        n3575), .ZN(n3572) );
  OAI22_X1 U2553 ( .A1(n14266), .A2(n12293), .B1(n14230), .B2(n12287), .ZN(
        n3575) );
  AOI221_X1 U2554 ( .B1(n12305), .B2(n11630), .C1(n12299), .C2(n11450), .A(
        n3556), .ZN(n3553) );
  OAI22_X1 U2555 ( .A1(n14265), .A2(n12293), .B1(n14229), .B2(n12287), .ZN(
        n3556) );
  AOI221_X1 U2556 ( .B1(n12306), .B2(n11631), .C1(n12300), .C2(n11451), .A(
        n3537), .ZN(n3534) );
  OAI22_X1 U2557 ( .A1(n14264), .A2(n12294), .B1(n14228), .B2(n12288), .ZN(
        n3537) );
  AOI221_X1 U2558 ( .B1(n12306), .B2(n11632), .C1(n12300), .C2(n11452), .A(
        n3518), .ZN(n3515) );
  OAI22_X1 U2559 ( .A1(n14263), .A2(n12294), .B1(n14227), .B2(n12288), .ZN(
        n3518) );
  AOI221_X1 U2560 ( .B1(n12306), .B2(n11633), .C1(n12300), .C2(n11453), .A(
        n3499), .ZN(n3496) );
  OAI22_X1 U2561 ( .A1(n14262), .A2(n12294), .B1(n14226), .B2(n12288), .ZN(
        n3499) );
  AOI221_X1 U2562 ( .B1(n12306), .B2(n11634), .C1(n12300), .C2(n11454), .A(
        n3480), .ZN(n3477) );
  OAI22_X1 U2563 ( .A1(n14261), .A2(n12294), .B1(n14225), .B2(n12288), .ZN(
        n3480) );
  AOI221_X1 U2564 ( .B1(n12306), .B2(n11635), .C1(n12300), .C2(n11455), .A(
        n3461), .ZN(n3458) );
  OAI22_X1 U2565 ( .A1(n14260), .A2(n12294), .B1(n14224), .B2(n12288), .ZN(
        n3461) );
  AOI221_X1 U2566 ( .B1(n12306), .B2(n11636), .C1(n12300), .C2(n11456), .A(
        n3442), .ZN(n3439) );
  OAI22_X1 U2567 ( .A1(n14259), .A2(n12294), .B1(n14223), .B2(n12288), .ZN(
        n3442) );
  AOI221_X1 U2568 ( .B1(n12306), .B2(n11637), .C1(n12300), .C2(n11457), .A(
        n3423), .ZN(n3420) );
  OAI22_X1 U2569 ( .A1(n14258), .A2(n12294), .B1(n14222), .B2(n12288), .ZN(
        n3423) );
  AOI221_X1 U2570 ( .B1(n12306), .B2(n11638), .C1(n12300), .C2(n11458), .A(
        n3404), .ZN(n3401) );
  OAI22_X1 U2571 ( .A1(n14257), .A2(n12294), .B1(n14221), .B2(n12288), .ZN(
        n3404) );
  AOI221_X1 U2572 ( .B1(n12306), .B2(n11639), .C1(n12300), .C2(n11459), .A(
        n3385), .ZN(n3382) );
  OAI22_X1 U2573 ( .A1(n14256), .A2(n12294), .B1(n14220), .B2(n12288), .ZN(
        n3385) );
  AOI221_X1 U2574 ( .B1(n12306), .B2(n11640), .C1(n12300), .C2(n11460), .A(
        n3366), .ZN(n3363) );
  OAI22_X1 U2575 ( .A1(n14255), .A2(n12294), .B1(n14219), .B2(n12288), .ZN(
        n3366) );
  AOI221_X1 U2576 ( .B1(n12306), .B2(n11641), .C1(n12300), .C2(n11461), .A(
        n3347), .ZN(n3344) );
  OAI22_X1 U2577 ( .A1(n14254), .A2(n12294), .B1(n14218), .B2(n12288), .ZN(
        n3347) );
  AOI221_X1 U2578 ( .B1(n12307), .B2(n13835), .C1(n12301), .C2(n13839), .A(
        n3309), .ZN(n3306) );
  OAI22_X1 U2579 ( .A1(n13847), .A2(n12295), .B1(n13843), .B2(n12289), .ZN(
        n3309) );
  AOI221_X1 U2580 ( .B1(n12307), .B2(n13834), .C1(n12301), .C2(n13838), .A(
        n3290), .ZN(n3287) );
  OAI22_X1 U2581 ( .A1(n13846), .A2(n12295), .B1(n13842), .B2(n12289), .ZN(
        n3290) );
  AOI221_X1 U2582 ( .B1(n12307), .B2(n13833), .C1(n12301), .C2(n13837), .A(
        n3271), .ZN(n3268) );
  OAI22_X1 U2583 ( .A1(n13845), .A2(n12295), .B1(n13841), .B2(n12289), .ZN(
        n3271) );
  AOI221_X1 U2584 ( .B1(n12307), .B2(n13832), .C1(n12301), .C2(n13836), .A(
        n3226), .ZN(n3217) );
  OAI22_X1 U2585 ( .A1(n13844), .A2(n12295), .B1(n13840), .B2(n12289), .ZN(
        n3226) );
  AOI221_X1 U2586 ( .B1(n12278), .B2(n11642), .C1(n12272), .C2(n11462), .A(
        n4456), .ZN(n4445) );
  OAI22_X1 U2587 ( .A1(n13539), .A2(n12266), .B1(n13494), .B2(n12260), .ZN(
        n4456) );
  AOI221_X1 U2588 ( .B1(n12182), .B2(n14153), .C1(n12176), .C2(n14154), .A(
        n4468), .ZN(n4461) );
  OAI22_X1 U2589 ( .A1(n13746), .A2(n12170), .B1(n13730), .B2(n12164), .ZN(
        n4468) );
  AOI221_X1 U2590 ( .B1(n12278), .B2(n11643), .C1(n12272), .C2(n11463), .A(
        n4431), .ZN(n4426) );
  OAI22_X1 U2591 ( .A1(n13538), .A2(n12266), .B1(n13493), .B2(n12260), .ZN(
        n4431) );
  AOI221_X1 U2592 ( .B1(n12182), .B2(n14082), .C1(n12176), .C2(n14129), .A(
        n4439), .ZN(n4434) );
  OAI22_X1 U2593 ( .A1(n13745), .A2(n12170), .B1(n13729), .B2(n12164), .ZN(
        n4439) );
  AOI221_X1 U2594 ( .B1(n12278), .B2(n11644), .C1(n12272), .C2(n11464), .A(
        n4412), .ZN(n4407) );
  OAI22_X1 U2595 ( .A1(n13537), .A2(n12266), .B1(n13492), .B2(n12260), .ZN(
        n4412) );
  AOI221_X1 U2596 ( .B1(n12182), .B2(n14081), .C1(n12176), .C2(n14128), .A(
        n4420), .ZN(n4415) );
  OAI22_X1 U2597 ( .A1(n13744), .A2(n12170), .B1(n13728), .B2(n12164), .ZN(
        n4420) );
  AOI221_X1 U2598 ( .B1(n12278), .B2(n11645), .C1(n12272), .C2(n11465), .A(
        n4393), .ZN(n4388) );
  OAI22_X1 U2599 ( .A1(n13536), .A2(n12266), .B1(n13491), .B2(n12260), .ZN(
        n4393) );
  AOI221_X1 U2600 ( .B1(n12182), .B2(n14079), .C1(n12176), .C2(n14126), .A(
        n4401), .ZN(n4396) );
  OAI22_X1 U2601 ( .A1(n13743), .A2(n12170), .B1(n13727), .B2(n12164), .ZN(
        n4401) );
  AOI221_X1 U2602 ( .B1(n12278), .B2(n11646), .C1(n12272), .C2(n11466), .A(
        n4374), .ZN(n4369) );
  OAI22_X1 U2603 ( .A1(n14360), .A2(n12266), .B1(n13490), .B2(n12260), .ZN(
        n4374) );
  AOI221_X1 U2604 ( .B1(n12182), .B2(n14080), .C1(n12176), .C2(n14127), .A(
        n4382), .ZN(n4377) );
  OAI22_X1 U2605 ( .A1(n13892), .A2(n12170), .B1(n13726), .B2(n12164), .ZN(
        n4382) );
  AOI221_X1 U2606 ( .B1(n12278), .B2(n11647), .C1(n12272), .C2(n11467), .A(
        n4355), .ZN(n4350) );
  OAI22_X1 U2607 ( .A1(n14359), .A2(n12266), .B1(n13489), .B2(n12260), .ZN(
        n4355) );
  AOI221_X1 U2608 ( .B1(n12182), .B2(n14078), .C1(n12176), .C2(n14125), .A(
        n4363), .ZN(n4358) );
  OAI22_X1 U2609 ( .A1(n13891), .A2(n12170), .B1(n13725), .B2(n12164), .ZN(
        n4363) );
  AOI221_X1 U2610 ( .B1(n12278), .B2(n11648), .C1(n12272), .C2(n11468), .A(
        n4336), .ZN(n4331) );
  OAI22_X1 U2611 ( .A1(n14358), .A2(n12266), .B1(n13488), .B2(n12260), .ZN(
        n4336) );
  AOI221_X1 U2612 ( .B1(n12182), .B2(n14077), .C1(n12176), .C2(n14124), .A(
        n4344), .ZN(n4339) );
  OAI22_X1 U2613 ( .A1(n13890), .A2(n12170), .B1(n13724), .B2(n12164), .ZN(
        n4344) );
  AOI221_X1 U2614 ( .B1(n12278), .B2(n11649), .C1(n12272), .C2(n11469), .A(
        n4317), .ZN(n4312) );
  OAI22_X1 U2615 ( .A1(n14340), .A2(n12266), .B1(n13487), .B2(n12260), .ZN(
        n4317) );
  AOI221_X1 U2616 ( .B1(n12182), .B2(n14076), .C1(n12176), .C2(n14123), .A(
        n4325), .ZN(n4320) );
  OAI22_X1 U2617 ( .A1(n13889), .A2(n12170), .B1(n13723), .B2(n12164), .ZN(
        n4325) );
  AOI221_X1 U2618 ( .B1(n12278), .B2(n11650), .C1(n12272), .C2(n11470), .A(
        n4298), .ZN(n4293) );
  OAI22_X1 U2619 ( .A1(n14339), .A2(n12266), .B1(n13486), .B2(n12260), .ZN(
        n4298) );
  AOI221_X1 U2620 ( .B1(n12182), .B2(n14075), .C1(n12176), .C2(n14122), .A(
        n4306), .ZN(n4301) );
  OAI22_X1 U2621 ( .A1(n13888), .A2(n12170), .B1(n13722), .B2(n12164), .ZN(
        n4306) );
  AOI221_X1 U2622 ( .B1(n12278), .B2(n11651), .C1(n12272), .C2(n11471), .A(
        n4279), .ZN(n4274) );
  OAI22_X1 U2623 ( .A1(n14338), .A2(n12266), .B1(n13485), .B2(n12260), .ZN(
        n4279) );
  AOI221_X1 U2624 ( .B1(n12182), .B2(n14074), .C1(n12176), .C2(n14121), .A(
        n4287), .ZN(n4282) );
  OAI22_X1 U2625 ( .A1(n13887), .A2(n12170), .B1(n13721), .B2(n12164), .ZN(
        n4287) );
  AOI221_X1 U2626 ( .B1(n12278), .B2(n11652), .C1(n12272), .C2(n11472), .A(
        n4260), .ZN(n4255) );
  OAI22_X1 U2627 ( .A1(n14337), .A2(n12266), .B1(n13484), .B2(n12260), .ZN(
        n4260) );
  AOI221_X1 U2628 ( .B1(n12182), .B2(n14073), .C1(n12176), .C2(n14120), .A(
        n4268), .ZN(n4263) );
  OAI22_X1 U2629 ( .A1(n13886), .A2(n12170), .B1(n13720), .B2(n12164), .ZN(
        n4268) );
  AOI221_X1 U2630 ( .B1(n12278), .B2(n11653), .C1(n12272), .C2(n11473), .A(
        n4241), .ZN(n4236) );
  OAI22_X1 U2631 ( .A1(n14336), .A2(n12266), .B1(n13483), .B2(n12260), .ZN(
        n4241) );
  AOI221_X1 U2632 ( .B1(n12182), .B2(n14072), .C1(n12176), .C2(n14119), .A(
        n4249), .ZN(n4244) );
  OAI22_X1 U2633 ( .A1(n13885), .A2(n12170), .B1(n13719), .B2(n12164), .ZN(
        n4249) );
  AOI221_X1 U2634 ( .B1(n12279), .B2(n11654), .C1(n12273), .C2(n11474), .A(
        n4222), .ZN(n4217) );
  OAI22_X1 U2635 ( .A1(n14335), .A2(n12267), .B1(n13482), .B2(n12261), .ZN(
        n4222) );
  AOI221_X1 U2636 ( .B1(n12183), .B2(n14071), .C1(n12177), .C2(n14118), .A(
        n4230), .ZN(n4225) );
  OAI22_X1 U2637 ( .A1(n13884), .A2(n12171), .B1(n13718), .B2(n12165), .ZN(
        n4230) );
  AOI221_X1 U2638 ( .B1(n12279), .B2(n11655), .C1(n12273), .C2(n11475), .A(
        n4203), .ZN(n4198) );
  OAI22_X1 U2639 ( .A1(n14334), .A2(n12267), .B1(n13481), .B2(n12261), .ZN(
        n4203) );
  AOI221_X1 U2640 ( .B1(n12183), .B2(n14070), .C1(n12177), .C2(n14117), .A(
        n4211), .ZN(n4206) );
  OAI22_X1 U2641 ( .A1(n13883), .A2(n12171), .B1(n13717), .B2(n12165), .ZN(
        n4211) );
  AOI221_X1 U2642 ( .B1(n12279), .B2(n11656), .C1(n12273), .C2(n11476), .A(
        n4184), .ZN(n4179) );
  OAI22_X1 U2643 ( .A1(n14333), .A2(n12267), .B1(n13480), .B2(n12261), .ZN(
        n4184) );
  AOI221_X1 U2644 ( .B1(n12183), .B2(n14069), .C1(n12177), .C2(n14116), .A(
        n4192), .ZN(n4187) );
  OAI22_X1 U2645 ( .A1(n13882), .A2(n12171), .B1(n13716), .B2(n12165), .ZN(
        n4192) );
  AOI221_X1 U2646 ( .B1(n12279), .B2(n11657), .C1(n12273), .C2(n11477), .A(
        n4165), .ZN(n4160) );
  OAI22_X1 U2647 ( .A1(n14332), .A2(n12267), .B1(n13479), .B2(n12261), .ZN(
        n4165) );
  AOI221_X1 U2648 ( .B1(n12183), .B2(n14068), .C1(n12177), .C2(n14115), .A(
        n4173), .ZN(n4168) );
  OAI22_X1 U2649 ( .A1(n13881), .A2(n12171), .B1(n13715), .B2(n12165), .ZN(
        n4173) );
  AOI221_X1 U2650 ( .B1(n12279), .B2(n11658), .C1(n12273), .C2(n11478), .A(
        n4146), .ZN(n4141) );
  OAI22_X1 U2651 ( .A1(n13535), .A2(n12267), .B1(n13478), .B2(n12261), .ZN(
        n4146) );
  AOI221_X1 U2652 ( .B1(n12183), .B2(n14067), .C1(n12177), .C2(n14114), .A(
        n4154), .ZN(n4149) );
  OAI22_X1 U2653 ( .A1(n13880), .A2(n12171), .B1(n13714), .B2(n12165), .ZN(
        n4154) );
  AOI221_X1 U2654 ( .B1(n12279), .B2(n11659), .C1(n12273), .C2(n11479), .A(
        n4127), .ZN(n4122) );
  OAI22_X1 U2655 ( .A1(n14331), .A2(n12267), .B1(n13477), .B2(n12261), .ZN(
        n4127) );
  AOI221_X1 U2656 ( .B1(n12183), .B2(n14066), .C1(n12177), .C2(n14113), .A(
        n4135), .ZN(n4130) );
  OAI22_X1 U2657 ( .A1(n13879), .A2(n12171), .B1(n13713), .B2(n12165), .ZN(
        n4135) );
  AOI221_X1 U2658 ( .B1(n12279), .B2(n11660), .C1(n12273), .C2(n11480), .A(
        n4108), .ZN(n4103) );
  OAI22_X1 U2659 ( .A1(n14330), .A2(n12267), .B1(n13476), .B2(n12261), .ZN(
        n4108) );
  AOI221_X1 U2660 ( .B1(n12183), .B2(n14065), .C1(n12177), .C2(n14112), .A(
        n4116), .ZN(n4111) );
  OAI22_X1 U2661 ( .A1(n13878), .A2(n12171), .B1(n13712), .B2(n12165), .ZN(
        n4116) );
  AOI221_X1 U2662 ( .B1(n12279), .B2(n11661), .C1(n12273), .C2(n11481), .A(
        n4089), .ZN(n4084) );
  OAI22_X1 U2663 ( .A1(n14329), .A2(n12267), .B1(n13475), .B2(n12261), .ZN(
        n4089) );
  AOI221_X1 U2664 ( .B1(n12183), .B2(n14064), .C1(n12177), .C2(n14111), .A(
        n4097), .ZN(n4092) );
  OAI22_X1 U2665 ( .A1(n13877), .A2(n12171), .B1(n13711), .B2(n12165), .ZN(
        n4097) );
  AOI221_X1 U2666 ( .B1(n12279), .B2(n11662), .C1(n12273), .C2(n11482), .A(
        n4070), .ZN(n4065) );
  OAI22_X1 U2667 ( .A1(n13534), .A2(n12267), .B1(n13474), .B2(n12261), .ZN(
        n4070) );
  AOI221_X1 U2668 ( .B1(n12183), .B2(n14063), .C1(n12177), .C2(n14110), .A(
        n4078), .ZN(n4073) );
  OAI22_X1 U2669 ( .A1(n13876), .A2(n12171), .B1(n13710), .B2(n12165), .ZN(
        n4078) );
  AOI221_X1 U2670 ( .B1(n12279), .B2(n11663), .C1(n12273), .C2(n11483), .A(
        n4051), .ZN(n4046) );
  OAI22_X1 U2671 ( .A1(n13533), .A2(n12267), .B1(n13473), .B2(n12261), .ZN(
        n4051) );
  AOI221_X1 U2672 ( .B1(n12183), .B2(n14062), .C1(n12177), .C2(n14109), .A(
        n4059), .ZN(n4054) );
  OAI22_X1 U2673 ( .A1(n13875), .A2(n12171), .B1(n13709), .B2(n12165), .ZN(
        n4059) );
  AOI221_X1 U2674 ( .B1(n12279), .B2(n11664), .C1(n12273), .C2(n11484), .A(
        n4032), .ZN(n4027) );
  OAI22_X1 U2675 ( .A1(n13532), .A2(n12267), .B1(n13472), .B2(n12261), .ZN(
        n4032) );
  AOI221_X1 U2676 ( .B1(n12183), .B2(n14061), .C1(n12177), .C2(n14108), .A(
        n4040), .ZN(n4035) );
  OAI22_X1 U2677 ( .A1(n13874), .A2(n12171), .B1(n13708), .B2(n12165), .ZN(
        n4040) );
  AOI221_X1 U2678 ( .B1(n12279), .B2(n11665), .C1(n12273), .C2(n11485), .A(
        n4013), .ZN(n4008) );
  OAI22_X1 U2679 ( .A1(n13531), .A2(n12267), .B1(n13471), .B2(n12261), .ZN(
        n4013) );
  AOI221_X1 U2680 ( .B1(n12183), .B2(n14060), .C1(n12177), .C2(n14107), .A(
        n4021), .ZN(n4016) );
  OAI22_X1 U2681 ( .A1(n13873), .A2(n12171), .B1(n13707), .B2(n12165), .ZN(
        n4021) );
  AOI221_X1 U2682 ( .B1(n12280), .B2(n11666), .C1(n12274), .C2(n11486), .A(
        n3994), .ZN(n3989) );
  OAI22_X1 U2683 ( .A1(n13530), .A2(n12268), .B1(n13470), .B2(n12262), .ZN(
        n3994) );
  AOI221_X1 U2684 ( .B1(n12184), .B2(n13928), .C1(n12178), .C2(n13988), .A(
        n4002), .ZN(n3997) );
  OAI22_X1 U2685 ( .A1(n13872), .A2(n12172), .B1(n13706), .B2(n12166), .ZN(
        n4002) );
  AOI221_X1 U2686 ( .B1(n12280), .B2(n11667), .C1(n12274), .C2(n11487), .A(
        n3975), .ZN(n3970) );
  OAI22_X1 U2687 ( .A1(n13529), .A2(n12268), .B1(n13469), .B2(n12262), .ZN(
        n3975) );
  AOI221_X1 U2688 ( .B1(n12184), .B2(n13927), .C1(n12178), .C2(n13987), .A(
        n3983), .ZN(n3978) );
  OAI22_X1 U2689 ( .A1(n13871), .A2(n12172), .B1(n13705), .B2(n12166), .ZN(
        n3983) );
  AOI221_X1 U2690 ( .B1(n12280), .B2(n11668), .C1(n12274), .C2(n11488), .A(
        n3956), .ZN(n3951) );
  OAI22_X1 U2691 ( .A1(n13528), .A2(n12268), .B1(n13468), .B2(n12262), .ZN(
        n3956) );
  AOI221_X1 U2692 ( .B1(n12184), .B2(n13926), .C1(n12178), .C2(n13986), .A(
        n3964), .ZN(n3959) );
  OAI22_X1 U2693 ( .A1(n13870), .A2(n12172), .B1(n13704), .B2(n12166), .ZN(
        n3964) );
  AOI221_X1 U2694 ( .B1(n12280), .B2(n11669), .C1(n12274), .C2(n11489), .A(
        n3937), .ZN(n3932) );
  OAI22_X1 U2695 ( .A1(n13527), .A2(n12268), .B1(n13467), .B2(n12262), .ZN(
        n3937) );
  AOI221_X1 U2696 ( .B1(n12184), .B2(n13925), .C1(n12178), .C2(n13985), .A(
        n3945), .ZN(n3940) );
  OAI22_X1 U2697 ( .A1(n13869), .A2(n12172), .B1(n13703), .B2(n12166), .ZN(
        n3945) );
  AOI221_X1 U2698 ( .B1(n12280), .B2(n11670), .C1(n12274), .C2(n11490), .A(
        n3918), .ZN(n3913) );
  OAI22_X1 U2699 ( .A1(n13526), .A2(n12268), .B1(n13466), .B2(n12262), .ZN(
        n3918) );
  AOI221_X1 U2700 ( .B1(n12184), .B2(n13924), .C1(n12178), .C2(n13984), .A(
        n3926), .ZN(n3921) );
  OAI22_X1 U2701 ( .A1(n14059), .A2(n12172), .B1(n13702), .B2(n12166), .ZN(
        n3926) );
  AOI221_X1 U2702 ( .B1(n12280), .B2(n11671), .C1(n12274), .C2(n11491), .A(
        n3899), .ZN(n3894) );
  OAI22_X1 U2703 ( .A1(n13525), .A2(n12268), .B1(n13465), .B2(n12262), .ZN(
        n3899) );
  AOI221_X1 U2704 ( .B1(n12184), .B2(n13923), .C1(n12178), .C2(n13983), .A(
        n3907), .ZN(n3902) );
  OAI22_X1 U2705 ( .A1(n14058), .A2(n12172), .B1(n13701), .B2(n12166), .ZN(
        n3907) );
  AOI221_X1 U2706 ( .B1(n12280), .B2(n11672), .C1(n12274), .C2(n11492), .A(
        n3880), .ZN(n3875) );
  OAI22_X1 U2707 ( .A1(n13524), .A2(n12268), .B1(n13464), .B2(n12262), .ZN(
        n3880) );
  AOI221_X1 U2708 ( .B1(n12184), .B2(n13922), .C1(n12178), .C2(n13982), .A(
        n3888), .ZN(n3883) );
  OAI22_X1 U2709 ( .A1(n14057), .A2(n12172), .B1(n13700), .B2(n12166), .ZN(
        n3888) );
  AOI221_X1 U2710 ( .B1(n12280), .B2(n11673), .C1(n12274), .C2(n11493), .A(
        n3861), .ZN(n3856) );
  OAI22_X1 U2711 ( .A1(n13523), .A2(n12268), .B1(n13463), .B2(n12262), .ZN(
        n3861) );
  AOI221_X1 U2712 ( .B1(n12184), .B2(n13921), .C1(n12178), .C2(n13981), .A(
        n3869), .ZN(n3864) );
  OAI22_X1 U2713 ( .A1(n14056), .A2(n12172), .B1(n13699), .B2(n12166), .ZN(
        n3869) );
  AOI221_X1 U2714 ( .B1(n12280), .B2(n11674), .C1(n12274), .C2(n11494), .A(
        n3842), .ZN(n3837) );
  OAI22_X1 U2715 ( .A1(n13522), .A2(n12268), .B1(n13462), .B2(n12262), .ZN(
        n3842) );
  AOI221_X1 U2716 ( .B1(n12184), .B2(n13920), .C1(n12178), .C2(n13980), .A(
        n3850), .ZN(n3845) );
  OAI22_X1 U2717 ( .A1(n14055), .A2(n12172), .B1(n13698), .B2(n12166), .ZN(
        n3850) );
  AOI221_X1 U2718 ( .B1(n12280), .B2(n11675), .C1(n12274), .C2(n11495), .A(
        n3823), .ZN(n3818) );
  OAI22_X1 U2719 ( .A1(n13521), .A2(n12268), .B1(n13461), .B2(n12262), .ZN(
        n3823) );
  AOI221_X1 U2720 ( .B1(n12184), .B2(n13919), .C1(n12178), .C2(n13979), .A(
        n3831), .ZN(n3826) );
  OAI22_X1 U2721 ( .A1(n14054), .A2(n12172), .B1(n13697), .B2(n12166), .ZN(
        n3831) );
  AOI221_X1 U2722 ( .B1(n12280), .B2(n11676), .C1(n12274), .C2(n11496), .A(
        n3804), .ZN(n3799) );
  OAI22_X1 U2723 ( .A1(n13520), .A2(n12268), .B1(n13460), .B2(n12262), .ZN(
        n3804) );
  AOI221_X1 U2724 ( .B1(n12184), .B2(n13918), .C1(n12178), .C2(n13978), .A(
        n3812), .ZN(n3807) );
  OAI22_X1 U2725 ( .A1(n14053), .A2(n12172), .B1(n13696), .B2(n12166), .ZN(
        n3812) );
  AOI221_X1 U2726 ( .B1(n12280), .B2(n11677), .C1(n12274), .C2(n11497), .A(
        n3785), .ZN(n3780) );
  OAI22_X1 U2727 ( .A1(n13519), .A2(n12268), .B1(n13459), .B2(n12262), .ZN(
        n3785) );
  AOI221_X1 U2728 ( .B1(n12184), .B2(n13917), .C1(n12178), .C2(n13977), .A(
        n3793), .ZN(n3788) );
  OAI22_X1 U2729 ( .A1(n14052), .A2(n12172), .B1(n13695), .B2(n12166), .ZN(
        n3793) );
  AOI221_X1 U2730 ( .B1(n12281), .B2(n11678), .C1(n12275), .C2(n11498), .A(
        n3766), .ZN(n3761) );
  OAI22_X1 U2731 ( .A1(n13518), .A2(n12269), .B1(n13458), .B2(n12263), .ZN(
        n3766) );
  AOI221_X1 U2732 ( .B1(n12185), .B2(n13916), .C1(n12179), .C2(n13976), .A(
        n3774), .ZN(n3769) );
  OAI22_X1 U2733 ( .A1(n14051), .A2(n12173), .B1(n13694), .B2(n12167), .ZN(
        n3774) );
  AOI221_X1 U2734 ( .B1(n12281), .B2(n11679), .C1(n12275), .C2(n11499), .A(
        n3747), .ZN(n3742) );
  OAI22_X1 U2735 ( .A1(n13517), .A2(n12269), .B1(n13457), .B2(n12263), .ZN(
        n3747) );
  AOI221_X1 U2736 ( .B1(n12185), .B2(n13915), .C1(n12179), .C2(n13975), .A(
        n3755), .ZN(n3750) );
  OAI22_X1 U2737 ( .A1(n14050), .A2(n12173), .B1(n13693), .B2(n12167), .ZN(
        n3755) );
  AOI221_X1 U2738 ( .B1(n12281), .B2(n11680), .C1(n12275), .C2(n11500), .A(
        n3728), .ZN(n3723) );
  OAI22_X1 U2739 ( .A1(n13516), .A2(n12269), .B1(n13456), .B2(n12263), .ZN(
        n3728) );
  AOI221_X1 U2740 ( .B1(n12185), .B2(n13914), .C1(n12179), .C2(n13974), .A(
        n3736), .ZN(n3731) );
  OAI22_X1 U2741 ( .A1(n14049), .A2(n12173), .B1(n13692), .B2(n12167), .ZN(
        n3736) );
  AOI221_X1 U2742 ( .B1(n12281), .B2(n11681), .C1(n12275), .C2(n11501), .A(
        n3709), .ZN(n3704) );
  OAI22_X1 U2743 ( .A1(n14460), .A2(n12269), .B1(n13455), .B2(n12263), .ZN(
        n3709) );
  AOI221_X1 U2744 ( .B1(n12185), .B2(n13913), .C1(n12179), .C2(n13973), .A(
        n3717), .ZN(n3712) );
  OAI22_X1 U2745 ( .A1(n14048), .A2(n12173), .B1(n13691), .B2(n12167), .ZN(
        n3717) );
  AOI221_X1 U2746 ( .B1(n12281), .B2(n11682), .C1(n12275), .C2(n11502), .A(
        n3690), .ZN(n3685) );
  OAI22_X1 U2747 ( .A1(n14459), .A2(n12269), .B1(n13454), .B2(n12263), .ZN(
        n3690) );
  AOI221_X1 U2748 ( .B1(n12185), .B2(n13912), .C1(n12179), .C2(n13972), .A(
        n3698), .ZN(n3693) );
  OAI22_X1 U2749 ( .A1(n14047), .A2(n12173), .B1(n13690), .B2(n12167), .ZN(
        n3698) );
  AOI221_X1 U2750 ( .B1(n12281), .B2(n11683), .C1(n12275), .C2(n11503), .A(
        n3671), .ZN(n3666) );
  OAI22_X1 U2751 ( .A1(n14458), .A2(n12269), .B1(n13453), .B2(n12263), .ZN(
        n3671) );
  AOI221_X1 U2752 ( .B1(n12185), .B2(n13911), .C1(n12179), .C2(n13971), .A(
        n3679), .ZN(n3674) );
  OAI22_X1 U2753 ( .A1(n14046), .A2(n12173), .B1(n13689), .B2(n12167), .ZN(
        n3679) );
  AOI221_X1 U2754 ( .B1(n12281), .B2(n11684), .C1(n12275), .C2(n11504), .A(
        n3652), .ZN(n3647) );
  OAI22_X1 U2755 ( .A1(n14457), .A2(n12269), .B1(n13452), .B2(n12263), .ZN(
        n3652) );
  AOI221_X1 U2756 ( .B1(n12185), .B2(n13910), .C1(n12179), .C2(n13970), .A(
        n3660), .ZN(n3655) );
  OAI22_X1 U2757 ( .A1(n14045), .A2(n12173), .B1(n13688), .B2(n12167), .ZN(
        n3660) );
  AOI221_X1 U2758 ( .B1(n12281), .B2(n11685), .C1(n12275), .C2(n11505), .A(
        n3633), .ZN(n3628) );
  OAI22_X1 U2759 ( .A1(n13515), .A2(n12269), .B1(n13451), .B2(n12263), .ZN(
        n3633) );
  AOI221_X1 U2760 ( .B1(n12185), .B2(n13909), .C1(n12179), .C2(n13969), .A(
        n3641), .ZN(n3636) );
  OAI22_X1 U2761 ( .A1(n14044), .A2(n12173), .B1(n13687), .B2(n12167), .ZN(
        n3641) );
  AOI221_X1 U2762 ( .B1(n12281), .B2(n11686), .C1(n12275), .C2(n11506), .A(
        n3614), .ZN(n3609) );
  OAI22_X1 U2763 ( .A1(n13514), .A2(n12269), .B1(n13450), .B2(n12263), .ZN(
        n3614) );
  AOI221_X1 U2764 ( .B1(n12185), .B2(n13908), .C1(n12179), .C2(n13968), .A(
        n3622), .ZN(n3617) );
  OAI22_X1 U2765 ( .A1(n14043), .A2(n12173), .B1(n13686), .B2(n12167), .ZN(
        n3622) );
  AOI221_X1 U2766 ( .B1(n12281), .B2(n11687), .C1(n12275), .C2(n11507), .A(
        n3595), .ZN(n3590) );
  OAI22_X1 U2767 ( .A1(n13513), .A2(n12269), .B1(n13449), .B2(n12263), .ZN(
        n3595) );
  AOI221_X1 U2768 ( .B1(n12185), .B2(n13907), .C1(n12179), .C2(n13967), .A(
        n3603), .ZN(n3598) );
  OAI22_X1 U2769 ( .A1(n14042), .A2(n12173), .B1(n13685), .B2(n12167), .ZN(
        n3603) );
  AOI221_X1 U2770 ( .B1(n12281), .B2(n11688), .C1(n12275), .C2(n11508), .A(
        n3576), .ZN(n3571) );
  OAI22_X1 U2771 ( .A1(n13512), .A2(n12269), .B1(n13448), .B2(n12263), .ZN(
        n3576) );
  AOI221_X1 U2772 ( .B1(n12185), .B2(n13906), .C1(n12179), .C2(n13966), .A(
        n3584), .ZN(n3579) );
  OAI22_X1 U2773 ( .A1(n14041), .A2(n12173), .B1(n13684), .B2(n12167), .ZN(
        n3584) );
  AOI221_X1 U2774 ( .B1(n12281), .B2(n11689), .C1(n12275), .C2(n11509), .A(
        n3557), .ZN(n3552) );
  OAI22_X1 U2775 ( .A1(n13511), .A2(n12269), .B1(n13447), .B2(n12263), .ZN(
        n3557) );
  AOI221_X1 U2776 ( .B1(n12185), .B2(n13905), .C1(n12179), .C2(n13965), .A(
        n3565), .ZN(n3560) );
  OAI22_X1 U2777 ( .A1(n14040), .A2(n12173), .B1(n13683), .B2(n12167), .ZN(
        n3565) );
  AOI221_X1 U2778 ( .B1(n12282), .B2(n11690), .C1(n12276), .C2(n11510), .A(
        n3538), .ZN(n3533) );
  OAI22_X1 U2779 ( .A1(n13510), .A2(n12270), .B1(n13446), .B2(n12264), .ZN(
        n3538) );
  AOI221_X1 U2780 ( .B1(n12186), .B2(n13904), .C1(n12180), .C2(n13964), .A(
        n3546), .ZN(n3541) );
  OAI22_X1 U2781 ( .A1(n14039), .A2(n12174), .B1(n13682), .B2(n12168), .ZN(
        n3546) );
  AOI221_X1 U2782 ( .B1(n12282), .B2(n11691), .C1(n12276), .C2(n11511), .A(
        n3519), .ZN(n3514) );
  OAI22_X1 U2783 ( .A1(n13509), .A2(n12270), .B1(n13445), .B2(n12264), .ZN(
        n3519) );
  AOI221_X1 U2784 ( .B1(n12186), .B2(n13903), .C1(n12180), .C2(n13963), .A(
        n3527), .ZN(n3522) );
  OAI22_X1 U2785 ( .A1(n14038), .A2(n12174), .B1(n13681), .B2(n12168), .ZN(
        n3527) );
  AOI221_X1 U2786 ( .B1(n12282), .B2(n11692), .C1(n12276), .C2(n11512), .A(
        n3500), .ZN(n3495) );
  OAI22_X1 U2787 ( .A1(n13508), .A2(n12270), .B1(n13444), .B2(n12264), .ZN(
        n3500) );
  AOI221_X1 U2788 ( .B1(n12186), .B2(n13902), .C1(n12180), .C2(n13962), .A(
        n3508), .ZN(n3503) );
  OAI22_X1 U2789 ( .A1(n14037), .A2(n12174), .B1(n13680), .B2(n12168), .ZN(
        n3508) );
  AOI221_X1 U2790 ( .B1(n12282), .B2(n11693), .C1(n12276), .C2(n11513), .A(
        n3481), .ZN(n3476) );
  OAI22_X1 U2791 ( .A1(n13507), .A2(n12270), .B1(n13443), .B2(n12264), .ZN(
        n3481) );
  AOI221_X1 U2792 ( .B1(n12186), .B2(n13901), .C1(n12180), .C2(n13961), .A(
        n3489), .ZN(n3484) );
  OAI22_X1 U2793 ( .A1(n14036), .A2(n12174), .B1(n13679), .B2(n12168), .ZN(
        n3489) );
  AOI221_X1 U2794 ( .B1(n12282), .B2(n11694), .C1(n12276), .C2(n11514), .A(
        n3462), .ZN(n3457) );
  OAI22_X1 U2795 ( .A1(n13506), .A2(n12270), .B1(n13442), .B2(n12264), .ZN(
        n3462) );
  AOI221_X1 U2796 ( .B1(n12186), .B2(n13900), .C1(n12180), .C2(n13960), .A(
        n3470), .ZN(n3465) );
  OAI22_X1 U2797 ( .A1(n13742), .A2(n12174), .B1(n13678), .B2(n12168), .ZN(
        n3470) );
  AOI221_X1 U2798 ( .B1(n12282), .B2(n11695), .C1(n12276), .C2(n11515), .A(
        n3443), .ZN(n3438) );
  OAI22_X1 U2799 ( .A1(n13505), .A2(n12270), .B1(n13441), .B2(n12264), .ZN(
        n3443) );
  AOI221_X1 U2800 ( .B1(n12186), .B2(n13899), .C1(n12180), .C2(n13959), .A(
        n3451), .ZN(n3446) );
  OAI22_X1 U2801 ( .A1(n13741), .A2(n12174), .B1(n13677), .B2(n12168), .ZN(
        n3451) );
  AOI221_X1 U2802 ( .B1(n12282), .B2(n11696), .C1(n12276), .C2(n11516), .A(
        n3424), .ZN(n3419) );
  OAI22_X1 U2803 ( .A1(n13504), .A2(n12270), .B1(n13440), .B2(n12264), .ZN(
        n3424) );
  AOI221_X1 U2804 ( .B1(n12186), .B2(n13898), .C1(n12180), .C2(n13958), .A(
        n3432), .ZN(n3427) );
  OAI22_X1 U2805 ( .A1(n13740), .A2(n12174), .B1(n13676), .B2(n12168), .ZN(
        n3432) );
  AOI221_X1 U2806 ( .B1(n12282), .B2(n11697), .C1(n12276), .C2(n11517), .A(
        n3405), .ZN(n3400) );
  OAI22_X1 U2807 ( .A1(n13503), .A2(n12270), .B1(n13439), .B2(n12264), .ZN(
        n3405) );
  AOI221_X1 U2808 ( .B1(n12186), .B2(n13897), .C1(n12180), .C2(n13957), .A(
        n3413), .ZN(n3408) );
  OAI22_X1 U2809 ( .A1(n13739), .A2(n12174), .B1(n13675), .B2(n12168), .ZN(
        n3413) );
  AOI221_X1 U2810 ( .B1(n12282), .B2(n11698), .C1(n12276), .C2(n11518), .A(
        n3386), .ZN(n3381) );
  OAI22_X1 U2811 ( .A1(n13502), .A2(n12270), .B1(n13438), .B2(n12264), .ZN(
        n3386) );
  AOI221_X1 U2812 ( .B1(n12186), .B2(n13896), .C1(n12180), .C2(n13956), .A(
        n3394), .ZN(n3389) );
  OAI22_X1 U2813 ( .A1(n13738), .A2(n12174), .B1(n13674), .B2(n12168), .ZN(
        n3394) );
  AOI221_X1 U2814 ( .B1(n12282), .B2(n11699), .C1(n12276), .C2(n11519), .A(
        n3367), .ZN(n3362) );
  OAI22_X1 U2815 ( .A1(n13501), .A2(n12270), .B1(n13437), .B2(n12264), .ZN(
        n3367) );
  AOI221_X1 U2816 ( .B1(n12186), .B2(n13895), .C1(n12180), .C2(n13955), .A(
        n3375), .ZN(n3370) );
  OAI22_X1 U2817 ( .A1(n13737), .A2(n12174), .B1(n13673), .B2(n12168), .ZN(
        n3375) );
  AOI221_X1 U2818 ( .B1(n12282), .B2(n11700), .C1(n12276), .C2(n11520), .A(
        n3348), .ZN(n3343) );
  OAI22_X1 U2819 ( .A1(n13500), .A2(n12270), .B1(n13436), .B2(n12264), .ZN(
        n3348) );
  AOI221_X1 U2820 ( .B1(n12186), .B2(n13894), .C1(n12180), .C2(n13954), .A(
        n3356), .ZN(n3351) );
  OAI22_X1 U2821 ( .A1(n13736), .A2(n12174), .B1(n13672), .B2(n12168), .ZN(
        n3356) );
  AOI221_X1 U2822 ( .B1(n12282), .B2(n11701), .C1(n12276), .C2(n11521), .A(
        n3329), .ZN(n3324) );
  OAI22_X1 U2823 ( .A1(n13499), .A2(n12270), .B1(n13435), .B2(n12264), .ZN(
        n3329) );
  AOI221_X1 U2824 ( .B1(n12186), .B2(n13893), .C1(n12180), .C2(n13953), .A(
        n3337), .ZN(n3332) );
  OAI22_X1 U2825 ( .A1(n13735), .A2(n12174), .B1(n13671), .B2(n12168), .ZN(
        n3337) );
  AOI221_X1 U2826 ( .B1(n12187), .B2(n13819), .C1(n12181), .C2(n13823), .A(
        n3318), .ZN(n3313) );
  OAI22_X1 U2827 ( .A1(n13734), .A2(n12175), .B1(n13670), .B2(n12169), .ZN(
        n3318) );
  AOI221_X1 U2828 ( .B1(n12283), .B2(n13860), .C1(n12277), .C2(n13856), .A(
        n3310), .ZN(n3305) );
  OAI22_X1 U2829 ( .A1(n13498), .A2(n12271), .B1(n13434), .B2(n12265), .ZN(
        n3310) );
  AOI221_X1 U2830 ( .B1(n12187), .B2(n13818), .C1(n12181), .C2(n13822), .A(
        n3299), .ZN(n3294) );
  OAI22_X1 U2831 ( .A1(n13733), .A2(n12175), .B1(n13669), .B2(n12169), .ZN(
        n3299) );
  AOI221_X1 U2832 ( .B1(n12283), .B2(n13859), .C1(n12277), .C2(n13855), .A(
        n3291), .ZN(n3286) );
  OAI22_X1 U2833 ( .A1(n13497), .A2(n12271), .B1(n13433), .B2(n12265), .ZN(
        n3291) );
  AOI221_X1 U2834 ( .B1(n12187), .B2(n13817), .C1(n12181), .C2(n13821), .A(
        n3280), .ZN(n3275) );
  OAI22_X1 U2835 ( .A1(n13732), .A2(n12175), .B1(n13668), .B2(n12169), .ZN(
        n3280) );
  AOI221_X1 U2836 ( .B1(n12283), .B2(n13858), .C1(n12277), .C2(n13854), .A(
        n3272), .ZN(n3267) );
  OAI22_X1 U2837 ( .A1(n13496), .A2(n12271), .B1(n13432), .B2(n12265), .ZN(
        n3272) );
  AOI221_X1 U2838 ( .B1(n12187), .B2(n13816), .C1(n12181), .C2(n13820), .A(
        n3255), .ZN(n3240) );
  OAI22_X1 U2839 ( .A1(n13731), .A2(n12175), .B1(n13667), .B2(n12169), .ZN(
        n3255) );
  AOI221_X1 U2840 ( .B1(n12283), .B2(n13857), .C1(n12277), .C2(n13853), .A(
        n3231), .ZN(n3216) );
  OAI22_X1 U2841 ( .A1(n13495), .A2(n12271), .B1(n13431), .B2(n12265), .ZN(
        n3231) );
  AOI221_X1 U2842 ( .B1(n12254), .B2(n11702), .C1(n12248), .C2(n11522), .A(
        n4459), .ZN(n4444) );
  OAI22_X1 U2843 ( .A1(n13650), .A2(n12242), .B1(n13603), .B2(n12236), .ZN(
        n4459) );
  AOI221_X1 U2844 ( .B1(n12158), .B2(n14155), .C1(n12152), .C2(n13831), .A(
        n4471), .ZN(n4460) );
  OAI22_X1 U2845 ( .A1(n13815), .A2(n12146), .B1(n13810), .B2(n12140), .ZN(
        n4471) );
  AOI221_X1 U2846 ( .B1(n12254), .B2(n11703), .C1(n12248), .C2(n11523), .A(
        n4432), .ZN(n4425) );
  OAI22_X1 U2847 ( .A1(n13649), .A2(n12242), .B1(n13602), .B2(n12236), .ZN(
        n4432) );
  AOI221_X1 U2848 ( .B1(n12158), .B2(n14152), .C1(n12152), .C2(n13830), .A(
        n4440), .ZN(n4433) );
  OAI22_X1 U2849 ( .A1(n13814), .A2(n12146), .B1(n13809), .B2(n12140), .ZN(
        n4440) );
  AOI221_X1 U2850 ( .B1(n12254), .B2(n11704), .C1(n12248), .C2(n11524), .A(
        n4413), .ZN(n4406) );
  OAI22_X1 U2851 ( .A1(n13648), .A2(n12242), .B1(n13601), .B2(n12236), .ZN(
        n4413) );
  AOI221_X1 U2852 ( .B1(n12158), .B2(n14151), .C1(n12152), .C2(n13829), .A(
        n4421), .ZN(n4414) );
  OAI22_X1 U2853 ( .A1(n13813), .A2(n12146), .B1(n13808), .B2(n12140), .ZN(
        n4421) );
  AOI221_X1 U2854 ( .B1(n12254), .B2(n11705), .C1(n12248), .C2(n11525), .A(
        n4394), .ZN(n4387) );
  OAI22_X1 U2855 ( .A1(n13647), .A2(n12242), .B1(n13600), .B2(n12236), .ZN(
        n4394) );
  AOI221_X1 U2856 ( .B1(n12158), .B2(n14149), .C1(n12152), .C2(n13828), .A(
        n4402), .ZN(n4395) );
  OAI22_X1 U2857 ( .A1(n13812), .A2(n12146), .B1(n13807), .B2(n12140), .ZN(
        n4402) );
  AOI221_X1 U2858 ( .B1(n12254), .B2(n11706), .C1(n12248), .C2(n11526), .A(
        n4375), .ZN(n4368) );
  OAI22_X1 U2859 ( .A1(n14357), .A2(n12242), .B1(n13599), .B2(n12236), .ZN(
        n4375) );
  AOI221_X1 U2860 ( .B1(n12158), .B2(n14150), .C1(n12152), .C2(n14215), .A(
        n4383), .ZN(n4376) );
  OAI22_X1 U2861 ( .A1(n13811), .A2(n12146), .B1(n13806), .B2(n12140), .ZN(
        n4383) );
  AOI221_X1 U2862 ( .B1(n12254), .B2(n11707), .C1(n12248), .C2(n11527), .A(
        n4356), .ZN(n4349) );
  OAI22_X1 U2863 ( .A1(n14356), .A2(n12242), .B1(n13598), .B2(n12236), .ZN(
        n4356) );
  AOI221_X1 U2864 ( .B1(n12158), .B2(n14148), .C1(n12152), .C2(n14214), .A(
        n4364), .ZN(n4357) );
  OAI22_X1 U2865 ( .A1(n14035), .A2(n12146), .B1(n13805), .B2(n12140), .ZN(
        n4364) );
  AOI221_X1 U2866 ( .B1(n12254), .B2(n11708), .C1(n12248), .C2(n11528), .A(
        n4337), .ZN(n4330) );
  OAI22_X1 U2867 ( .A1(n14355), .A2(n12242), .B1(n13597), .B2(n12236), .ZN(
        n4337) );
  AOI221_X1 U2868 ( .B1(n12158), .B2(n14147), .C1(n12152), .C2(n14213), .A(
        n4345), .ZN(n4338) );
  OAI22_X1 U2869 ( .A1(n14034), .A2(n12146), .B1(n13804), .B2(n12140), .ZN(
        n4345) );
  AOI221_X1 U2870 ( .B1(n12254), .B2(n11709), .C1(n12248), .C2(n11529), .A(
        n4318), .ZN(n4311) );
  OAI22_X1 U2871 ( .A1(n14354), .A2(n12242), .B1(n13596), .B2(n12236), .ZN(
        n4318) );
  AOI221_X1 U2872 ( .B1(n12158), .B2(n14146), .C1(n12152), .C2(n14212), .A(
        n4326), .ZN(n4319) );
  OAI22_X1 U2873 ( .A1(n14033), .A2(n12146), .B1(n13803), .B2(n12140), .ZN(
        n4326) );
  AOI221_X1 U2874 ( .B1(n12254), .B2(n11710), .C1(n12248), .C2(n11530), .A(
        n4299), .ZN(n4292) );
  OAI22_X1 U2875 ( .A1(n14353), .A2(n12242), .B1(n13595), .B2(n12236), .ZN(
        n4299) );
  AOI221_X1 U2876 ( .B1(n12158), .B2(n14145), .C1(n12152), .C2(n14211), .A(
        n4307), .ZN(n4300) );
  OAI22_X1 U2877 ( .A1(n14032), .A2(n12146), .B1(n13802), .B2(n12140), .ZN(
        n4307) );
  AOI221_X1 U2878 ( .B1(n12254), .B2(n11711), .C1(n12248), .C2(n11531), .A(
        n4280), .ZN(n4273) );
  OAI22_X1 U2879 ( .A1(n14352), .A2(n12242), .B1(n13594), .B2(n12236), .ZN(
        n4280) );
  AOI221_X1 U2880 ( .B1(n12158), .B2(n14144), .C1(n12152), .C2(n14210), .A(
        n4288), .ZN(n4281) );
  OAI22_X1 U2881 ( .A1(n14031), .A2(n12146), .B1(n13801), .B2(n12140), .ZN(
        n4288) );
  AOI221_X1 U2882 ( .B1(n12254), .B2(n11712), .C1(n12248), .C2(n11532), .A(
        n4261), .ZN(n4254) );
  OAI22_X1 U2883 ( .A1(n14351), .A2(n12242), .B1(n13593), .B2(n12236), .ZN(
        n4261) );
  AOI221_X1 U2884 ( .B1(n12158), .B2(n14143), .C1(n12152), .C2(n14209), .A(
        n4269), .ZN(n4262) );
  OAI22_X1 U2885 ( .A1(n14030), .A2(n12146), .B1(n13800), .B2(n12140), .ZN(
        n4269) );
  AOI221_X1 U2886 ( .B1(n12254), .B2(n11713), .C1(n12248), .C2(n11533), .A(
        n4242), .ZN(n4235) );
  OAI22_X1 U2887 ( .A1(n14350), .A2(n12242), .B1(n13592), .B2(n12236), .ZN(
        n4242) );
  AOI221_X1 U2888 ( .B1(n12158), .B2(n14142), .C1(n12152), .C2(n14208), .A(
        n4250), .ZN(n4243) );
  OAI22_X1 U2889 ( .A1(n14029), .A2(n12146), .B1(n13799), .B2(n12140), .ZN(
        n4250) );
  AOI221_X1 U2890 ( .B1(n12255), .B2(n11714), .C1(n12249), .C2(n11534), .A(
        n4223), .ZN(n4216) );
  OAI22_X1 U2891 ( .A1(n14349), .A2(n12243), .B1(n13591), .B2(n12237), .ZN(
        n4223) );
  AOI221_X1 U2892 ( .B1(n12159), .B2(n14141), .C1(n12153), .C2(n14207), .A(
        n4231), .ZN(n4224) );
  OAI22_X1 U2893 ( .A1(n14028), .A2(n12147), .B1(n13798), .B2(n12141), .ZN(
        n4231) );
  AOI221_X1 U2894 ( .B1(n12255), .B2(n11715), .C1(n12249), .C2(n11535), .A(
        n4204), .ZN(n4197) );
  OAI22_X1 U2895 ( .A1(n14348), .A2(n12243), .B1(n13590), .B2(n12237), .ZN(
        n4204) );
  AOI221_X1 U2896 ( .B1(n12159), .B2(n14140), .C1(n12153), .C2(n14206), .A(
        n4212), .ZN(n4205) );
  OAI22_X1 U2897 ( .A1(n14027), .A2(n12147), .B1(n13797), .B2(n12141), .ZN(
        n4212) );
  AOI221_X1 U2898 ( .B1(n12255), .B2(n11716), .C1(n12249), .C2(n11536), .A(
        n4185), .ZN(n4178) );
  OAI22_X1 U2899 ( .A1(n14347), .A2(n12243), .B1(n13589), .B2(n12237), .ZN(
        n4185) );
  AOI221_X1 U2900 ( .B1(n12159), .B2(n14139), .C1(n12153), .C2(n14205), .A(
        n4193), .ZN(n4186) );
  OAI22_X1 U2901 ( .A1(n14026), .A2(n12147), .B1(n13796), .B2(n12141), .ZN(
        n4193) );
  AOI221_X1 U2902 ( .B1(n12255), .B2(n11717), .C1(n12249), .C2(n11537), .A(
        n4166), .ZN(n4159) );
  OAI22_X1 U2903 ( .A1(n14346), .A2(n12243), .B1(n13588), .B2(n12237), .ZN(
        n4166) );
  AOI221_X1 U2904 ( .B1(n12159), .B2(n14138), .C1(n12153), .C2(n14204), .A(
        n4174), .ZN(n4167) );
  OAI22_X1 U2905 ( .A1(n14025), .A2(n12147), .B1(n13795), .B2(n12141), .ZN(
        n4174) );
  AOI221_X1 U2906 ( .B1(n12255), .B2(n11718), .C1(n12249), .C2(n11538), .A(
        n4147), .ZN(n4140) );
  OAI22_X1 U2907 ( .A1(n13646), .A2(n12243), .B1(n13587), .B2(n12237), .ZN(
        n4147) );
  AOI221_X1 U2908 ( .B1(n12159), .B2(n14137), .C1(n12153), .C2(n14203), .A(
        n4155), .ZN(n4148) );
  OAI22_X1 U2909 ( .A1(n13952), .A2(n12147), .B1(n13794), .B2(n12141), .ZN(
        n4155) );
  AOI221_X1 U2910 ( .B1(n12255), .B2(n11719), .C1(n12249), .C2(n11539), .A(
        n4128), .ZN(n4121) );
  OAI22_X1 U2911 ( .A1(n14345), .A2(n12243), .B1(n13586), .B2(n12237), .ZN(
        n4128) );
  AOI221_X1 U2912 ( .B1(n12159), .B2(n14136), .C1(n12153), .C2(n14202), .A(
        n4136), .ZN(n4129) );
  OAI22_X1 U2913 ( .A1(n13951), .A2(n12147), .B1(n13793), .B2(n12141), .ZN(
        n4136) );
  AOI221_X1 U2914 ( .B1(n12255), .B2(n11720), .C1(n12249), .C2(n11540), .A(
        n4109), .ZN(n4102) );
  OAI22_X1 U2915 ( .A1(n14344), .A2(n12243), .B1(n13585), .B2(n12237), .ZN(
        n4109) );
  AOI221_X1 U2916 ( .B1(n12159), .B2(n14135), .C1(n12153), .C2(n14201), .A(
        n4117), .ZN(n4110) );
  OAI22_X1 U2917 ( .A1(n13950), .A2(n12147), .B1(n13792), .B2(n12141), .ZN(
        n4117) );
  AOI221_X1 U2918 ( .B1(n12255), .B2(n11721), .C1(n12249), .C2(n11541), .A(
        n4090), .ZN(n4083) );
  OAI22_X1 U2919 ( .A1(n14343), .A2(n12243), .B1(n13584), .B2(n12237), .ZN(
        n4090) );
  AOI221_X1 U2920 ( .B1(n12159), .B2(n14134), .C1(n12153), .C2(n14200), .A(
        n4098), .ZN(n4091) );
  OAI22_X1 U2921 ( .A1(n13949), .A2(n12147), .B1(n13791), .B2(n12141), .ZN(
        n4098) );
  AOI221_X1 U2922 ( .B1(n12255), .B2(n11722), .C1(n12249), .C2(n11542), .A(
        n4071), .ZN(n4064) );
  OAI22_X1 U2923 ( .A1(n14342), .A2(n12243), .B1(n13583), .B2(n12237), .ZN(
        n4071) );
  AOI221_X1 U2924 ( .B1(n12159), .B2(n14133), .C1(n12153), .C2(n14199), .A(
        n4079), .ZN(n4072) );
  OAI22_X1 U2925 ( .A1(n13948), .A2(n12147), .B1(n13790), .B2(n12141), .ZN(
        n4079) );
  AOI221_X1 U2926 ( .B1(n12255), .B2(n11723), .C1(n12249), .C2(n11543), .A(
        n4052), .ZN(n4045) );
  OAI22_X1 U2927 ( .A1(n14341), .A2(n12243), .B1(n13582), .B2(n12237), .ZN(
        n4052) );
  AOI221_X1 U2928 ( .B1(n12159), .B2(n14132), .C1(n12153), .C2(n14198), .A(
        n4060), .ZN(n4053) );
  OAI22_X1 U2929 ( .A1(n13947), .A2(n12147), .B1(n13789), .B2(n12141), .ZN(
        n4060) );
  AOI221_X1 U2930 ( .B1(n12255), .B2(n11724), .C1(n12249), .C2(n11544), .A(
        n4033), .ZN(n4026) );
  OAI22_X1 U2931 ( .A1(n13645), .A2(n12243), .B1(n13581), .B2(n12237), .ZN(
        n4033) );
  AOI221_X1 U2932 ( .B1(n12159), .B2(n14131), .C1(n12153), .C2(n14197), .A(
        n4041), .ZN(n4034) );
  OAI22_X1 U2933 ( .A1(n13946), .A2(n12147), .B1(n13788), .B2(n12141), .ZN(
        n4041) );
  AOI221_X1 U2934 ( .B1(n12255), .B2(n11725), .C1(n12249), .C2(n11545), .A(
        n4014), .ZN(n4007) );
  OAI22_X1 U2935 ( .A1(n13644), .A2(n12243), .B1(n13580), .B2(n12237), .ZN(
        n4014) );
  AOI221_X1 U2936 ( .B1(n12159), .B2(n14130), .C1(n12153), .C2(n14196), .A(
        n4022), .ZN(n4015) );
  OAI22_X1 U2937 ( .A1(n13945), .A2(n12147), .B1(n13787), .B2(n12141), .ZN(
        n4022) );
  AOI221_X1 U2938 ( .B1(n12256), .B2(n11726), .C1(n12250), .C2(n11546), .A(
        n3995), .ZN(n3988) );
  OAI22_X1 U2939 ( .A1(n13643), .A2(n12244), .B1(n13579), .B2(n12238), .ZN(
        n3995) );
  AOI221_X1 U2940 ( .B1(n12160), .B2(n14024), .C1(n12154), .C2(n14195), .A(
        n4003), .ZN(n3996) );
  OAI22_X1 U2941 ( .A1(n13944), .A2(n12148), .B1(n13786), .B2(n12142), .ZN(
        n4003) );
  AOI221_X1 U2942 ( .B1(n12256), .B2(n11727), .C1(n12250), .C2(n11547), .A(
        n3976), .ZN(n3969) );
  OAI22_X1 U2943 ( .A1(n13642), .A2(n12244), .B1(n13578), .B2(n12238), .ZN(
        n3976) );
  AOI221_X1 U2944 ( .B1(n12160), .B2(n14023), .C1(n12154), .C2(n14194), .A(
        n3984), .ZN(n3977) );
  OAI22_X1 U2945 ( .A1(n13943), .A2(n12148), .B1(n13785), .B2(n12142), .ZN(
        n3984) );
  AOI221_X1 U2946 ( .B1(n12256), .B2(n11728), .C1(n12250), .C2(n11548), .A(
        n3957), .ZN(n3950) );
  OAI22_X1 U2947 ( .A1(n13641), .A2(n12244), .B1(n13577), .B2(n12238), .ZN(
        n3957) );
  AOI221_X1 U2948 ( .B1(n12160), .B2(n14022), .C1(n12154), .C2(n14193), .A(
        n3965), .ZN(n3958) );
  OAI22_X1 U2949 ( .A1(n13942), .A2(n12148), .B1(n13784), .B2(n12142), .ZN(
        n3965) );
  AOI221_X1 U2950 ( .B1(n12256), .B2(n11729), .C1(n12250), .C2(n11549), .A(
        n3938), .ZN(n3931) );
  OAI22_X1 U2951 ( .A1(n13640), .A2(n12244), .B1(n13576), .B2(n12238), .ZN(
        n3938) );
  AOI221_X1 U2952 ( .B1(n12160), .B2(n14021), .C1(n12154), .C2(n14192), .A(
        n3946), .ZN(n3939) );
  OAI22_X1 U2953 ( .A1(n13941), .A2(n12148), .B1(n13783), .B2(n12142), .ZN(
        n3946) );
  AOI221_X1 U2954 ( .B1(n12256), .B2(n11730), .C1(n12250), .C2(n11550), .A(
        n3919), .ZN(n3912) );
  OAI22_X1 U2955 ( .A1(n13639), .A2(n12244), .B1(n13575), .B2(n12238), .ZN(
        n3919) );
  AOI221_X1 U2956 ( .B1(n12160), .B2(n14020), .C1(n12154), .C2(n14191), .A(
        n3927), .ZN(n3920) );
  OAI22_X1 U2957 ( .A1(n13940), .A2(n12148), .B1(n13782), .B2(n12142), .ZN(
        n3927) );
  AOI221_X1 U2958 ( .B1(n12256), .B2(n11731), .C1(n12250), .C2(n11551), .A(
        n3900), .ZN(n3893) );
  OAI22_X1 U2959 ( .A1(n13638), .A2(n12244), .B1(n13574), .B2(n12238), .ZN(
        n3900) );
  AOI221_X1 U2960 ( .B1(n12160), .B2(n14019), .C1(n12154), .C2(n14190), .A(
        n3908), .ZN(n3901) );
  OAI22_X1 U2961 ( .A1(n13939), .A2(n12148), .B1(n13781), .B2(n12142), .ZN(
        n3908) );
  AOI221_X1 U2962 ( .B1(n12256), .B2(n11732), .C1(n12250), .C2(n11552), .A(
        n3881), .ZN(n3874) );
  OAI22_X1 U2963 ( .A1(n13637), .A2(n12244), .B1(n13573), .B2(n12238), .ZN(
        n3881) );
  AOI221_X1 U2964 ( .B1(n12160), .B2(n14018), .C1(n12154), .C2(n14189), .A(
        n3889), .ZN(n3882) );
  OAI22_X1 U2965 ( .A1(n13938), .A2(n12148), .B1(n13780), .B2(n12142), .ZN(
        n3889) );
  AOI221_X1 U2966 ( .B1(n12256), .B2(n11733), .C1(n12250), .C2(n11553), .A(
        n3862), .ZN(n3855) );
  OAI22_X1 U2967 ( .A1(n13636), .A2(n12244), .B1(n13572), .B2(n12238), .ZN(
        n3862) );
  AOI221_X1 U2968 ( .B1(n12160), .B2(n14017), .C1(n12154), .C2(n14188), .A(
        n3870), .ZN(n3863) );
  OAI22_X1 U2969 ( .A1(n13937), .A2(n12148), .B1(n13779), .B2(n12142), .ZN(
        n3870) );
  AOI221_X1 U2970 ( .B1(n12256), .B2(n11734), .C1(n12250), .C2(n11554), .A(
        n3843), .ZN(n3836) );
  OAI22_X1 U2971 ( .A1(n13635), .A2(n12244), .B1(n13571), .B2(n12238), .ZN(
        n3843) );
  AOI221_X1 U2972 ( .B1(n12160), .B2(n14016), .C1(n12154), .C2(n14187), .A(
        n3851), .ZN(n3844) );
  OAI22_X1 U2973 ( .A1(n13936), .A2(n12148), .B1(n13778), .B2(n12142), .ZN(
        n3851) );
  AOI221_X1 U2974 ( .B1(n12256), .B2(n11735), .C1(n12250), .C2(n11555), .A(
        n3824), .ZN(n3817) );
  OAI22_X1 U2975 ( .A1(n13634), .A2(n12244), .B1(n13570), .B2(n12238), .ZN(
        n3824) );
  AOI221_X1 U2976 ( .B1(n12160), .B2(n14015), .C1(n12154), .C2(n14186), .A(
        n3832), .ZN(n3825) );
  OAI22_X1 U2977 ( .A1(n13935), .A2(n12148), .B1(n13777), .B2(n12142), .ZN(
        n3832) );
  AOI221_X1 U2978 ( .B1(n12256), .B2(n11736), .C1(n12250), .C2(n11556), .A(
        n3805), .ZN(n3798) );
  OAI22_X1 U2979 ( .A1(n13633), .A2(n12244), .B1(n13569), .B2(n12238), .ZN(
        n3805) );
  AOI221_X1 U2980 ( .B1(n12160), .B2(n14014), .C1(n12154), .C2(n14185), .A(
        n3813), .ZN(n3806) );
  OAI22_X1 U2981 ( .A1(n13934), .A2(n12148), .B1(n13776), .B2(n12142), .ZN(
        n3813) );
  AOI221_X1 U2982 ( .B1(n12256), .B2(n11737), .C1(n12250), .C2(n11557), .A(
        n3786), .ZN(n3779) );
  OAI22_X1 U2983 ( .A1(n13632), .A2(n12244), .B1(n13568), .B2(n12238), .ZN(
        n3786) );
  AOI221_X1 U2984 ( .B1(n12160), .B2(n14013), .C1(n12154), .C2(n14184), .A(
        n3794), .ZN(n3787) );
  OAI22_X1 U2985 ( .A1(n13933), .A2(n12148), .B1(n13775), .B2(n12142), .ZN(
        n3794) );
  AOI221_X1 U2986 ( .B1(n12257), .B2(n11738), .C1(n12251), .C2(n11558), .A(
        n3767), .ZN(n3760) );
  OAI22_X1 U2987 ( .A1(n13631), .A2(n12245), .B1(n13567), .B2(n12239), .ZN(
        n3767) );
  AOI221_X1 U2988 ( .B1(n12161), .B2(n14012), .C1(n12155), .C2(n14183), .A(
        n3775), .ZN(n3768) );
  OAI22_X1 U2989 ( .A1(n13932), .A2(n12149), .B1(n13774), .B2(n12143), .ZN(
        n3775) );
  AOI221_X1 U2990 ( .B1(n12257), .B2(n11739), .C1(n12251), .C2(n11559), .A(
        n3748), .ZN(n3741) );
  OAI22_X1 U2991 ( .A1(n13630), .A2(n12245), .B1(n13566), .B2(n12239), .ZN(
        n3748) );
  AOI221_X1 U2992 ( .B1(n12161), .B2(n14011), .C1(n12155), .C2(n14182), .A(
        n3756), .ZN(n3749) );
  OAI22_X1 U2993 ( .A1(n13931), .A2(n12149), .B1(n13773), .B2(n12143), .ZN(
        n3756) );
  AOI221_X1 U2994 ( .B1(n12257), .B2(n11740), .C1(n12251), .C2(n11560), .A(
        n3729), .ZN(n3722) );
  OAI22_X1 U2995 ( .A1(n13629), .A2(n12245), .B1(n13565), .B2(n12239), .ZN(
        n3729) );
  AOI221_X1 U2996 ( .B1(n12161), .B2(n14010), .C1(n12155), .C2(n14181), .A(
        n3737), .ZN(n3730) );
  OAI22_X1 U2997 ( .A1(n13930), .A2(n12149), .B1(n13772), .B2(n12143), .ZN(
        n3737) );
  AOI221_X1 U2998 ( .B1(n12257), .B2(n11741), .C1(n12251), .C2(n11561), .A(
        n3710), .ZN(n3703) );
  OAI22_X1 U2999 ( .A1(n13628), .A2(n12245), .B1(n13564), .B2(n12239), .ZN(
        n3710) );
  AOI221_X1 U3000 ( .B1(n12161), .B2(n14009), .C1(n12155), .C2(n14180), .A(
        n3718), .ZN(n3711) );
  OAI22_X1 U3001 ( .A1(n13929), .A2(n12149), .B1(n13771), .B2(n12143), .ZN(
        n3718) );
  AOI221_X1 U3002 ( .B1(n12257), .B2(n11742), .C1(n12251), .C2(n11562), .A(
        n3691), .ZN(n3684) );
  OAI22_X1 U3003 ( .A1(n13627), .A2(n12245), .B1(n13563), .B2(n12239), .ZN(
        n3691) );
  AOI221_X1 U3004 ( .B1(n12161), .B2(n14008), .C1(n12155), .C2(n14179), .A(
        n3699), .ZN(n3692) );
  OAI22_X1 U3005 ( .A1(n14106), .A2(n12149), .B1(n13770), .B2(n12143), .ZN(
        n3699) );
  AOI221_X1 U3006 ( .B1(n12257), .B2(n11743), .C1(n12251), .C2(n11563), .A(
        n3672), .ZN(n3665) );
  OAI22_X1 U3007 ( .A1(n13626), .A2(n12245), .B1(n13562), .B2(n12239), .ZN(
        n3672) );
  AOI221_X1 U3008 ( .B1(n12161), .B2(n14007), .C1(n12155), .C2(n14178), .A(
        n3680), .ZN(n3673) );
  OAI22_X1 U3009 ( .A1(n14105), .A2(n12149), .B1(n13769), .B2(n12143), .ZN(
        n3680) );
  AOI221_X1 U3010 ( .B1(n12257), .B2(n11744), .C1(n12251), .C2(n11564), .A(
        n3653), .ZN(n3646) );
  OAI22_X1 U3011 ( .A1(n13625), .A2(n12245), .B1(n13561), .B2(n12239), .ZN(
        n3653) );
  AOI221_X1 U3012 ( .B1(n12161), .B2(n14006), .C1(n12155), .C2(n14177), .A(
        n3661), .ZN(n3654) );
  OAI22_X1 U3013 ( .A1(n14104), .A2(n12149), .B1(n13768), .B2(n12143), .ZN(
        n3661) );
  AOI221_X1 U3014 ( .B1(n12257), .B2(n11745), .C1(n12251), .C2(n11565), .A(
        n3634), .ZN(n3627) );
  OAI22_X1 U3015 ( .A1(n13624), .A2(n12245), .B1(n13560), .B2(n12239), .ZN(
        n3634) );
  AOI221_X1 U3016 ( .B1(n12161), .B2(n14005), .C1(n12155), .C2(n14176), .A(
        n3642), .ZN(n3635) );
  OAI22_X1 U3017 ( .A1(n14103), .A2(n12149), .B1(n13767), .B2(n12143), .ZN(
        n3642) );
  AOI221_X1 U3018 ( .B1(n12257), .B2(n11746), .C1(n12251), .C2(n11566), .A(
        n3615), .ZN(n3608) );
  OAI22_X1 U3019 ( .A1(n13623), .A2(n12245), .B1(n13559), .B2(n12239), .ZN(
        n3615) );
  AOI221_X1 U3020 ( .B1(n12161), .B2(n14004), .C1(n12155), .C2(n14175), .A(
        n3623), .ZN(n3616) );
  OAI22_X1 U3021 ( .A1(n14102), .A2(n12149), .B1(n13766), .B2(n12143), .ZN(
        n3623) );
  AOI221_X1 U3022 ( .B1(n12257), .B2(n11747), .C1(n12251), .C2(n11567), .A(
        n3596), .ZN(n3589) );
  OAI22_X1 U3023 ( .A1(n13622), .A2(n12245), .B1(n13558), .B2(n12239), .ZN(
        n3596) );
  AOI221_X1 U3024 ( .B1(n12161), .B2(n14003), .C1(n12155), .C2(n14174), .A(
        n3604), .ZN(n3597) );
  OAI22_X1 U3025 ( .A1(n14101), .A2(n12149), .B1(n13765), .B2(n12143), .ZN(
        n3604) );
  AOI221_X1 U3026 ( .B1(n12257), .B2(n11748), .C1(n12251), .C2(n11568), .A(
        n3577), .ZN(n3570) );
  OAI22_X1 U3027 ( .A1(n13621), .A2(n12245), .B1(n13557), .B2(n12239), .ZN(
        n3577) );
  AOI221_X1 U3028 ( .B1(n12161), .B2(n14002), .C1(n12155), .C2(n14173), .A(
        n3585), .ZN(n3578) );
  OAI22_X1 U3029 ( .A1(n14100), .A2(n12149), .B1(n13764), .B2(n12143), .ZN(
        n3585) );
  AOI221_X1 U3030 ( .B1(n12257), .B2(n11749), .C1(n12251), .C2(n11569), .A(
        n3558), .ZN(n3551) );
  OAI22_X1 U3031 ( .A1(n13620), .A2(n12245), .B1(n13556), .B2(n12239), .ZN(
        n3558) );
  AOI221_X1 U3032 ( .B1(n12161), .B2(n14001), .C1(n12155), .C2(n14172), .A(
        n3566), .ZN(n3559) );
  OAI22_X1 U3033 ( .A1(n14099), .A2(n12149), .B1(n13763), .B2(n12143), .ZN(
        n3566) );
  AOI221_X1 U3034 ( .B1(n12258), .B2(n11750), .C1(n12252), .C2(n11570), .A(
        n3539), .ZN(n3532) );
  OAI22_X1 U3035 ( .A1(n13619), .A2(n12246), .B1(n13555), .B2(n12240), .ZN(
        n3539) );
  AOI221_X1 U3036 ( .B1(n12162), .B2(n14000), .C1(n12156), .C2(n14171), .A(
        n3547), .ZN(n3540) );
  OAI22_X1 U3037 ( .A1(n14098), .A2(n12150), .B1(n13762), .B2(n12144), .ZN(
        n3547) );
  AOI221_X1 U3038 ( .B1(n12258), .B2(n11751), .C1(n12252), .C2(n11571), .A(
        n3520), .ZN(n3513) );
  OAI22_X1 U3039 ( .A1(n13618), .A2(n12246), .B1(n13554), .B2(n12240), .ZN(
        n3520) );
  AOI221_X1 U3040 ( .B1(n12162), .B2(n13999), .C1(n12156), .C2(n14170), .A(
        n3528), .ZN(n3521) );
  OAI22_X1 U3041 ( .A1(n14097), .A2(n12150), .B1(n13761), .B2(n12144), .ZN(
        n3528) );
  AOI221_X1 U3042 ( .B1(n12258), .B2(n11752), .C1(n12252), .C2(n11572), .A(
        n3501), .ZN(n3494) );
  OAI22_X1 U3043 ( .A1(n13617), .A2(n12246), .B1(n13553), .B2(n12240), .ZN(
        n3501) );
  AOI221_X1 U3044 ( .B1(n12162), .B2(n13998), .C1(n12156), .C2(n14169), .A(
        n3509), .ZN(n3502) );
  OAI22_X1 U3045 ( .A1(n14096), .A2(n12150), .B1(n13760), .B2(n12144), .ZN(
        n3509) );
  AOI221_X1 U3046 ( .B1(n12258), .B2(n11753), .C1(n12252), .C2(n11573), .A(
        n3482), .ZN(n3475) );
  OAI22_X1 U3047 ( .A1(n13616), .A2(n12246), .B1(n13552), .B2(n12240), .ZN(
        n3482) );
  AOI221_X1 U3048 ( .B1(n12162), .B2(n13997), .C1(n12156), .C2(n14168), .A(
        n3490), .ZN(n3483) );
  OAI22_X1 U3049 ( .A1(n14095), .A2(n12150), .B1(n13759), .B2(n12144), .ZN(
        n3490) );
  AOI221_X1 U3050 ( .B1(n12258), .B2(n11754), .C1(n12252), .C2(n11574), .A(
        n3463), .ZN(n3456) );
  OAI22_X1 U3051 ( .A1(n13615), .A2(n12246), .B1(n13551), .B2(n12240), .ZN(
        n3463) );
  AOI221_X1 U3052 ( .B1(n12162), .B2(n13996), .C1(n12156), .C2(n14167), .A(
        n3471), .ZN(n3464) );
  OAI22_X1 U3053 ( .A1(n14094), .A2(n12150), .B1(n13758), .B2(n12144), .ZN(
        n3471) );
  AOI221_X1 U3054 ( .B1(n12258), .B2(n11755), .C1(n12252), .C2(n11575), .A(
        n3444), .ZN(n3437) );
  OAI22_X1 U3055 ( .A1(n13614), .A2(n12246), .B1(n13550), .B2(n12240), .ZN(
        n3444) );
  AOI221_X1 U3056 ( .B1(n12162), .B2(n13995), .C1(n12156), .C2(n14166), .A(
        n3452), .ZN(n3445) );
  OAI22_X1 U3057 ( .A1(n14093), .A2(n12150), .B1(n13757), .B2(n12144), .ZN(
        n3452) );
  AOI221_X1 U3058 ( .B1(n12258), .B2(n11756), .C1(n12252), .C2(n11576), .A(
        n3425), .ZN(n3418) );
  OAI22_X1 U3059 ( .A1(n13613), .A2(n12246), .B1(n13549), .B2(n12240), .ZN(
        n3425) );
  AOI221_X1 U3060 ( .B1(n12162), .B2(n13994), .C1(n12156), .C2(n14165), .A(
        n3433), .ZN(n3426) );
  OAI22_X1 U3061 ( .A1(n14092), .A2(n12150), .B1(n13756), .B2(n12144), .ZN(
        n3433) );
  AOI221_X1 U3062 ( .B1(n12258), .B2(n11757), .C1(n12252), .C2(n11577), .A(
        n3406), .ZN(n3399) );
  OAI22_X1 U3063 ( .A1(n13612), .A2(n12246), .B1(n13548), .B2(n12240), .ZN(
        n3406) );
  AOI221_X1 U3064 ( .B1(n12162), .B2(n13993), .C1(n12156), .C2(n14164), .A(
        n3414), .ZN(n3407) );
  OAI22_X1 U3065 ( .A1(n14091), .A2(n12150), .B1(n13755), .B2(n12144), .ZN(
        n3414) );
  AOI221_X1 U3066 ( .B1(n12258), .B2(n11758), .C1(n12252), .C2(n11578), .A(
        n3387), .ZN(n3380) );
  OAI22_X1 U3067 ( .A1(n13611), .A2(n12246), .B1(n13547), .B2(n12240), .ZN(
        n3387) );
  AOI221_X1 U3068 ( .B1(n12162), .B2(n13992), .C1(n12156), .C2(n14163), .A(
        n3395), .ZN(n3388) );
  OAI22_X1 U3069 ( .A1(n14090), .A2(n12150), .B1(n13754), .B2(n12144), .ZN(
        n3395) );
  AOI221_X1 U3070 ( .B1(n12258), .B2(n11759), .C1(n12252), .C2(n11579), .A(
        n3368), .ZN(n3361) );
  OAI22_X1 U3071 ( .A1(n13610), .A2(n12246), .B1(n13546), .B2(n12240), .ZN(
        n3368) );
  AOI221_X1 U3072 ( .B1(n12162), .B2(n13991), .C1(n12156), .C2(n14162), .A(
        n3376), .ZN(n3369) );
  OAI22_X1 U3073 ( .A1(n14089), .A2(n12150), .B1(n13753), .B2(n12144), .ZN(
        n3376) );
  AOI221_X1 U3074 ( .B1(n12258), .B2(n11760), .C1(n12252), .C2(n11580), .A(
        n3349), .ZN(n3342) );
  OAI22_X1 U3075 ( .A1(n13609), .A2(n12246), .B1(n13545), .B2(n12240), .ZN(
        n3349) );
  AOI221_X1 U3076 ( .B1(n12162), .B2(n13990), .C1(n12156), .C2(n14161), .A(
        n3357), .ZN(n3350) );
  OAI22_X1 U3077 ( .A1(n14088), .A2(n12150), .B1(n13752), .B2(n12144), .ZN(
        n3357) );
  AOI221_X1 U3078 ( .B1(n12258), .B2(n11761), .C1(n12252), .C2(n11581), .A(
        n3330), .ZN(n3323) );
  OAI22_X1 U3079 ( .A1(n13608), .A2(n12246), .B1(n13544), .B2(n12240), .ZN(
        n3330) );
  AOI221_X1 U3080 ( .B1(n12162), .B2(n13989), .C1(n12156), .C2(n14160), .A(
        n3338), .ZN(n3331) );
  OAI22_X1 U3081 ( .A1(n14087), .A2(n12150), .B1(n13751), .B2(n12144), .ZN(
        n3338) );
  AOI221_X1 U3082 ( .B1(n12163), .B2(n13827), .C1(n12157), .C2(n14159), .A(
        n3319), .ZN(n3312) );
  OAI22_X1 U3083 ( .A1(n14086), .A2(n12151), .B1(n13750), .B2(n12145), .ZN(
        n3319) );
  AOI221_X1 U3084 ( .B1(n12259), .B2(n13864), .C1(n12253), .C2(n13868), .A(
        n3311), .ZN(n3304) );
  OAI22_X1 U3085 ( .A1(n13607), .A2(n12247), .B1(n13543), .B2(n12241), .ZN(
        n3311) );
  AOI221_X1 U3086 ( .B1(n12163), .B2(n13826), .C1(n12157), .C2(n14158), .A(
        n3300), .ZN(n3293) );
  OAI22_X1 U3087 ( .A1(n14085), .A2(n12151), .B1(n13749), .B2(n12145), .ZN(
        n3300) );
  AOI221_X1 U3088 ( .B1(n12259), .B2(n13863), .C1(n12253), .C2(n13867), .A(
        n3292), .ZN(n3285) );
  OAI22_X1 U3089 ( .A1(n13606), .A2(n12247), .B1(n13542), .B2(n12241), .ZN(
        n3292) );
  AOI221_X1 U3090 ( .B1(n12163), .B2(n13825), .C1(n12157), .C2(n14157), .A(
        n3281), .ZN(n3274) );
  OAI22_X1 U3091 ( .A1(n14084), .A2(n12151), .B1(n13748), .B2(n12145), .ZN(
        n3281) );
  AOI221_X1 U3092 ( .B1(n12259), .B2(n13862), .C1(n12253), .C2(n13866), .A(
        n3273), .ZN(n3266) );
  OAI22_X1 U3093 ( .A1(n13605), .A2(n12247), .B1(n13541), .B2(n12241), .ZN(
        n3273) );
  AOI221_X1 U3094 ( .B1(n12163), .B2(n13824), .C1(n12157), .C2(n14156), .A(
        n3260), .ZN(n3239) );
  OAI22_X1 U3095 ( .A1(n14083), .A2(n12151), .B1(n13747), .B2(n12145), .ZN(
        n3260) );
  AOI221_X1 U3096 ( .B1(n12259), .B2(n13861), .C1(n12253), .C2(n13865), .A(
        n3236), .ZN(n3215) );
  OAI22_X1 U3097 ( .A1(n13604), .A2(n12247), .B1(n13540), .B2(n12241), .ZN(
        n3236) );
  NAND2_X1 U3098 ( .A1(n4450), .A2(n4466), .ZN(n3246) );
  NAND2_X1 U3099 ( .A1(n4450), .A2(n4465), .ZN(n3247) );
  NAND2_X1 U3100 ( .A1(n4454), .A2(n4466), .ZN(n3251) );
  NAND2_X1 U3101 ( .A1(n4454), .A2(n4465), .ZN(n3252) );
  AOI221_X1 U3102 ( .B1(n12302), .B2(n11762), .C1(n12296), .C2(n11582), .A(
        n4430), .ZN(n4427) );
  OAI22_X1 U3103 ( .A1(n14408), .A2(n12290), .B1(n14385), .B2(n12284), .ZN(
        n4430) );
  AOI221_X1 U3104 ( .B1(n12302), .B2(n11763), .C1(n12296), .C2(n11583), .A(
        n4354), .ZN(n4351) );
  OAI22_X1 U3105 ( .A1(n14404), .A2(n12290), .B1(n14381), .B2(n12284), .ZN(
        n4354) );
  AOI221_X1 U3106 ( .B1(n12302), .B2(n11764), .C1(n12296), .C2(n11584), .A(
        n4335), .ZN(n4332) );
  OAI22_X1 U3107 ( .A1(n14403), .A2(n12290), .B1(n14380), .B2(n12284), .ZN(
        n4335) );
  AOI221_X1 U3108 ( .B1(n12306), .B2(n11765), .C1(n12300), .C2(n11585), .A(
        n3328), .ZN(n3325) );
  OAI22_X1 U3109 ( .A1(n14253), .A2(n12294), .B1(n14217), .B2(n12288), .ZN(
        n3328) );
  BUF_X1 U3110 ( .A(n1892), .Z(n13210) );
  BUF_X1 U3111 ( .A(n1891), .Z(n13213) );
  BUF_X1 U3112 ( .A(n1890), .Z(n13216) );
  BUF_X1 U3113 ( .A(n1889), .Z(n13219) );
  BUF_X1 U3114 ( .A(n1888), .Z(n13222) );
  BUF_X1 U3115 ( .A(n1887), .Z(n13225) );
  BUF_X1 U3116 ( .A(n1881), .Z(n13243) );
  BUF_X1 U3117 ( .A(n1880), .Z(n13246) );
  BUF_X1 U3118 ( .A(n1879), .Z(n13249) );
  BUF_X1 U3119 ( .A(n1878), .Z(n13252) );
  BUF_X1 U3120 ( .A(n1877), .Z(n13255) );
  BUF_X1 U3121 ( .A(n1876), .Z(n13258) );
  BUF_X1 U3122 ( .A(n1875), .Z(n13261) );
  BUF_X1 U3123 ( .A(n1874), .Z(n13264) );
  BUF_X1 U3124 ( .A(n1873), .Z(n13267) );
  BUF_X1 U3125 ( .A(n1872), .Z(n13270) );
  BUF_X1 U3126 ( .A(n1871), .Z(n13273) );
  BUF_X1 U3127 ( .A(n1870), .Z(n13276) );
  BUF_X1 U3128 ( .A(n1869), .Z(n13279) );
  BUF_X1 U3129 ( .A(n1868), .Z(n13282) );
  BUF_X1 U3130 ( .A(n1867), .Z(n13285) );
  BUF_X1 U3131 ( .A(n1866), .Z(n13288) );
  BUF_X1 U3132 ( .A(n1865), .Z(n13291) );
  BUF_X1 U3133 ( .A(n1864), .Z(n13294) );
  BUF_X1 U3134 ( .A(n1863), .Z(n13297) );
  BUF_X1 U3135 ( .A(n1862), .Z(n13300) );
  BUF_X1 U3136 ( .A(n1861), .Z(n13303) );
  BUF_X1 U3137 ( .A(n1860), .Z(n13306) );
  BUF_X1 U3138 ( .A(n1859), .Z(n13309) );
  BUF_X1 U3139 ( .A(n1858), .Z(n13312) );
  BUF_X1 U3140 ( .A(n1857), .Z(n13315) );
  BUF_X1 U3141 ( .A(n1856), .Z(n13318) );
  BUF_X1 U3142 ( .A(n1855), .Z(n13321) );
  BUF_X1 U3143 ( .A(n1854), .Z(n13324) );
  BUF_X1 U3144 ( .A(n1853), .Z(n13327) );
  BUF_X1 U3145 ( .A(n1852), .Z(n13330) );
  BUF_X1 U3146 ( .A(n1851), .Z(n13333) );
  BUF_X1 U3147 ( .A(n1850), .Z(n13336) );
  BUF_X1 U3148 ( .A(n1849), .Z(n13339) );
  BUF_X1 U3149 ( .A(n1848), .Z(n13342) );
  BUF_X1 U3150 ( .A(n1847), .Z(n13345) );
  BUF_X1 U3151 ( .A(n1846), .Z(n13348) );
  BUF_X1 U3152 ( .A(n1845), .Z(n13351) );
  BUF_X1 U3153 ( .A(n1844), .Z(n13354) );
  BUF_X1 U3154 ( .A(n1843), .Z(n13357) );
  BUF_X1 U3155 ( .A(n1841), .Z(n13380) );
  BUF_X1 U3156 ( .A(n1876), .Z(n13257) );
  BUF_X1 U3157 ( .A(n1875), .Z(n13260) );
  BUF_X1 U3158 ( .A(n1874), .Z(n13263) );
  BUF_X1 U3159 ( .A(n1873), .Z(n13266) );
  BUF_X1 U3160 ( .A(n1872), .Z(n13269) );
  BUF_X1 U3161 ( .A(n1871), .Z(n13272) );
  BUF_X1 U3162 ( .A(n1870), .Z(n13275) );
  BUF_X1 U3163 ( .A(n1869), .Z(n13278) );
  BUF_X1 U3164 ( .A(n1868), .Z(n13281) );
  BUF_X1 U3165 ( .A(n1867), .Z(n13284) );
  BUF_X1 U3166 ( .A(n1866), .Z(n13287) );
  BUF_X1 U3167 ( .A(n1865), .Z(n13290) );
  BUF_X1 U3168 ( .A(n1864), .Z(n13293) );
  BUF_X1 U3169 ( .A(n1863), .Z(n13296) );
  BUF_X1 U3170 ( .A(n1862), .Z(n13299) );
  BUF_X1 U3171 ( .A(n1861), .Z(n13302) );
  BUF_X1 U3172 ( .A(n1860), .Z(n13305) );
  BUF_X1 U3173 ( .A(n1850), .Z(n13335) );
  BUF_X1 U3174 ( .A(n1849), .Z(n13338) );
  BUF_X1 U3175 ( .A(n1848), .Z(n13341) );
  BUF_X1 U3176 ( .A(n1847), .Z(n13344) );
  BUF_X1 U3177 ( .A(n1846), .Z(n13347) );
  BUF_X1 U3178 ( .A(n1845), .Z(n13350) );
  BUF_X1 U3179 ( .A(n1844), .Z(n13353) );
  BUF_X1 U3180 ( .A(n1843), .Z(n13356) );
  BUF_X1 U3181 ( .A(n1893), .Z(n13206) );
  BUF_X1 U3182 ( .A(n1892), .Z(n13209) );
  BUF_X1 U3183 ( .A(n1891), .Z(n13212) );
  BUF_X1 U3184 ( .A(n1890), .Z(n13215) );
  BUF_X1 U3185 ( .A(n1889), .Z(n13218) );
  BUF_X1 U3186 ( .A(n1888), .Z(n13221) );
  BUF_X1 U3187 ( .A(n1887), .Z(n13224) );
  BUF_X1 U3188 ( .A(n1886), .Z(n13227) );
  BUF_X1 U3189 ( .A(n1885), .Z(n13230) );
  BUF_X1 U3190 ( .A(n1884), .Z(n13233) );
  BUF_X1 U3191 ( .A(n1883), .Z(n13236) );
  BUF_X1 U3192 ( .A(n1882), .Z(n13239) );
  BUF_X1 U3193 ( .A(n1881), .Z(n13242) );
  BUF_X1 U3194 ( .A(n1880), .Z(n13245) );
  BUF_X1 U3195 ( .A(n1879), .Z(n13248) );
  BUF_X1 U3196 ( .A(n1878), .Z(n13251) );
  BUF_X1 U3197 ( .A(n1877), .Z(n13254) );
  BUF_X1 U3198 ( .A(n1859), .Z(n13308) );
  BUF_X1 U3199 ( .A(n1858), .Z(n13311) );
  BUF_X1 U3200 ( .A(n1857), .Z(n13314) );
  BUF_X1 U3201 ( .A(n1856), .Z(n13317) );
  BUF_X1 U3202 ( .A(n1855), .Z(n13320) );
  BUF_X1 U3203 ( .A(n1854), .Z(n13323) );
  BUF_X1 U3204 ( .A(n1853), .Z(n13326) );
  BUF_X1 U3205 ( .A(n1852), .Z(n13329) );
  BUF_X1 U3206 ( .A(n1851), .Z(n13332) );
  BUF_X1 U3207 ( .A(n1841), .Z(n13379) );
  NAND2_X1 U3208 ( .A1(n4469), .A2(n4450), .ZN(n3257) );
  NAND2_X1 U3209 ( .A1(n4470), .A2(n4450), .ZN(n3256) );
  NAND2_X1 U3210 ( .A1(n4449), .A2(n4450), .ZN(n3223) );
  NAND2_X1 U3211 ( .A1(n4451), .A2(n4450), .ZN(n3222) );
  NAND2_X1 U3212 ( .A1(n4469), .A2(n4454), .ZN(n3262) );
  NAND2_X1 U3213 ( .A1(n4470), .A2(n4454), .ZN(n3261) );
  NAND2_X1 U3214 ( .A1(n4449), .A2(n4454), .ZN(n3228) );
  NAND2_X1 U3215 ( .A1(n4451), .A2(n4454), .ZN(n3227) );
  NAND2_X1 U3216 ( .A1(n4458), .A2(n4452), .ZN(n3232) );
  NAND2_X1 U3217 ( .A1(n4457), .A2(n4452), .ZN(n3233) );
  NAND2_X1 U3218 ( .A1(n4458), .A2(n4455), .ZN(n3237) );
  NAND2_X1 U3219 ( .A1(n4457), .A2(n4455), .ZN(n3238) );
  BUF_X1 U3220 ( .A(n1905), .Z(n13171) );
  BUF_X1 U3221 ( .A(n1904), .Z(n13174) );
  BUF_X1 U3222 ( .A(n1903), .Z(n13177) );
  BUF_X1 U3223 ( .A(n1902), .Z(n13180) );
  BUF_X1 U3224 ( .A(n1901), .Z(n13183) );
  BUF_X1 U3225 ( .A(n1900), .Z(n13186) );
  BUF_X1 U3226 ( .A(n1893), .Z(n13207) );
  BUF_X1 U3227 ( .A(n1886), .Z(n13228) );
  BUF_X1 U3228 ( .A(n1885), .Z(n13231) );
  BUF_X1 U3229 ( .A(n1884), .Z(n13234) );
  BUF_X1 U3230 ( .A(n1883), .Z(n13237) );
  BUF_X1 U3231 ( .A(n1882), .Z(n13240) );
  BUF_X1 U3232 ( .A(n1899), .Z(n13189) );
  BUF_X1 U3233 ( .A(n1898), .Z(n13192) );
  BUF_X1 U3234 ( .A(n1897), .Z(n13195) );
  BUF_X1 U3235 ( .A(n1896), .Z(n13198) );
  BUF_X1 U3236 ( .A(n1895), .Z(n13201) );
  BUF_X1 U3237 ( .A(n1894), .Z(n13204) );
  BUF_X1 U3238 ( .A(n1905), .Z(n13172) );
  BUF_X1 U3239 ( .A(n1904), .Z(n13175) );
  BUF_X1 U3240 ( .A(n1903), .Z(n13178) );
  BUF_X1 U3241 ( .A(n1902), .Z(n13181) );
  BUF_X1 U3242 ( .A(n1901), .Z(n13184) );
  BUF_X1 U3243 ( .A(n1900), .Z(n13187) );
  BUF_X1 U3244 ( .A(n1899), .Z(n13190) );
  BUF_X1 U3245 ( .A(n1898), .Z(n13193) );
  BUF_X1 U3246 ( .A(n1897), .Z(n13196) );
  BUF_X1 U3247 ( .A(n1896), .Z(n13199) );
  BUF_X1 U3248 ( .A(n1895), .Z(n13202) );
  BUF_X1 U3249 ( .A(n1894), .Z(n13205) );
  BUF_X1 U3250 ( .A(n1893), .Z(n13208) );
  BUF_X1 U3251 ( .A(n1892), .Z(n13211) );
  BUF_X1 U3252 ( .A(n1891), .Z(n13214) );
  BUF_X1 U3253 ( .A(n1890), .Z(n13217) );
  BUF_X1 U3254 ( .A(n1889), .Z(n13220) );
  BUF_X1 U3255 ( .A(n1888), .Z(n13223) );
  BUF_X1 U3256 ( .A(n1887), .Z(n13226) );
  BUF_X1 U3257 ( .A(n1886), .Z(n13229) );
  BUF_X1 U3258 ( .A(n1885), .Z(n13232) );
  BUF_X1 U3259 ( .A(n1884), .Z(n13235) );
  BUF_X1 U3260 ( .A(n1883), .Z(n13238) );
  BUF_X1 U3261 ( .A(n1882), .Z(n13241) );
  BUF_X1 U3262 ( .A(n1881), .Z(n13244) );
  BUF_X1 U3263 ( .A(n1880), .Z(n13247) );
  BUF_X1 U3264 ( .A(n1879), .Z(n13250) );
  BUF_X1 U3265 ( .A(n1878), .Z(n13253) );
  BUF_X1 U3266 ( .A(n1877), .Z(n13256) );
  BUF_X1 U3267 ( .A(n1876), .Z(n13259) );
  BUF_X1 U3268 ( .A(n1875), .Z(n13262) );
  BUF_X1 U3269 ( .A(n1874), .Z(n13265) );
  BUF_X1 U3270 ( .A(n1873), .Z(n13268) );
  BUF_X1 U3271 ( .A(n1872), .Z(n13271) );
  BUF_X1 U3272 ( .A(n1871), .Z(n13274) );
  BUF_X1 U3273 ( .A(n1870), .Z(n13277) );
  BUF_X1 U3274 ( .A(n1869), .Z(n13280) );
  BUF_X1 U3275 ( .A(n1868), .Z(n13283) );
  BUF_X1 U3276 ( .A(n1867), .Z(n13286) );
  BUF_X1 U3277 ( .A(n1866), .Z(n13289) );
  BUF_X1 U3278 ( .A(n1865), .Z(n13292) );
  BUF_X1 U3279 ( .A(n1864), .Z(n13295) );
  BUF_X1 U3280 ( .A(n1863), .Z(n13298) );
  BUF_X1 U3281 ( .A(n1862), .Z(n13301) );
  BUF_X1 U3282 ( .A(n1861), .Z(n13304) );
  BUF_X1 U3283 ( .A(n1860), .Z(n13307) );
  BUF_X1 U3284 ( .A(n1859), .Z(n13310) );
  BUF_X1 U3285 ( .A(n1858), .Z(n13313) );
  BUF_X1 U3286 ( .A(n1857), .Z(n13316) );
  BUF_X1 U3287 ( .A(n1856), .Z(n13319) );
  BUF_X1 U3288 ( .A(n1855), .Z(n13322) );
  BUF_X1 U3289 ( .A(n1854), .Z(n13325) );
  BUF_X1 U3290 ( .A(n1853), .Z(n13328) );
  BUF_X1 U3291 ( .A(n1852), .Z(n13331) );
  BUF_X1 U3292 ( .A(n1851), .Z(n13334) );
  BUF_X1 U3293 ( .A(n1850), .Z(n13337) );
  BUF_X1 U3294 ( .A(n1849), .Z(n13340) );
  BUF_X1 U3295 ( .A(n1848), .Z(n13343) );
  BUF_X1 U3296 ( .A(n1847), .Z(n13346) );
  BUF_X1 U3297 ( .A(n1846), .Z(n13349) );
  BUF_X1 U3298 ( .A(n1845), .Z(n13352) );
  BUF_X1 U3299 ( .A(n1844), .Z(n13355) );
  BUF_X1 U3300 ( .A(n1843), .Z(n13358) );
  BUF_X1 U3301 ( .A(n1841), .Z(n13381) );
  BUF_X1 U3302 ( .A(n1905), .Z(n13170) );
  BUF_X1 U3303 ( .A(n1904), .Z(n13173) );
  BUF_X1 U3304 ( .A(n1903), .Z(n13176) );
  BUF_X1 U3305 ( .A(n1902), .Z(n13179) );
  BUF_X1 U3306 ( .A(n1901), .Z(n13182) );
  BUF_X1 U3307 ( .A(n1900), .Z(n13185) );
  BUF_X1 U3308 ( .A(n1899), .Z(n13188) );
  BUF_X1 U3309 ( .A(n1898), .Z(n13191) );
  BUF_X1 U3310 ( .A(n1897), .Z(n13194) );
  BUF_X1 U3311 ( .A(n1896), .Z(n13197) );
  BUF_X1 U3312 ( .A(n1895), .Z(n13200) );
  BUF_X1 U3313 ( .A(n1894), .Z(n13203) );
  BUF_X1 U3314 ( .A(n3211), .Z(n12332) );
  AND2_X1 U3315 ( .A1(n4466), .A2(n4452), .ZN(n3244) );
  AND2_X1 U3316 ( .A1(n4452), .A2(n4465), .ZN(n3243) );
  AND2_X1 U3317 ( .A1(n4455), .A2(n4465), .ZN(n3248) );
  AND2_X1 U3318 ( .A1(n4455), .A2(n4466), .ZN(n3249) );
  AND2_X1 U3319 ( .A1(n4457), .A2(n4450), .ZN(n3229) );
  AND2_X1 U3320 ( .A1(n4458), .A2(n4450), .ZN(n3230) );
  AND2_X1 U3321 ( .A1(n4457), .A2(n4454), .ZN(n3234) );
  AND2_X1 U3322 ( .A1(n4458), .A2(n4454), .ZN(n3235) );
  AND2_X1 U3323 ( .A1(n4469), .A2(n4452), .ZN(n3253) );
  AND2_X1 U3324 ( .A1(n4469), .A2(n4455), .ZN(n3258) );
  AND2_X1 U3325 ( .A1(n4449), .A2(n4452), .ZN(n3219) );
  AND2_X1 U3326 ( .A1(n4451), .A2(n4452), .ZN(n3220) );
  AND2_X1 U3327 ( .A1(n4449), .A2(n4455), .ZN(n3224) );
  AND2_X1 U3328 ( .A1(n4451), .A2(n4455), .ZN(n3225) );
  AND2_X1 U3329 ( .A1(n4470), .A2(n4452), .ZN(n3254) );
  BUF_X1 U3330 ( .A(n3211), .Z(n12333) );
  BUF_X1 U3331 ( .A(n1950), .Z(n12537) );
  BUF_X1 U3332 ( .A(n1950), .Z(n12538) );
  AOI221_X1 U3333 ( .B1(n12435), .B2(n4642), .C1(n12429), .C2(n4643), .A(n3203), .ZN(n3202) );
  OAI22_X1 U3334 ( .A1(n8577), .A2(n12423), .B1(n8578), .B2(n12417), .ZN(n3203) );
  AOI221_X1 U3335 ( .B1(n12435), .B2(n4646), .C1(n12429), .C2(n4647), .A(n3176), .ZN(n3175) );
  OAI22_X1 U3336 ( .A1(n8560), .A2(n12423), .B1(n8561), .B2(n12417), .ZN(n3176) );
  AOI221_X1 U3337 ( .B1(n12435), .B2(n4652), .C1(n12429), .C2(n4653), .A(n3157), .ZN(n3156) );
  OAI22_X1 U3338 ( .A1(n8543), .A2(n12423), .B1(n8544), .B2(n12417), .ZN(n3157) );
  AOI221_X1 U3339 ( .B1(n12435), .B2(n4654), .C1(n12429), .C2(n4655), .A(n3138), .ZN(n3137) );
  OAI22_X1 U3340 ( .A1(n8526), .A2(n12423), .B1(n8527), .B2(n12417), .ZN(n3138) );
  AOI221_X1 U3341 ( .B1(n12435), .B2(n8599), .C1(n12429), .C2(n8600), .A(n3119), .ZN(n3118) );
  OAI22_X1 U3342 ( .A1(n8509), .A2(n12423), .B1(n8510), .B2(n12417), .ZN(n3119) );
  AOI221_X1 U3343 ( .B1(n12435), .B2(n8603), .C1(n12429), .C2(n8604), .A(n3100), .ZN(n3099) );
  OAI22_X1 U3344 ( .A1(n8492), .A2(n12423), .B1(n8493), .B2(n12417), .ZN(n3100) );
  AOI221_X1 U3345 ( .B1(n12435), .B2(n8611), .C1(n12429), .C2(n8612), .A(n3081), .ZN(n3080) );
  OAI22_X1 U3346 ( .A1(n8475), .A2(n12423), .B1(n8476), .B2(n12417), .ZN(n3081) );
  AOI221_X1 U3347 ( .B1(n12435), .B2(n8617), .C1(n12429), .C2(n8618), .A(n3062), .ZN(n3061) );
  OAI22_X1 U3348 ( .A1(n8458), .A2(n12423), .B1(n8459), .B2(n12417), .ZN(n3062) );
  AOI221_X1 U3349 ( .B1(n12435), .B2(n8619), .C1(n12429), .C2(n8620), .A(n3043), .ZN(n3042) );
  OAI22_X1 U3350 ( .A1(n8441), .A2(n12423), .B1(n8442), .B2(n12417), .ZN(n3043) );
  AOI221_X1 U3351 ( .B1(n12435), .B2(n8621), .C1(n12429), .C2(n8622), .A(n3024), .ZN(n3023) );
  OAI22_X1 U3352 ( .A1(n8424), .A2(n12423), .B1(n8425), .B2(n12417), .ZN(n3024) );
  AOI221_X1 U3353 ( .B1(n12435), .B2(n8623), .C1(n12429), .C2(n8624), .A(n3005), .ZN(n3004) );
  OAI22_X1 U3354 ( .A1(n8407), .A2(n12423), .B1(n8408), .B2(n12417), .ZN(n3005) );
  AOI221_X1 U3355 ( .B1(n12435), .B2(n8625), .C1(n12429), .C2(n8626), .A(n2986), .ZN(n2985) );
  OAI22_X1 U3356 ( .A1(n8390), .A2(n12423), .B1(n8391), .B2(n12417), .ZN(n2986) );
  AOI221_X1 U3357 ( .B1(n12436), .B2(n8627), .C1(n12430), .C2(n8628), .A(n2967), .ZN(n2966) );
  OAI22_X1 U3358 ( .A1(n8373), .A2(n12424), .B1(n8374), .B2(n12418), .ZN(n2967) );
  AOI221_X1 U3359 ( .B1(n12436), .B2(n8629), .C1(n12430), .C2(n8630), .A(n2948), .ZN(n2947) );
  OAI22_X1 U3360 ( .A1(n8356), .A2(n12424), .B1(n8357), .B2(n12418), .ZN(n2948) );
  AOI221_X1 U3361 ( .B1(n12436), .B2(n8631), .C1(n12430), .C2(n8632), .A(n2929), .ZN(n2928) );
  OAI22_X1 U3362 ( .A1(n8339), .A2(n12424), .B1(n8340), .B2(n12418), .ZN(n2929) );
  AOI221_X1 U3363 ( .B1(n12436), .B2(n8633), .C1(n12430), .C2(n8634), .A(n2910), .ZN(n2909) );
  OAI22_X1 U3364 ( .A1(n8322), .A2(n12424), .B1(n8323), .B2(n12418), .ZN(n2910) );
  AOI221_X1 U3365 ( .B1(n12436), .B2(n8635), .C1(n12430), .C2(n8636), .A(n2891), .ZN(n2890) );
  OAI22_X1 U3366 ( .A1(n8305), .A2(n12424), .B1(n8306), .B2(n12418), .ZN(n2891) );
  AOI221_X1 U3367 ( .B1(n12436), .B2(n8637), .C1(n12430), .C2(n8638), .A(n2872), .ZN(n2871) );
  OAI22_X1 U3368 ( .A1(n8288), .A2(n12424), .B1(n8289), .B2(n12418), .ZN(n2872) );
  AOI221_X1 U3369 ( .B1(n12436), .B2(n8639), .C1(n12430), .C2(n8640), .A(n2853), .ZN(n2852) );
  OAI22_X1 U3370 ( .A1(n8271), .A2(n12424), .B1(n8272), .B2(n12418), .ZN(n2853) );
  AOI221_X1 U3371 ( .B1(n12436), .B2(n8641), .C1(n12430), .C2(n8642), .A(n2834), .ZN(n2833) );
  OAI22_X1 U3372 ( .A1(n8254), .A2(n12424), .B1(n8255), .B2(n12418), .ZN(n2834) );
  AOI221_X1 U3373 ( .B1(n12436), .B2(n8643), .C1(n12430), .C2(n8644), .A(n2815), .ZN(n2814) );
  OAI22_X1 U3374 ( .A1(n8237), .A2(n12424), .B1(n8238), .B2(n12418), .ZN(n2815) );
  AOI221_X1 U3375 ( .B1(n12436), .B2(n8645), .C1(n12430), .C2(n8646), .A(n2796), .ZN(n2795) );
  OAI22_X1 U3376 ( .A1(n8220), .A2(n12424), .B1(n8221), .B2(n12418), .ZN(n2796) );
  AOI221_X1 U3377 ( .B1(n12436), .B2(n8647), .C1(n12430), .C2(n8648), .A(n2777), .ZN(n2776) );
  OAI22_X1 U3378 ( .A1(n8203), .A2(n12424), .B1(n8204), .B2(n12418), .ZN(n2777) );
  AOI221_X1 U3379 ( .B1(n12436), .B2(n8649), .C1(n12430), .C2(n8650), .A(n2758), .ZN(n2757) );
  OAI22_X1 U3380 ( .A1(n8186), .A2(n12424), .B1(n8187), .B2(n12418), .ZN(n2758) );
  AOI221_X1 U3381 ( .B1(n12437), .B2(n8651), .C1(n12431), .C2(n8652), .A(n2739), .ZN(n2738) );
  OAI22_X1 U3382 ( .A1(n8169), .A2(n12425), .B1(n8170), .B2(n12419), .ZN(n2739) );
  AOI221_X1 U3383 ( .B1(n12437), .B2(n8653), .C1(n12431), .C2(n8654), .A(n2720), .ZN(n2719) );
  OAI22_X1 U3384 ( .A1(n8152), .A2(n12425), .B1(n8153), .B2(n12419), .ZN(n2720) );
  AOI221_X1 U3385 ( .B1(n12437), .B2(n8655), .C1(n12431), .C2(n8656), .A(n2701), .ZN(n2700) );
  OAI22_X1 U3386 ( .A1(n8135), .A2(n12425), .B1(n8136), .B2(n12419), .ZN(n2701) );
  AOI221_X1 U3387 ( .B1(n12437), .B2(n8657), .C1(n12431), .C2(n8658), .A(n2682), .ZN(n2681) );
  OAI22_X1 U3388 ( .A1(n8118), .A2(n12425), .B1(n8119), .B2(n12419), .ZN(n2682) );
  AOI221_X1 U3389 ( .B1(n12437), .B2(n8659), .C1(n12431), .C2(n8660), .A(n2663), .ZN(n2662) );
  OAI22_X1 U3390 ( .A1(n8101), .A2(n12425), .B1(n8102), .B2(n12419), .ZN(n2663) );
  AOI221_X1 U3391 ( .B1(n12437), .B2(n8661), .C1(n12431), .C2(n8662), .A(n2644), .ZN(n2643) );
  OAI22_X1 U3392 ( .A1(n8084), .A2(n12425), .B1(n8085), .B2(n12419), .ZN(n2644) );
  AOI221_X1 U3393 ( .B1(n12437), .B2(n8663), .C1(n12431), .C2(n8664), .A(n2625), .ZN(n2624) );
  OAI22_X1 U3394 ( .A1(n8067), .A2(n12425), .B1(n8068), .B2(n12419), .ZN(n2625) );
  AOI221_X1 U3395 ( .B1(n12437), .B2(n8665), .C1(n12431), .C2(n8666), .A(n2606), .ZN(n2605) );
  OAI22_X1 U3396 ( .A1(n8050), .A2(n12425), .B1(n8051), .B2(n12419), .ZN(n2606) );
  AOI221_X1 U3397 ( .B1(n12437), .B2(n8667), .C1(n12431), .C2(n8668), .A(n2587), .ZN(n2586) );
  OAI22_X1 U3398 ( .A1(n8033), .A2(n12425), .B1(n8034), .B2(n12419), .ZN(n2587) );
  AOI221_X1 U3399 ( .B1(n12437), .B2(n8669), .C1(n12431), .C2(n8670), .A(n2568), .ZN(n2567) );
  OAI22_X1 U3400 ( .A1(n8016), .A2(n12425), .B1(n8017), .B2(n12419), .ZN(n2568) );
  AOI221_X1 U3401 ( .B1(n12437), .B2(n8671), .C1(n12431), .C2(n8672), .A(n2549), .ZN(n2548) );
  OAI22_X1 U3402 ( .A1(n7999), .A2(n12425), .B1(n8000), .B2(n12419), .ZN(n2549) );
  AOI221_X1 U3403 ( .B1(n12437), .B2(n8673), .C1(n12431), .C2(n8674), .A(n2530), .ZN(n2529) );
  OAI22_X1 U3404 ( .A1(n7982), .A2(n12425), .B1(n7983), .B2(n12419), .ZN(n2530) );
  AOI221_X1 U3405 ( .B1(n12438), .B2(n8675), .C1(n12432), .C2(n8676), .A(n2511), .ZN(n2510) );
  OAI22_X1 U3406 ( .A1(n7965), .A2(n12426), .B1(n7966), .B2(n12420), .ZN(n2511) );
  AOI221_X1 U3407 ( .B1(n12438), .B2(n8677), .C1(n12432), .C2(n8678), .A(n2492), .ZN(n2491) );
  OAI22_X1 U3408 ( .A1(n7948), .A2(n12426), .B1(n7949), .B2(n12420), .ZN(n2492) );
  AOI221_X1 U3409 ( .B1(n12438), .B2(n8679), .C1(n12432), .C2(n8680), .A(n2473), .ZN(n2472) );
  OAI22_X1 U3410 ( .A1(n7931), .A2(n12426), .B1(n7932), .B2(n12420), .ZN(n2473) );
  AOI221_X1 U3411 ( .B1(n12438), .B2(n8681), .C1(n12432), .C2(n8682), .A(n2454), .ZN(n2453) );
  OAI22_X1 U3412 ( .A1(n7914), .A2(n12426), .B1(n7915), .B2(n12420), .ZN(n2454) );
  AOI221_X1 U3413 ( .B1(n12438), .B2(n8683), .C1(n12432), .C2(n8684), .A(n2435), .ZN(n2434) );
  OAI22_X1 U3414 ( .A1(n7897), .A2(n12426), .B1(n7898), .B2(n12420), .ZN(n2435) );
  AOI221_X1 U3415 ( .B1(n12438), .B2(n8685), .C1(n12432), .C2(n8686), .A(n2416), .ZN(n2415) );
  OAI22_X1 U3416 ( .A1(n7880), .A2(n12426), .B1(n7881), .B2(n12420), .ZN(n2416) );
  AOI221_X1 U3417 ( .B1(n12438), .B2(n8687), .C1(n12432), .C2(n8688), .A(n2397), .ZN(n2396) );
  OAI22_X1 U3418 ( .A1(n7863), .A2(n12426), .B1(n7864), .B2(n12420), .ZN(n2397) );
  AOI221_X1 U3419 ( .B1(n12438), .B2(n8689), .C1(n12432), .C2(n8690), .A(n2378), .ZN(n2377) );
  OAI22_X1 U3420 ( .A1(n7846), .A2(n12426), .B1(n7847), .B2(n12420), .ZN(n2378) );
  AOI221_X1 U3421 ( .B1(n12438), .B2(n8691), .C1(n12432), .C2(n8692), .A(n2359), .ZN(n2358) );
  OAI22_X1 U3422 ( .A1(n7829), .A2(n12426), .B1(n7830), .B2(n12420), .ZN(n2359) );
  AOI221_X1 U3423 ( .B1(n12438), .B2(n8693), .C1(n12432), .C2(n8694), .A(n2340), .ZN(n2339) );
  OAI22_X1 U3424 ( .A1(n7812), .A2(n12426), .B1(n7813), .B2(n12420), .ZN(n2340) );
  AOI221_X1 U3425 ( .B1(n12438), .B2(n8695), .C1(n12432), .C2(n8696), .A(n2321), .ZN(n2320) );
  OAI22_X1 U3426 ( .A1(n7795), .A2(n12426), .B1(n7796), .B2(n12420), .ZN(n2321) );
  AOI221_X1 U3427 ( .B1(n12438), .B2(n4656), .C1(n12432), .C2(n4657), .A(n2302), .ZN(n2301) );
  OAI22_X1 U3428 ( .A1(n7778), .A2(n12426), .B1(n7779), .B2(n12420), .ZN(n2302) );
  AOI221_X1 U3429 ( .B1(n12439), .B2(n4658), .C1(n12433), .C2(n4659), .A(n2283), .ZN(n2282) );
  OAI22_X1 U3430 ( .A1(n7761), .A2(n12427), .B1(n7762), .B2(n12421), .ZN(n2283) );
  AOI221_X1 U3431 ( .B1(n12439), .B2(n4660), .C1(n12433), .C2(n4661), .A(n2264), .ZN(n2263) );
  OAI22_X1 U3432 ( .A1(n7744), .A2(n12427), .B1(n7745), .B2(n12421), .ZN(n2264) );
  AOI221_X1 U3433 ( .B1(n12439), .B2(n4662), .C1(n12433), .C2(n4663), .A(n2245), .ZN(n2244) );
  OAI22_X1 U3434 ( .A1(n7642), .A2(n12427), .B1(n7643), .B2(n12421), .ZN(n2245) );
  AOI221_X1 U3435 ( .B1(n12439), .B2(n4664), .C1(n12433), .C2(n4665), .A(n2226), .ZN(n2225) );
  OAI22_X1 U3436 ( .A1(n7625), .A2(n12427), .B1(n7626), .B2(n12421), .ZN(n2226) );
  AOI221_X1 U3437 ( .B1(n12439), .B2(n4666), .C1(n12433), .C2(n4667), .A(n2207), .ZN(n2206) );
  OAI22_X1 U3438 ( .A1(n7521), .A2(n12427), .B1(n7522), .B2(n12421), .ZN(n2207) );
  AOI221_X1 U3439 ( .B1(n12439), .B2(n4668), .C1(n12433), .C2(n4669), .A(n2188), .ZN(n2187) );
  OAI22_X1 U3440 ( .A1(n7504), .A2(n12427), .B1(n7505), .B2(n12421), .ZN(n2188) );
  AOI221_X1 U3441 ( .B1(n12439), .B2(n4670), .C1(n12433), .C2(n4671), .A(n2169), .ZN(n2168) );
  OAI22_X1 U3442 ( .A1(n7402), .A2(n12427), .B1(n7403), .B2(n12421), .ZN(n2169) );
  AOI221_X1 U3443 ( .B1(n12439), .B2(n4672), .C1(n12433), .C2(n4673), .A(n2150), .ZN(n2149) );
  OAI22_X1 U3444 ( .A1(n7385), .A2(n12427), .B1(n7386), .B2(n12421), .ZN(n2150) );
  AOI221_X1 U3445 ( .B1(n12439), .B2(n4674), .C1(n12433), .C2(n4675), .A(n2131), .ZN(n2130) );
  OAI22_X1 U3446 ( .A1(n7368), .A2(n12427), .B1(n7369), .B2(n12421), .ZN(n2131) );
  AOI221_X1 U3447 ( .B1(n12439), .B2(n4676), .C1(n12433), .C2(n4677), .A(n2112), .ZN(n2111) );
  OAI22_X1 U3448 ( .A1(n7269), .A2(n12427), .B1(n7270), .B2(n12421), .ZN(n2112) );
  AOI221_X1 U3449 ( .B1(n12439), .B2(n4678), .C1(n12433), .C2(n4679), .A(n2093), .ZN(n2092) );
  OAI22_X1 U3450 ( .A1(n7252), .A2(n12427), .B1(n7253), .B2(n12421), .ZN(n2093) );
  AOI221_X1 U3451 ( .B1(n12439), .B2(n4682), .C1(n12433), .C2(n4683), .A(n2074), .ZN(n2073) );
  OAI22_X1 U3452 ( .A1(n7235), .A2(n12427), .B1(n7236), .B2(n12421), .ZN(n2074) );
  AOI221_X1 U3453 ( .B1(n12440), .B2(n4472), .C1(n12434), .C2(n4473), .A(n2055), .ZN(n2054) );
  OAI22_X1 U3454 ( .A1(n7138), .A2(n12428), .B1(n7139), .B2(n12422), .ZN(n2055) );
  AOI221_X1 U3455 ( .B1(n12536), .B2(n9952), .C1(n12530), .C2(n9888), .A(n2047), .ZN(n2046) );
  OAI22_X1 U3456 ( .A1(n14435), .A2(n12524), .B1(n14412), .B2(n12518), .ZN(
        n2047) );
  AOI221_X1 U3457 ( .B1(n12440), .B2(n4474), .C1(n12434), .C2(n4475), .A(n2036), .ZN(n2035) );
  OAI22_X1 U3458 ( .A1(n7121), .A2(n12428), .B1(n7122), .B2(n12422), .ZN(n2036) );
  AOI221_X1 U3459 ( .B1(n12536), .B2(n9951), .C1(n12530), .C2(n9887), .A(n2028), .ZN(n2027) );
  OAI22_X1 U3460 ( .A1(n14434), .A2(n12524), .B1(n14411), .B2(n12518), .ZN(
        n2028) );
  AOI221_X1 U3461 ( .B1(n12440), .B2(n4476), .C1(n12434), .C2(n4477), .A(n2017), .ZN(n2016) );
  OAI22_X1 U3462 ( .A1(n4860), .A2(n12428), .B1(n4861), .B2(n12422), .ZN(n2017) );
  AOI221_X1 U3463 ( .B1(n12536), .B2(n9950), .C1(n12530), .C2(n9886), .A(n2009), .ZN(n2008) );
  OAI22_X1 U3464 ( .A1(n14433), .A2(n12524), .B1(n14410), .B2(n12518), .ZN(
        n2009) );
  AOI221_X1 U3465 ( .B1(n12440), .B2(n4478), .C1(n12434), .C2(n4479), .A(n1984), .ZN(n1981) );
  OAI22_X1 U3466 ( .A1(n4843), .A2(n12428), .B1(n4844), .B2(n12422), .ZN(n1984) );
  AOI221_X1 U3467 ( .B1(n12536), .B2(n9949), .C1(n12530), .C2(n9885), .A(n1960), .ZN(n1957) );
  OAI22_X1 U3468 ( .A1(n13392), .A2(n12524), .B1(n14409), .B2(n12518), .ZN(
        n1960) );
  AOI221_X1 U3469 ( .B1(n12411), .B2(n4480), .C1(n12405), .C2(n4481), .A(n3206), .ZN(n3201) );
  OAI22_X1 U3470 ( .A1(n8579), .A2(n12399), .B1(n8580), .B2(n12393), .ZN(n3206) );
  AOI221_X1 U3471 ( .B1(n12411), .B2(n4648), .C1(n12405), .C2(n4649), .A(n3177), .ZN(n3174) );
  OAI22_X1 U3472 ( .A1(n8562), .A2(n12399), .B1(n8563), .B2(n12393), .ZN(n3177) );
  AOI221_X1 U3473 ( .B1(n12411), .B2(n4482), .C1(n12405), .C2(n4483), .A(n3158), .ZN(n3155) );
  OAI22_X1 U3474 ( .A1(n8545), .A2(n12399), .B1(n8546), .B2(n12393), .ZN(n3158) );
  AOI221_X1 U3475 ( .B1(n12411), .B2(n4484), .C1(n12405), .C2(n4485), .A(n3139), .ZN(n3136) );
  OAI22_X1 U3476 ( .A1(n8528), .A2(n12399), .B1(n8529), .B2(n12393), .ZN(n3139) );
  AOI221_X1 U3477 ( .B1(n12411), .B2(n7080), .C1(n12405), .C2(n7081), .A(n3120), .ZN(n3117) );
  OAI22_X1 U3478 ( .A1(n8511), .A2(n12399), .B1(n8512), .B2(n12393), .ZN(n3120) );
  AOI221_X1 U3479 ( .B1(n12411), .B2(n8605), .C1(n12405), .C2(n8606), .A(n3101), .ZN(n3098) );
  OAI22_X1 U3480 ( .A1(n8494), .A2(n12399), .B1(n8495), .B2(n12393), .ZN(n3101) );
  AOI221_X1 U3481 ( .B1(n12411), .B2(n8613), .C1(n12405), .C2(n8614), .A(n3082), .ZN(n3079) );
  OAI22_X1 U3482 ( .A1(n8477), .A2(n12399), .B1(n8478), .B2(n12393), .ZN(n3082) );
  AOI221_X1 U3483 ( .B1(n12411), .B2(n7084), .C1(n12405), .C2(n7085), .A(n3063), .ZN(n3060) );
  OAI22_X1 U3484 ( .A1(n8460), .A2(n12399), .B1(n8461), .B2(n12393), .ZN(n3063) );
  AOI221_X1 U3485 ( .B1(n12411), .B2(n7088), .C1(n12405), .C2(n7089), .A(n3044), .ZN(n3041) );
  OAI22_X1 U3486 ( .A1(n8443), .A2(n12399), .B1(n8444), .B2(n12393), .ZN(n3044) );
  AOI221_X1 U3487 ( .B1(n12411), .B2(n7092), .C1(n12405), .C2(n7093), .A(n3025), .ZN(n3022) );
  OAI22_X1 U3488 ( .A1(n8426), .A2(n12399), .B1(n8427), .B2(n12393), .ZN(n3025) );
  AOI221_X1 U3489 ( .B1(n12411), .B2(n7096), .C1(n12405), .C2(n7097), .A(n3006), .ZN(n3003) );
  OAI22_X1 U3490 ( .A1(n8409), .A2(n12399), .B1(n8410), .B2(n12393), .ZN(n3006) );
  AOI221_X1 U3491 ( .B1(n12411), .B2(n7100), .C1(n12405), .C2(n7101), .A(n2987), .ZN(n2984) );
  OAI22_X1 U3492 ( .A1(n8392), .A2(n12399), .B1(n8393), .B2(n12393), .ZN(n2987) );
  AOI221_X1 U3493 ( .B1(n12412), .B2(n7104), .C1(n12406), .C2(n7105), .A(n2968), .ZN(n2965) );
  OAI22_X1 U3494 ( .A1(n8375), .A2(n12400), .B1(n8376), .B2(n12394), .ZN(n2968) );
  AOI221_X1 U3495 ( .B1(n12412), .B2(n7130), .C1(n12406), .C2(n7131), .A(n2949), .ZN(n2946) );
  OAI22_X1 U3496 ( .A1(n8358), .A2(n12400), .B1(n8359), .B2(n12394), .ZN(n2949) );
  AOI221_X1 U3497 ( .B1(n12412), .B2(n7154), .C1(n12406), .C2(n7155), .A(n2930), .ZN(n2927) );
  OAI22_X1 U3498 ( .A1(n8341), .A2(n12400), .B1(n8342), .B2(n12394), .ZN(n2930) );
  AOI221_X1 U3499 ( .B1(n12412), .B2(n7158), .C1(n12406), .C2(n7159), .A(n2911), .ZN(n2908) );
  OAI22_X1 U3500 ( .A1(n8324), .A2(n12400), .B1(n8325), .B2(n12394), .ZN(n2911) );
  AOI221_X1 U3501 ( .B1(n12412), .B2(n7162), .C1(n12406), .C2(n7163), .A(n2892), .ZN(n2889) );
  OAI22_X1 U3502 ( .A1(n8307), .A2(n12400), .B1(n8308), .B2(n12394), .ZN(n2892) );
  AOI221_X1 U3503 ( .B1(n12412), .B2(n7166), .C1(n12406), .C2(n7167), .A(n2873), .ZN(n2870) );
  OAI22_X1 U3504 ( .A1(n8290), .A2(n12400), .B1(n8291), .B2(n12394), .ZN(n2873) );
  AOI221_X1 U3505 ( .B1(n12412), .B2(n7170), .C1(n12406), .C2(n7171), .A(n2854), .ZN(n2851) );
  OAI22_X1 U3506 ( .A1(n8273), .A2(n12400), .B1(n8274), .B2(n12394), .ZN(n2854) );
  AOI221_X1 U3507 ( .B1(n12412), .B2(n7174), .C1(n12406), .C2(n7175), .A(n2835), .ZN(n2832) );
  OAI22_X1 U3508 ( .A1(n8256), .A2(n12400), .B1(n8257), .B2(n12394), .ZN(n2835) );
  AOI221_X1 U3509 ( .B1(n12412), .B2(n7178), .C1(n12406), .C2(n7179), .A(n2816), .ZN(n2813) );
  OAI22_X1 U3510 ( .A1(n8239), .A2(n12400), .B1(n8240), .B2(n12394), .ZN(n2816) );
  AOI221_X1 U3511 ( .B1(n12412), .B2(n7182), .C1(n12406), .C2(n7183), .A(n2797), .ZN(n2794) );
  OAI22_X1 U3512 ( .A1(n8222), .A2(n12400), .B1(n8223), .B2(n12394), .ZN(n2797) );
  AOI221_X1 U3513 ( .B1(n12412), .B2(n7186), .C1(n12406), .C2(n7187), .A(n2778), .ZN(n2775) );
  OAI22_X1 U3514 ( .A1(n8205), .A2(n12400), .B1(n8206), .B2(n12394), .ZN(n2778) );
  AOI221_X1 U3515 ( .B1(n12412), .B2(n7190), .C1(n12406), .C2(n7191), .A(n2759), .ZN(n2756) );
  OAI22_X1 U3516 ( .A1(n8188), .A2(n12400), .B1(n8189), .B2(n12394), .ZN(n2759) );
  AOI221_X1 U3517 ( .B1(n12413), .B2(n7194), .C1(n12407), .C2(n7195), .A(n2740), .ZN(n2737) );
  OAI22_X1 U3518 ( .A1(n8171), .A2(n12401), .B1(n8172), .B2(n12395), .ZN(n2740) );
  AOI221_X1 U3519 ( .B1(n12413), .B2(n7198), .C1(n12407), .C2(n7199), .A(n2721), .ZN(n2718) );
  OAI22_X1 U3520 ( .A1(n8154), .A2(n12401), .B1(n8155), .B2(n12395), .ZN(n2721) );
  AOI221_X1 U3521 ( .B1(n12413), .B2(n7202), .C1(n12407), .C2(n8708), .A(n2702), .ZN(n2699) );
  OAI22_X1 U3522 ( .A1(n8137), .A2(n12401), .B1(n8138), .B2(n12395), .ZN(n2702) );
  AOI221_X1 U3523 ( .B1(n12413), .B2(n7205), .C1(n12407), .C2(n8707), .A(n2683), .ZN(n2680) );
  OAI22_X1 U3524 ( .A1(n8120), .A2(n12401), .B1(n8121), .B2(n12395), .ZN(n2683) );
  AOI221_X1 U3525 ( .B1(n12413), .B2(n7208), .C1(n12407), .C2(n8706), .A(n2664), .ZN(n2661) );
  OAI22_X1 U3526 ( .A1(n8103), .A2(n12401), .B1(n8104), .B2(n12395), .ZN(n2664) );
  AOI221_X1 U3527 ( .B1(n12413), .B2(n7211), .C1(n12407), .C2(n8705), .A(n2645), .ZN(n2642) );
  OAI22_X1 U3528 ( .A1(n8086), .A2(n12401), .B1(n8087), .B2(n12395), .ZN(n2645) );
  AOI221_X1 U3529 ( .B1(n12413), .B2(n7214), .C1(n12407), .C2(n8704), .A(n2626), .ZN(n2623) );
  OAI22_X1 U3530 ( .A1(n8069), .A2(n12401), .B1(n8070), .B2(n12395), .ZN(n2626) );
  AOI221_X1 U3531 ( .B1(n12413), .B2(n7217), .C1(n12407), .C2(n8703), .A(n2607), .ZN(n2604) );
  OAI22_X1 U3532 ( .A1(n8052), .A2(n12401), .B1(n8053), .B2(n12395), .ZN(n2607) );
  AOI221_X1 U3533 ( .B1(n12413), .B2(n7220), .C1(n12407), .C2(n8702), .A(n2588), .ZN(n2585) );
  OAI22_X1 U3534 ( .A1(n8035), .A2(n12401), .B1(n8036), .B2(n12395), .ZN(n2588) );
  AOI221_X1 U3535 ( .B1(n12413), .B2(n7223), .C1(n12407), .C2(n8701), .A(n2569), .ZN(n2566) );
  OAI22_X1 U3536 ( .A1(n8018), .A2(n12401), .B1(n8019), .B2(n12395), .ZN(n2569) );
  AOI221_X1 U3537 ( .B1(n12413), .B2(n7226), .C1(n12407), .C2(n8700), .A(n2550), .ZN(n2547) );
  OAI22_X1 U3538 ( .A1(n8001), .A2(n12401), .B1(n8002), .B2(n12395), .ZN(n2550) );
  AOI221_X1 U3539 ( .B1(n12413), .B2(n7229), .C1(n12407), .C2(n8699), .A(n2531), .ZN(n2528) );
  OAI22_X1 U3540 ( .A1(n7984), .A2(n12401), .B1(n7985), .B2(n12395), .ZN(n2531) );
  AOI221_X1 U3541 ( .B1(n12414), .B2(n7232), .C1(n12408), .C2(n8698), .A(n2512), .ZN(n2509) );
  OAI22_X1 U3542 ( .A1(n7967), .A2(n12402), .B1(n7968), .B2(n12396), .ZN(n2512) );
  AOI221_X1 U3543 ( .B1(n12414), .B2(n7245), .C1(n12408), .C2(n8697), .A(n2493), .ZN(n2490) );
  OAI22_X1 U3544 ( .A1(n7950), .A2(n12402), .B1(n7951), .B2(n12396), .ZN(n2493) );
  AOI221_X1 U3545 ( .B1(n12414), .B2(n7278), .C1(n12408), .C2(n7279), .A(n2474), .ZN(n2471) );
  OAI22_X1 U3546 ( .A1(n7933), .A2(n12402), .B1(n7934), .B2(n12396), .ZN(n2474) );
  AOI221_X1 U3547 ( .B1(n12414), .B2(n7282), .C1(n12408), .C2(n7283), .A(n2455), .ZN(n2452) );
  OAI22_X1 U3548 ( .A1(n7916), .A2(n12402), .B1(n7917), .B2(n12396), .ZN(n2455) );
  AOI221_X1 U3549 ( .B1(n12414), .B2(n7286), .C1(n12408), .C2(n7287), .A(n2436), .ZN(n2433) );
  OAI22_X1 U3550 ( .A1(n7899), .A2(n12402), .B1(n7900), .B2(n12396), .ZN(n2436) );
  AOI221_X1 U3551 ( .B1(n12414), .B2(n7290), .C1(n12408), .C2(n7291), .A(n2417), .ZN(n2414) );
  OAI22_X1 U3552 ( .A1(n7882), .A2(n12402), .B1(n7883), .B2(n12396), .ZN(n2417) );
  AOI221_X1 U3553 ( .B1(n12414), .B2(n7294), .C1(n12408), .C2(n7295), .A(n2398), .ZN(n2395) );
  OAI22_X1 U3554 ( .A1(n7865), .A2(n12402), .B1(n7866), .B2(n12396), .ZN(n2398) );
  AOI221_X1 U3555 ( .B1(n12414), .B2(n7298), .C1(n12408), .C2(n7299), .A(n2379), .ZN(n2376) );
  OAI22_X1 U3556 ( .A1(n7848), .A2(n12402), .B1(n7849), .B2(n12396), .ZN(n2379) );
  AOI221_X1 U3557 ( .B1(n12414), .B2(n7302), .C1(n12408), .C2(n7303), .A(n2360), .ZN(n2357) );
  OAI22_X1 U3558 ( .A1(n7831), .A2(n12402), .B1(n7832), .B2(n12396), .ZN(n2360) );
  AOI221_X1 U3559 ( .B1(n12414), .B2(n7306), .C1(n12408), .C2(n7307), .A(n2341), .ZN(n2338) );
  OAI22_X1 U3560 ( .A1(n7814), .A2(n12402), .B1(n7815), .B2(n12396), .ZN(n2341) );
  AOI221_X1 U3561 ( .B1(n12414), .B2(n7310), .C1(n12408), .C2(n7311), .A(n2322), .ZN(n2319) );
  OAI22_X1 U3562 ( .A1(n7797), .A2(n12402), .B1(n7798), .B2(n12396), .ZN(n2322) );
  AOI221_X1 U3563 ( .B1(n12414), .B2(n7314), .C1(n12408), .C2(n7315), .A(n2303), .ZN(n2300) );
  OAI22_X1 U3564 ( .A1(n7780), .A2(n12402), .B1(n7781), .B2(n12396), .ZN(n2303) );
  AOI221_X1 U3565 ( .B1(n12415), .B2(n7318), .C1(n12409), .C2(n7319), .A(n2284), .ZN(n2281) );
  OAI22_X1 U3566 ( .A1(n7763), .A2(n12403), .B1(n7764), .B2(n12397), .ZN(n2284) );
  AOI221_X1 U3567 ( .B1(n12415), .B2(n7322), .C1(n12409), .C2(n7323), .A(n2265), .ZN(n2262) );
  OAI22_X1 U3568 ( .A1(n7746), .A2(n12403), .B1(n7747), .B2(n12397), .ZN(n2265) );
  AOI221_X1 U3569 ( .B1(n12415), .B2(n4486), .C1(n12409), .C2(n4487), .A(n2246), .ZN(n2243) );
  OAI22_X1 U3570 ( .A1(n7644), .A2(n12403), .B1(n7645), .B2(n12397), .ZN(n2246) );
  AOI221_X1 U3571 ( .B1(n12415), .B2(n4488), .C1(n12409), .C2(n4489), .A(n2227), .ZN(n2224) );
  OAI22_X1 U3572 ( .A1(n7627), .A2(n12403), .B1(n7628), .B2(n12397), .ZN(n2227) );
  AOI221_X1 U3573 ( .B1(n12415), .B2(n4490), .C1(n12409), .C2(n4491), .A(n2208), .ZN(n2205) );
  OAI22_X1 U3574 ( .A1(n7523), .A2(n12403), .B1(n7524), .B2(n12397), .ZN(n2208) );
  AOI221_X1 U3575 ( .B1(n12415), .B2(n4492), .C1(n12409), .C2(n4493), .A(n2189), .ZN(n2186) );
  OAI22_X1 U3576 ( .A1(n7506), .A2(n12403), .B1(n7507), .B2(n12397), .ZN(n2189) );
  AOI221_X1 U3577 ( .B1(n12415), .B2(n4494), .C1(n12409), .C2(n4495), .A(n2170), .ZN(n2167) );
  OAI22_X1 U3578 ( .A1(n7404), .A2(n12403), .B1(n7490), .B2(n12397), .ZN(n2170) );
  AOI221_X1 U3579 ( .B1(n12415), .B2(n4496), .C1(n12409), .C2(n4497), .A(n2151), .ZN(n2148) );
  OAI22_X1 U3580 ( .A1(n7387), .A2(n12403), .B1(n7388), .B2(n12397), .ZN(n2151) );
  AOI221_X1 U3581 ( .B1(n12415), .B2(n4498), .C1(n12409), .C2(n4499), .A(n2132), .ZN(n2129) );
  OAI22_X1 U3582 ( .A1(n7370), .A2(n12403), .B1(n7371), .B2(n12397), .ZN(n2132) );
  AOI221_X1 U3583 ( .B1(n12415), .B2(n4500), .C1(n12409), .C2(n4501), .A(n2113), .ZN(n2110) );
  OAI22_X1 U3584 ( .A1(n7271), .A2(n12403), .B1(n7272), .B2(n12397), .ZN(n2113) );
  AOI221_X1 U3585 ( .B1(n12415), .B2(n4502), .C1(n12409), .C2(n4503), .A(n2094), .ZN(n2091) );
  OAI22_X1 U3586 ( .A1(n7254), .A2(n12403), .B1(n7255), .B2(n12397), .ZN(n2094) );
  AOI221_X1 U3587 ( .B1(n12415), .B2(n4684), .C1(n12409), .C2(n4685), .A(n2075), .ZN(n2072) );
  OAI22_X1 U3588 ( .A1(n7237), .A2(n12403), .B1(n7238), .B2(n12397), .ZN(n2075) );
  AOI221_X1 U3589 ( .B1(n12416), .B2(n4504), .C1(n12410), .C2(n4505), .A(n2056), .ZN(n2053) );
  OAI22_X1 U3590 ( .A1(n7140), .A2(n12404), .B1(n7141), .B2(n12398), .ZN(n2056) );
  AOI221_X1 U3591 ( .B1(n12416), .B2(n4506), .C1(n12410), .C2(n4507), .A(n2037), .ZN(n2034) );
  OAI22_X1 U3592 ( .A1(n7123), .A2(n12404), .B1(n7124), .B2(n12398), .ZN(n2037) );
  AOI221_X1 U3593 ( .B1(n12416), .B2(n4508), .C1(n12410), .C2(n4509), .A(n2018), .ZN(n2015) );
  OAI22_X1 U3594 ( .A1(n7106), .A2(n12404), .B1(n7107), .B2(n12398), .ZN(n2018) );
  AOI221_X1 U3595 ( .B1(n12416), .B2(n4510), .C1(n12410), .C2(n4511), .A(n1989), .ZN(n1980) );
  OAI22_X1 U3596 ( .A1(n4845), .A2(n12404), .B1(n4846), .B2(n12398), .ZN(n1989) );
  AOI221_X1 U3597 ( .B1(n12531), .B2(n11766), .C1(n12525), .C2(n9948), .A(
        n3187), .ZN(n3186) );
  OAI22_X1 U3598 ( .A1(n14216), .A2(n12519), .B1(n13430), .B2(n12513), .ZN(
        n3187) );
  AOI221_X1 U3599 ( .B1(n12531), .B2(n11767), .C1(n12525), .C2(n9947), .A(
        n3168), .ZN(n3167) );
  OAI22_X1 U3600 ( .A1(n14328), .A2(n12519), .B1(n13429), .B2(n12513), .ZN(
        n3168) );
  AOI221_X1 U3601 ( .B1(n12531), .B2(n11768), .C1(n12525), .C2(n9946), .A(
        n3149), .ZN(n3148) );
  OAI22_X1 U3602 ( .A1(n14327), .A2(n12519), .B1(n13428), .B2(n12513), .ZN(
        n3149) );
  AOI221_X1 U3603 ( .B1(n12531), .B2(n11769), .C1(n12525), .C2(n9945), .A(
        n3130), .ZN(n3129) );
  OAI22_X1 U3604 ( .A1(n14326), .A2(n12519), .B1(n13427), .B2(n12513), .ZN(
        n3130) );
  AOI221_X1 U3605 ( .B1(n12531), .B2(n11770), .C1(n12525), .C2(n9944), .A(
        n3111), .ZN(n3110) );
  OAI22_X1 U3606 ( .A1(n14325), .A2(n12519), .B1(n13426), .B2(n12513), .ZN(
        n3111) );
  AOI221_X1 U3607 ( .B1(n12531), .B2(n11771), .C1(n12525), .C2(n9943), .A(
        n3092), .ZN(n3091) );
  OAI22_X1 U3608 ( .A1(n14324), .A2(n12519), .B1(n13425), .B2(n12513), .ZN(
        n3092) );
  AOI221_X1 U3609 ( .B1(n12531), .B2(n11772), .C1(n12525), .C2(n9942), .A(
        n3073), .ZN(n3072) );
  OAI22_X1 U3610 ( .A1(n14311), .A2(n12519), .B1(n13424), .B2(n12513), .ZN(
        n3073) );
  AOI221_X1 U3611 ( .B1(n12531), .B2(n11773), .C1(n12525), .C2(n9941), .A(
        n3054), .ZN(n3053) );
  OAI22_X1 U3612 ( .A1(n14310), .A2(n12519), .B1(n13423), .B2(n12513), .ZN(
        n3054) );
  AOI221_X1 U3613 ( .B1(n12531), .B2(n11774), .C1(n12525), .C2(n9940), .A(
        n3035), .ZN(n3034) );
  OAI22_X1 U3614 ( .A1(n14323), .A2(n12519), .B1(n13422), .B2(n12513), .ZN(
        n3035) );
  AOI221_X1 U3615 ( .B1(n12531), .B2(n11775), .C1(n12525), .C2(n9939), .A(
        n3016), .ZN(n3015) );
  OAI22_X1 U3616 ( .A1(n14309), .A2(n12519), .B1(n13421), .B2(n12513), .ZN(
        n3016) );
  AOI221_X1 U3617 ( .B1(n12531), .B2(n11776), .C1(n12525), .C2(n9938), .A(
        n2997), .ZN(n2996) );
  OAI22_X1 U3618 ( .A1(n14308), .A2(n12519), .B1(n13420), .B2(n12513), .ZN(
        n2997) );
  AOI221_X1 U3619 ( .B1(n12531), .B2(n11777), .C1(n12525), .C2(n9937), .A(
        n2978), .ZN(n2977) );
  OAI22_X1 U3620 ( .A1(n14307), .A2(n12519), .B1(n13419), .B2(n12513), .ZN(
        n2978) );
  AOI221_X1 U3621 ( .B1(n12532), .B2(n11778), .C1(n12526), .C2(n9936), .A(
        n2959), .ZN(n2958) );
  OAI22_X1 U3622 ( .A1(n14306), .A2(n12520), .B1(n13418), .B2(n12514), .ZN(
        n2959) );
  AOI221_X1 U3623 ( .B1(n12532), .B2(n9999), .C1(n12526), .C2(n9935), .A(n2940), .ZN(n2939) );
  OAI22_X1 U3624 ( .A1(n14305), .A2(n12520), .B1(n13417), .B2(n12514), .ZN(
        n2940) );
  AOI221_X1 U3625 ( .B1(n12532), .B2(n9998), .C1(n12526), .C2(n9934), .A(n2921), .ZN(n2920) );
  OAI22_X1 U3626 ( .A1(n14304), .A2(n12520), .B1(n13416), .B2(n12514), .ZN(
        n2921) );
  AOI221_X1 U3627 ( .B1(n12532), .B2(n9997), .C1(n12526), .C2(n9933), .A(n2902), .ZN(n2901) );
  OAI22_X1 U3628 ( .A1(n14303), .A2(n12520), .B1(n13415), .B2(n12514), .ZN(
        n2902) );
  AOI221_X1 U3629 ( .B1(n12532), .B2(n9996), .C1(n12526), .C2(n9932), .A(n2883), .ZN(n2882) );
  OAI22_X1 U3630 ( .A1(n14302), .A2(n12520), .B1(n13414), .B2(n12514), .ZN(
        n2883) );
  AOI221_X1 U3631 ( .B1(n12532), .B2(n9995), .C1(n12526), .C2(n9931), .A(n2864), .ZN(n2863) );
  OAI22_X1 U3632 ( .A1(n14301), .A2(n12520), .B1(n13413), .B2(n12514), .ZN(
        n2864) );
  AOI221_X1 U3633 ( .B1(n12532), .B2(n9994), .C1(n12526), .C2(n9930), .A(n2845), .ZN(n2844) );
  OAI22_X1 U3634 ( .A1(n14300), .A2(n12520), .B1(n13412), .B2(n12514), .ZN(
        n2845) );
  AOI221_X1 U3635 ( .B1(n12532), .B2(n9993), .C1(n12526), .C2(n9929), .A(n2826), .ZN(n2825) );
  OAI22_X1 U3636 ( .A1(n14299), .A2(n12520), .B1(n13411), .B2(n12514), .ZN(
        n2826) );
  AOI221_X1 U3637 ( .B1(n12532), .B2(n9992), .C1(n12526), .C2(n9928), .A(n2807), .ZN(n2806) );
  OAI22_X1 U3638 ( .A1(n14298), .A2(n12520), .B1(n13410), .B2(n12514), .ZN(
        n2807) );
  AOI221_X1 U3639 ( .B1(n12532), .B2(n9991), .C1(n12526), .C2(n9927), .A(n2788), .ZN(n2787) );
  OAI22_X1 U3640 ( .A1(n14297), .A2(n12520), .B1(n13409), .B2(n12514), .ZN(
        n2788) );
  AOI221_X1 U3641 ( .B1(n12532), .B2(n9990), .C1(n12526), .C2(n9926), .A(n2769), .ZN(n2768) );
  OAI22_X1 U3642 ( .A1(n14296), .A2(n12520), .B1(n13408), .B2(n12514), .ZN(
        n2769) );
  AOI221_X1 U3643 ( .B1(n12532), .B2(n9989), .C1(n12526), .C2(n9925), .A(n2750), .ZN(n2749) );
  OAI22_X1 U3644 ( .A1(n14295), .A2(n12520), .B1(n13407), .B2(n12514), .ZN(
        n2750) );
  AOI221_X1 U3645 ( .B1(n12533), .B2(n9988), .C1(n12527), .C2(n9924), .A(n2731), .ZN(n2730) );
  OAI22_X1 U3646 ( .A1(n14294), .A2(n12521), .B1(n13406), .B2(n12515), .ZN(
        n2731) );
  AOI221_X1 U3647 ( .B1(n12533), .B2(n9987), .C1(n12527), .C2(n9923), .A(n2712), .ZN(n2711) );
  OAI22_X1 U3648 ( .A1(n14293), .A2(n12521), .B1(n13405), .B2(n12515), .ZN(
        n2712) );
  AOI221_X1 U3649 ( .B1(n12533), .B2(n9986), .C1(n12527), .C2(n9922), .A(n2693), .ZN(n2692) );
  OAI22_X1 U3650 ( .A1(n14292), .A2(n12521), .B1(n13404), .B2(n12515), .ZN(
        n2693) );
  AOI221_X1 U3651 ( .B1(n12533), .B2(n9985), .C1(n12527), .C2(n9921), .A(n2674), .ZN(n2673) );
  OAI22_X1 U3652 ( .A1(n14291), .A2(n12521), .B1(n13403), .B2(n12515), .ZN(
        n2674) );
  AOI221_X1 U3653 ( .B1(n12533), .B2(n9984), .C1(n12527), .C2(n9920), .A(n2655), .ZN(n2654) );
  OAI22_X1 U3654 ( .A1(n14290), .A2(n12521), .B1(n13402), .B2(n12515), .ZN(
        n2655) );
  AOI221_X1 U3655 ( .B1(n12533), .B2(n9983), .C1(n12527), .C2(n9919), .A(n2636), .ZN(n2635) );
  OAI22_X1 U3656 ( .A1(n14289), .A2(n12521), .B1(n14322), .B2(n12515), .ZN(
        n2636) );
  AOI221_X1 U3657 ( .B1(n12533), .B2(n9982), .C1(n12527), .C2(n9918), .A(n2617), .ZN(n2616) );
  OAI22_X1 U3658 ( .A1(n14456), .A2(n12521), .B1(n14321), .B2(n12515), .ZN(
        n2617) );
  AOI221_X1 U3659 ( .B1(n12533), .B2(n9981), .C1(n12527), .C2(n9917), .A(n2598), .ZN(n2597) );
  OAI22_X1 U3660 ( .A1(n14455), .A2(n12521), .B1(n14320), .B2(n12515), .ZN(
        n2598) );
  AOI221_X1 U3661 ( .B1(n12533), .B2(n9980), .C1(n12527), .C2(n9916), .A(n2579), .ZN(n2578) );
  OAI22_X1 U3662 ( .A1(n14454), .A2(n12521), .B1(n14319), .B2(n12515), .ZN(
        n2579) );
  AOI221_X1 U3663 ( .B1(n12533), .B2(n9979), .C1(n12527), .C2(n9915), .A(n2560), .ZN(n2559) );
  OAI22_X1 U3664 ( .A1(n14453), .A2(n12521), .B1(n14318), .B2(n12515), .ZN(
        n2560) );
  AOI221_X1 U3665 ( .B1(n12533), .B2(n9978), .C1(n12527), .C2(n9914), .A(n2541), .ZN(n2540) );
  OAI22_X1 U3666 ( .A1(n14452), .A2(n12521), .B1(n14317), .B2(n12515), .ZN(
        n2541) );
  AOI221_X1 U3667 ( .B1(n12533), .B2(n9977), .C1(n12527), .C2(n9913), .A(n2522), .ZN(n2521) );
  OAI22_X1 U3668 ( .A1(n14451), .A2(n12521), .B1(n14316), .B2(n12515), .ZN(
        n2522) );
  AOI221_X1 U3669 ( .B1(n12534), .B2(n9976), .C1(n12528), .C2(n9912), .A(n2503), .ZN(n2502) );
  OAI22_X1 U3670 ( .A1(n14450), .A2(n12522), .B1(n14315), .B2(n12516), .ZN(
        n2503) );
  AOI221_X1 U3671 ( .B1(n12534), .B2(n9975), .C1(n12528), .C2(n9911), .A(n2484), .ZN(n2483) );
  OAI22_X1 U3672 ( .A1(n14449), .A2(n12522), .B1(n14314), .B2(n12516), .ZN(
        n2484) );
  AOI221_X1 U3673 ( .B1(n12534), .B2(n9974), .C1(n12528), .C2(n9910), .A(n2465), .ZN(n2464) );
  OAI22_X1 U3674 ( .A1(n14448), .A2(n12522), .B1(n14313), .B2(n12516), .ZN(
        n2465) );
  AOI221_X1 U3675 ( .B1(n12534), .B2(n9973), .C1(n12528), .C2(n9909), .A(n2446), .ZN(n2445) );
  OAI22_X1 U3676 ( .A1(n14447), .A2(n12522), .B1(n14312), .B2(n12516), .ZN(
        n2446) );
  AOI221_X1 U3677 ( .B1(n12534), .B2(n9972), .C1(n12528), .C2(n9908), .A(n2427), .ZN(n2426) );
  OAI22_X1 U3678 ( .A1(n14446), .A2(n12522), .B1(n14432), .B2(n12516), .ZN(
        n2427) );
  AOI221_X1 U3679 ( .B1(n12534), .B2(n9971), .C1(n12528), .C2(n9907), .A(n2408), .ZN(n2407) );
  OAI22_X1 U3680 ( .A1(n14445), .A2(n12522), .B1(n14431), .B2(n12516), .ZN(
        n2408) );
  AOI221_X1 U3681 ( .B1(n12534), .B2(n9970), .C1(n12528), .C2(n9906), .A(n2389), .ZN(n2388) );
  OAI22_X1 U3682 ( .A1(n14444), .A2(n12522), .B1(n14430), .B2(n12516), .ZN(
        n2389) );
  AOI221_X1 U3683 ( .B1(n12534), .B2(n9969), .C1(n12528), .C2(n9905), .A(n2370), .ZN(n2369) );
  OAI22_X1 U3684 ( .A1(n14443), .A2(n12522), .B1(n14429), .B2(n12516), .ZN(
        n2370) );
  AOI221_X1 U3685 ( .B1(n12534), .B2(n9968), .C1(n12528), .C2(n9904), .A(n2351), .ZN(n2350) );
  OAI22_X1 U3686 ( .A1(n14442), .A2(n12522), .B1(n14428), .B2(n12516), .ZN(
        n2351) );
  AOI221_X1 U3687 ( .B1(n12534), .B2(n9967), .C1(n12528), .C2(n9903), .A(n2332), .ZN(n2331) );
  OAI22_X1 U3688 ( .A1(n14441), .A2(n12522), .B1(n14427), .B2(n12516), .ZN(
        n2332) );
  AOI221_X1 U3689 ( .B1(n12534), .B2(n9966), .C1(n12528), .C2(n9902), .A(n2313), .ZN(n2312) );
  OAI22_X1 U3690 ( .A1(n13401), .A2(n12522), .B1(n14426), .B2(n12516), .ZN(
        n2313) );
  AOI221_X1 U3691 ( .B1(n12534), .B2(n9965), .C1(n12528), .C2(n9901), .A(n2294), .ZN(n2293) );
  OAI22_X1 U3692 ( .A1(n13400), .A2(n12522), .B1(n14425), .B2(n12516), .ZN(
        n2294) );
  AOI221_X1 U3693 ( .B1(n12535), .B2(n9964), .C1(n12529), .C2(n9900), .A(n2275), .ZN(n2274) );
  OAI22_X1 U3694 ( .A1(n13399), .A2(n12523), .B1(n14424), .B2(n12517), .ZN(
        n2275) );
  AOI221_X1 U3695 ( .B1(n12535), .B2(n9963), .C1(n12529), .C2(n9899), .A(n2256), .ZN(n2255) );
  OAI22_X1 U3696 ( .A1(n13398), .A2(n12523), .B1(n14423), .B2(n12517), .ZN(
        n2256) );
  AOI221_X1 U3697 ( .B1(n12535), .B2(n9962), .C1(n12529), .C2(n9898), .A(n2237), .ZN(n2236) );
  OAI22_X1 U3698 ( .A1(n13397), .A2(n12523), .B1(n14422), .B2(n12517), .ZN(
        n2237) );
  AOI221_X1 U3699 ( .B1(n12535), .B2(n9961), .C1(n12529), .C2(n9897), .A(n2218), .ZN(n2217) );
  OAI22_X1 U3700 ( .A1(n13396), .A2(n12523), .B1(n14421), .B2(n12517), .ZN(
        n2218) );
  AOI221_X1 U3701 ( .B1(n12535), .B2(n9960), .C1(n12529), .C2(n9896), .A(n2199), .ZN(n2198) );
  OAI22_X1 U3702 ( .A1(n13395), .A2(n12523), .B1(n14420), .B2(n12517), .ZN(
        n2199) );
  AOI221_X1 U3703 ( .B1(n12535), .B2(n9959), .C1(n12529), .C2(n9895), .A(n2180), .ZN(n2179) );
  OAI22_X1 U3704 ( .A1(n13394), .A2(n12523), .B1(n14419), .B2(n12517), .ZN(
        n2180) );
  AOI221_X1 U3705 ( .B1(n12535), .B2(n9958), .C1(n12529), .C2(n9894), .A(n2161), .ZN(n2160) );
  OAI22_X1 U3706 ( .A1(n13393), .A2(n12523), .B1(n14418), .B2(n12517), .ZN(
        n2161) );
  AOI221_X1 U3707 ( .B1(n12535), .B2(n9957), .C1(n12529), .C2(n9893), .A(n2142), .ZN(n2141) );
  OAI22_X1 U3708 ( .A1(n14440), .A2(n12523), .B1(n14417), .B2(n12517), .ZN(
        n2142) );
  AOI221_X1 U3709 ( .B1(n12535), .B2(n9956), .C1(n12529), .C2(n9892), .A(n2123), .ZN(n2122) );
  OAI22_X1 U3710 ( .A1(n14439), .A2(n12523), .B1(n14416), .B2(n12517), .ZN(
        n2123) );
  AOI221_X1 U3711 ( .B1(n12535), .B2(n9955), .C1(n12529), .C2(n9891), .A(n2104), .ZN(n2103) );
  OAI22_X1 U3712 ( .A1(n14438), .A2(n12523), .B1(n14415), .B2(n12517), .ZN(
        n2104) );
  AOI221_X1 U3713 ( .B1(n12535), .B2(n9954), .C1(n12529), .C2(n9890), .A(n2085), .ZN(n2084) );
  OAI22_X1 U3714 ( .A1(n14437), .A2(n12523), .B1(n14414), .B2(n12517), .ZN(
        n2085) );
  AOI221_X1 U3715 ( .B1(n12535), .B2(n9953), .C1(n12529), .C2(n9889), .A(n2066), .ZN(n2065) );
  OAI22_X1 U3716 ( .A1(n14436), .A2(n12523), .B1(n14413), .B2(n12517), .ZN(
        n2066) );
  OAI22_X1 U3717 ( .A1(n13122), .A2(n13242), .B1(n13112), .B2(n11959), .ZN(
        n6806) );
  OAI22_X1 U3718 ( .A1(n13122), .A2(n13245), .B1(n13112), .B2(n11960), .ZN(
        n6807) );
  OAI22_X1 U3719 ( .A1(n13122), .A2(n13248), .B1(n13112), .B2(n11961), .ZN(
        n6808) );
  OAI22_X1 U3720 ( .A1(n13122), .A2(n13251), .B1(n13112), .B2(n11962), .ZN(
        n6809) );
  OAI22_X1 U3721 ( .A1(n13122), .A2(n13254), .B1(n13112), .B2(n11963), .ZN(
        n6810) );
  OAI22_X1 U3722 ( .A1(n13121), .A2(n13257), .B1(n13112), .B2(n11964), .ZN(
        n6811) );
  OAI22_X1 U3723 ( .A1(n13121), .A2(n13260), .B1(n13112), .B2(n11965), .ZN(
        n6812) );
  OAI22_X1 U3724 ( .A1(n13121), .A2(n13263), .B1(n13112), .B2(n11966), .ZN(
        n6813) );
  OAI22_X1 U3725 ( .A1(n13121), .A2(n13266), .B1(n13112), .B2(n11967), .ZN(
        n6814) );
  OAI22_X1 U3726 ( .A1(n13121), .A2(n13269), .B1(n13112), .B2(n11968), .ZN(
        n6815) );
  OAI22_X1 U3727 ( .A1(n13120), .A2(n13272), .B1(n13112), .B2(n11969), .ZN(
        n6816) );
  OAI22_X1 U3728 ( .A1(n13120), .A2(n13275), .B1(n13112), .B2(n11970), .ZN(
        n6817) );
  OAI22_X1 U3729 ( .A1(n13120), .A2(n13278), .B1(n13112), .B2(n11971), .ZN(
        n6818) );
  OAI22_X1 U3730 ( .A1(n13120), .A2(n13281), .B1(n13113), .B2(n11972), .ZN(
        n6819) );
  OAI22_X1 U3731 ( .A1(n13120), .A2(n13284), .B1(n13113), .B2(n11973), .ZN(
        n6820) );
  OAI22_X1 U3732 ( .A1(n13119), .A2(n13287), .B1(n13113), .B2(n11974), .ZN(
        n6821) );
  OAI22_X1 U3733 ( .A1(n13119), .A2(n13290), .B1(n13113), .B2(n11975), .ZN(
        n6822) );
  OAI22_X1 U3734 ( .A1(n13119), .A2(n13293), .B1(n13113), .B2(n11976), .ZN(
        n6823) );
  OAI22_X1 U3735 ( .A1(n13119), .A2(n13296), .B1(n13113), .B2(n11977), .ZN(
        n6824) );
  OAI22_X1 U3736 ( .A1(n13119), .A2(n13299), .B1(n13113), .B2(n11978), .ZN(
        n6825) );
  OAI22_X1 U3737 ( .A1(n13118), .A2(n13302), .B1(n13113), .B2(n11979), .ZN(
        n6826) );
  OAI22_X1 U3738 ( .A1(n13118), .A2(n13305), .B1(n13113), .B2(n11980), .ZN(
        n6827) );
  OAI22_X1 U3739 ( .A1(n13118), .A2(n13308), .B1(n13113), .B2(n11981), .ZN(
        n6828) );
  OAI22_X1 U3740 ( .A1(n13118), .A2(n13311), .B1(n13113), .B2(n11982), .ZN(
        n6829) );
  OAI22_X1 U3741 ( .A1(n13118), .A2(n13314), .B1(n13113), .B2(n11983), .ZN(
        n6830) );
  OAI22_X1 U3742 ( .A1(n13117), .A2(n13317), .B1(n13113), .B2(n11984), .ZN(
        n6831) );
  OAI22_X1 U3743 ( .A1(n13117), .A2(n13320), .B1(n13114), .B2(n11985), .ZN(
        n6832) );
  OAI22_X1 U3744 ( .A1(n13117), .A2(n13323), .B1(n13114), .B2(n11986), .ZN(
        n6833) );
  OAI22_X1 U3745 ( .A1(n13117), .A2(n13326), .B1(n13114), .B2(n11987), .ZN(
        n6834) );
  OAI22_X1 U3746 ( .A1(n13117), .A2(n13329), .B1(n13114), .B2(n11988), .ZN(
        n6835) );
  OAI22_X1 U3747 ( .A1(n13116), .A2(n13332), .B1(n13114), .B2(n11989), .ZN(
        n6836) );
  OAI22_X1 U3748 ( .A1(n13116), .A2(n13335), .B1(n13114), .B2(n11990), .ZN(
        n6837) );
  OAI22_X1 U3749 ( .A1(n13116), .A2(n13338), .B1(n13114), .B2(n11991), .ZN(
        n6838) );
  OAI22_X1 U3750 ( .A1(n13116), .A2(n13341), .B1(n13114), .B2(n11992), .ZN(
        n6839) );
  OAI22_X1 U3751 ( .A1(n13116), .A2(n13344), .B1(n13114), .B2(n11993), .ZN(
        n6840) );
  OAI22_X1 U3752 ( .A1(n13115), .A2(n13347), .B1(n13114), .B2(n11994), .ZN(
        n6841) );
  OAI22_X1 U3753 ( .A1(n13115), .A2(n13350), .B1(n13114), .B2(n11995), .ZN(
        n6842) );
  OAI22_X1 U3754 ( .A1(n13115), .A2(n13353), .B1(n13114), .B2(n11996), .ZN(
        n6843) );
  OAI22_X1 U3755 ( .A1(n13115), .A2(n13356), .B1(n13114), .B2(n11997), .ZN(
        n6844) );
  OAI22_X1 U3756 ( .A1(n13147), .A2(n13173), .B1(n13133), .B2(n11779), .ZN(
        n6847) );
  OAI22_X1 U3757 ( .A1(n13147), .A2(n13176), .B1(n13134), .B2(n11780), .ZN(
        n6848) );
  OAI22_X1 U3758 ( .A1(n13147), .A2(n13179), .B1(n13131), .B2(n11781), .ZN(
        n6849) );
  OAI22_X1 U3759 ( .A1(n13146), .A2(n13182), .B1(n13133), .B2(n11782), .ZN(
        n6850) );
  OAI22_X1 U3760 ( .A1(n13146), .A2(n13185), .B1(n13134), .B2(n11783), .ZN(
        n6851) );
  OAI22_X1 U3761 ( .A1(n13146), .A2(n13188), .B1(n13130), .B2(n11784), .ZN(
        n6852) );
  OAI22_X1 U3762 ( .A1(n13146), .A2(n13191), .B1(n1910), .B2(n11785), .ZN(
        n6853) );
  OAI22_X1 U3763 ( .A1(n13146), .A2(n13194), .B1(n1910), .B2(n11786), .ZN(
        n6854) );
  OAI22_X1 U3764 ( .A1(n13145), .A2(n13197), .B1(n1910), .B2(n11787), .ZN(
        n6855) );
  OAI22_X1 U3765 ( .A1(n13145), .A2(n13200), .B1(n1910), .B2(n11788), .ZN(
        n6856) );
  OAI22_X1 U3766 ( .A1(n13145), .A2(n13203), .B1(n1910), .B2(n11789), .ZN(
        n6857) );
  OAI22_X1 U3767 ( .A1(n13145), .A2(n13206), .B1(n13131), .B2(n11790), .ZN(
        n6858) );
  OAI22_X1 U3768 ( .A1(n13145), .A2(n13209), .B1(n13131), .B2(n11791), .ZN(
        n6859) );
  OAI22_X1 U3769 ( .A1(n13144), .A2(n13212), .B1(n13131), .B2(n11792), .ZN(
        n6860) );
  OAI22_X1 U3770 ( .A1(n13144), .A2(n13215), .B1(n13131), .B2(n11793), .ZN(
        n6861) );
  OAI22_X1 U3771 ( .A1(n13144), .A2(n13218), .B1(n13131), .B2(n11794), .ZN(
        n6862) );
  OAI22_X1 U3772 ( .A1(n13144), .A2(n13221), .B1(n13131), .B2(n11795), .ZN(
        n6863) );
  OAI22_X1 U3773 ( .A1(n13144), .A2(n13224), .B1(n13131), .B2(n11796), .ZN(
        n6864) );
  OAI22_X1 U3774 ( .A1(n13143), .A2(n13227), .B1(n13131), .B2(n11797), .ZN(
        n6865) );
  OAI22_X1 U3775 ( .A1(n13143), .A2(n13230), .B1(n13131), .B2(n11798), .ZN(
        n6866) );
  OAI22_X1 U3776 ( .A1(n13143), .A2(n13233), .B1(n13131), .B2(n11799), .ZN(
        n6867) );
  OAI22_X1 U3777 ( .A1(n13143), .A2(n13236), .B1(n13131), .B2(n11800), .ZN(
        n6868) );
  OAI22_X1 U3778 ( .A1(n13143), .A2(n13239), .B1(n13131), .B2(n11801), .ZN(
        n6869) );
  OAI22_X1 U3779 ( .A1(n13147), .A2(n13170), .B1(n1910), .B2(n11802), .ZN(
        n6846) );
  OAI22_X1 U3780 ( .A1(n12804), .A2(n13219), .B1(n12791), .B2(n11803), .ZN(
        n5774) );
  OAI22_X1 U3781 ( .A1(n12806), .A2(n13183), .B1(n12793), .B2(n11804), .ZN(
        n5762) );
  OAI22_X1 U3782 ( .A1(n12806), .A2(n13186), .B1(n12794), .B2(n11805), .ZN(
        n5763) );
  OAI22_X1 U3783 ( .A1(n12806), .A2(n13189), .B1(n12791), .B2(n11806), .ZN(
        n5764) );
  OAI22_X1 U3784 ( .A1(n12806), .A2(n13192), .B1(n12793), .B2(n11807), .ZN(
        n5765) );
  OAI22_X1 U3785 ( .A1(n12805), .A2(n13198), .B1(n12794), .B2(n11808), .ZN(
        n5767) );
  OAI22_X1 U3786 ( .A1(n12805), .A2(n13201), .B1(n12790), .B2(n11809), .ZN(
        n5768) );
  OAI22_X1 U3787 ( .A1(n12805), .A2(n13204), .B1(n1936), .B2(n11810), .ZN(
        n5769) );
  OAI22_X1 U3788 ( .A1(n12726), .A2(n13183), .B1(n12712), .B2(n11811), .ZN(
        n5506) );
  OAI22_X1 U3789 ( .A1(n12726), .A2(n13186), .B1(n12714), .B2(n11812), .ZN(
        n5507) );
  OAI22_X1 U3790 ( .A1(n12726), .A2(n13189), .B1(n12711), .B2(n11813), .ZN(
        n5508) );
  OAI22_X1 U3791 ( .A1(n12726), .A2(n13192), .B1(n12712), .B2(n11814), .ZN(
        n5509) );
  OAI22_X1 U3792 ( .A1(n12726), .A2(n13195), .B1(n12714), .B2(n11815), .ZN(
        n5510) );
  OAI22_X1 U3793 ( .A1(n12725), .A2(n13198), .B1(n12710), .B2(n11816), .ZN(
        n5511) );
  OAI22_X1 U3794 ( .A1(n12725), .A2(n13201), .B1(n1940), .B2(n11817), .ZN(
        n5512) );
  OAI22_X1 U3795 ( .A1(n12725), .A2(n13204), .B1(n1940), .B2(n11818), .ZN(
        n5513) );
  OAI22_X1 U3796 ( .A1(n12725), .A2(n13207), .B1(n12711), .B2(n11819), .ZN(
        n5514) );
  OAI22_X1 U3797 ( .A1(n12725), .A2(n13210), .B1(n12711), .B2(n11820), .ZN(
        n5515) );
  OAI22_X1 U3798 ( .A1(n12806), .A2(n13195), .B1(n1936), .B2(n11821), .ZN(
        n5766) );
  OAI22_X1 U3799 ( .A1(n12805), .A2(n13207), .B1(n12791), .B2(n11822), .ZN(
        n5770) );
  OAI22_X1 U3800 ( .A1(n12805), .A2(n13210), .B1(n12791), .B2(n11823), .ZN(
        n5771) );
  OAI22_X1 U3801 ( .A1(n12804), .A2(n13213), .B1(n12791), .B2(n11824), .ZN(
        n5772) );
  OAI22_X1 U3802 ( .A1(n12804), .A2(n13216), .B1(n12791), .B2(n11825), .ZN(
        n5773) );
  OAI22_X1 U3803 ( .A1(n12804), .A2(n13222), .B1(n12791), .B2(n11826), .ZN(
        n5775) );
  OAI22_X1 U3804 ( .A1(n12804), .A2(n13225), .B1(n12791), .B2(n11827), .ZN(
        n5776) );
  OAI22_X1 U3805 ( .A1(n12803), .A2(n13228), .B1(n12791), .B2(n11828), .ZN(
        n5777) );
  OAI22_X1 U3806 ( .A1(n12803), .A2(n13231), .B1(n12791), .B2(n11829), .ZN(
        n5778) );
  OAI22_X1 U3807 ( .A1(n12803), .A2(n13234), .B1(n12791), .B2(n11830), .ZN(
        n5779) );
  OAI22_X1 U3808 ( .A1(n12803), .A2(n13237), .B1(n12791), .B2(n11831), .ZN(
        n5780) );
  OAI22_X1 U3809 ( .A1(n12803), .A2(n13240), .B1(n12791), .B2(n11832), .ZN(
        n5781) );
  OAI22_X1 U3810 ( .A1(n12724), .A2(n13213), .B1(n12711), .B2(n11833), .ZN(
        n5516) );
  OAI22_X1 U3811 ( .A1(n12724), .A2(n13216), .B1(n12711), .B2(n11834), .ZN(
        n5517) );
  OAI22_X1 U3812 ( .A1(n12724), .A2(n13219), .B1(n12711), .B2(n11835), .ZN(
        n5518) );
  OAI22_X1 U3813 ( .A1(n12724), .A2(n13222), .B1(n12711), .B2(n11836), .ZN(
        n5519) );
  OAI22_X1 U3814 ( .A1(n12724), .A2(n13225), .B1(n12711), .B2(n11837), .ZN(
        n5520) );
  OAI22_X1 U3815 ( .A1(n12723), .A2(n13228), .B1(n12711), .B2(n11838), .ZN(
        n5521) );
  OAI22_X1 U3816 ( .A1(n12723), .A2(n13231), .B1(n12711), .B2(n11839), .ZN(
        n5522) );
  OAI22_X1 U3817 ( .A1(n12723), .A2(n13234), .B1(n12711), .B2(n11840), .ZN(
        n5523) );
  OAI22_X1 U3818 ( .A1(n12723), .A2(n13237), .B1(n12711), .B2(n11841), .ZN(
        n5524) );
  OAI22_X1 U3819 ( .A1(n12723), .A2(n13240), .B1(n12711), .B2(n11842), .ZN(
        n5525) );
  OAI22_X1 U3820 ( .A1(n12727), .A2(n13171), .B1(n1940), .B2(n11843), .ZN(
        n5502) );
  OAI22_X1 U3821 ( .A1(n12727), .A2(n13174), .B1(n1940), .B2(n11844), .ZN(
        n5503) );
  OAI22_X1 U3822 ( .A1(n12727), .A2(n13177), .B1(n1940), .B2(n11845), .ZN(
        n5504) );
  OAI22_X1 U3823 ( .A1(n12727), .A2(n13180), .B1(n1940), .B2(n11846), .ZN(
        n5505) );
  OAI22_X1 U3824 ( .A1(n12747), .A2(n13171), .B1(n12731), .B2(n11998), .ZN(
        n5566) );
  OAI22_X1 U3825 ( .A1(n12747), .A2(n13174), .B1(n12731), .B2(n11999), .ZN(
        n5567) );
  OAI22_X1 U3826 ( .A1(n12747), .A2(n13177), .B1(n12731), .B2(n12000), .ZN(
        n5568) );
  OAI22_X1 U3827 ( .A1(n12747), .A2(n13180), .B1(n12731), .B2(n12001), .ZN(
        n5569) );
  OAI22_X1 U3828 ( .A1(n12746), .A2(n13183), .B1(n12731), .B2(n12002), .ZN(
        n5570) );
  OAI22_X1 U3829 ( .A1(n12746), .A2(n13186), .B1(n12731), .B2(n12003), .ZN(
        n5571) );
  OAI22_X1 U3830 ( .A1(n12746), .A2(n13189), .B1(n12731), .B2(n12004), .ZN(
        n5572) );
  OAI22_X1 U3831 ( .A1(n12746), .A2(n13192), .B1(n12731), .B2(n12005), .ZN(
        n5573) );
  OAI22_X1 U3832 ( .A1(n12746), .A2(n13195), .B1(n12731), .B2(n12006), .ZN(
        n5574) );
  OAI22_X1 U3833 ( .A1(n12745), .A2(n13198), .B1(n12731), .B2(n12007), .ZN(
        n5575) );
  OAI22_X1 U3834 ( .A1(n12745), .A2(n13201), .B1(n12731), .B2(n12008), .ZN(
        n5576) );
  OAI22_X1 U3835 ( .A1(n12745), .A2(n13204), .B1(n12731), .B2(n12009), .ZN(
        n5577) );
  OAI22_X1 U3836 ( .A1(n12745), .A2(n13207), .B1(n12733), .B2(n12010), .ZN(
        n5578) );
  OAI22_X1 U3837 ( .A1(n12745), .A2(n13210), .B1(n12734), .B2(n12011), .ZN(
        n5579) );
  OAI22_X1 U3838 ( .A1(n12744), .A2(n13213), .B1(n12731), .B2(n12012), .ZN(
        n5580) );
  OAI22_X1 U3839 ( .A1(n12744), .A2(n13216), .B1(n12733), .B2(n12013), .ZN(
        n5581) );
  OAI22_X1 U3840 ( .A1(n12744), .A2(n13219), .B1(n12734), .B2(n12014), .ZN(
        n5582) );
  OAI22_X1 U3841 ( .A1(n12744), .A2(n13222), .B1(n12730), .B2(n12015), .ZN(
        n5583) );
  OAI22_X1 U3842 ( .A1(n12744), .A2(n13225), .B1(n1939), .B2(n12016), .ZN(
        n5584) );
  OAI22_X1 U3843 ( .A1(n12743), .A2(n13228), .B1(n1939), .B2(n12017), .ZN(
        n5585) );
  OAI22_X1 U3844 ( .A1(n12743), .A2(n13231), .B1(n1939), .B2(n12018), .ZN(
        n5586) );
  OAI22_X1 U3845 ( .A1(n12743), .A2(n13234), .B1(n1939), .B2(n12019), .ZN(
        n5587) );
  OAI22_X1 U3846 ( .A1(n12743), .A2(n13237), .B1(n1939), .B2(n12020), .ZN(
        n5588) );
  OAI22_X1 U3847 ( .A1(n12743), .A2(n13240), .B1(n1939), .B2(n12021), .ZN(
        n5589) );
  OAI22_X1 U3848 ( .A1(n12807), .A2(n13171), .B1(n1936), .B2(n11847), .ZN(
        n5758) );
  OAI22_X1 U3849 ( .A1(n12807), .A2(n13174), .B1(n1936), .B2(n11848), .ZN(
        n5759) );
  OAI22_X1 U3850 ( .A1(n12807), .A2(n13177), .B1(n1936), .B2(n11849), .ZN(
        n5760) );
  OAI22_X1 U3851 ( .A1(n12807), .A2(n13180), .B1(n1936), .B2(n11850), .ZN(
        n5761) );
  OAI22_X1 U3852 ( .A1(n12827), .A2(n13171), .B1(n12811), .B2(n12022), .ZN(
        n5822) );
  OAI22_X1 U3853 ( .A1(n12827), .A2(n13174), .B1(n12811), .B2(n12023), .ZN(
        n5823) );
  OAI22_X1 U3854 ( .A1(n12827), .A2(n13177), .B1(n12811), .B2(n12024), .ZN(
        n5824) );
  OAI22_X1 U3855 ( .A1(n12827), .A2(n13180), .B1(n12811), .B2(n12025), .ZN(
        n5825) );
  OAI22_X1 U3856 ( .A1(n12826), .A2(n13183), .B1(n12811), .B2(n12026), .ZN(
        n5826) );
  OAI22_X1 U3857 ( .A1(n12826), .A2(n13186), .B1(n12811), .B2(n12027), .ZN(
        n5827) );
  OAI22_X1 U3858 ( .A1(n12826), .A2(n13189), .B1(n12811), .B2(n12028), .ZN(
        n5828) );
  OAI22_X1 U3859 ( .A1(n12826), .A2(n13192), .B1(n12811), .B2(n12029), .ZN(
        n5829) );
  OAI22_X1 U3860 ( .A1(n12826), .A2(n13195), .B1(n12811), .B2(n12030), .ZN(
        n5830) );
  OAI22_X1 U3861 ( .A1(n12825), .A2(n13198), .B1(n12811), .B2(n12031), .ZN(
        n5831) );
  OAI22_X1 U3862 ( .A1(n12825), .A2(n13201), .B1(n12811), .B2(n12032), .ZN(
        n5832) );
  OAI22_X1 U3863 ( .A1(n12825), .A2(n13204), .B1(n12811), .B2(n12033), .ZN(
        n5833) );
  OAI22_X1 U3864 ( .A1(n12825), .A2(n13207), .B1(n12813), .B2(n12034), .ZN(
        n5834) );
  OAI22_X1 U3865 ( .A1(n12825), .A2(n13210), .B1(n12814), .B2(n12035), .ZN(
        n5835) );
  OAI22_X1 U3866 ( .A1(n12824), .A2(n13213), .B1(n12811), .B2(n12036), .ZN(
        n5836) );
  OAI22_X1 U3867 ( .A1(n12824), .A2(n13216), .B1(n12813), .B2(n12037), .ZN(
        n5837) );
  OAI22_X1 U3868 ( .A1(n12824), .A2(n13219), .B1(n12814), .B2(n12038), .ZN(
        n5838) );
  OAI22_X1 U3869 ( .A1(n12824), .A2(n13222), .B1(n12810), .B2(n12039), .ZN(
        n5839) );
  OAI22_X1 U3870 ( .A1(n12824), .A2(n13225), .B1(n1935), .B2(n12040), .ZN(
        n5840) );
  OAI22_X1 U3871 ( .A1(n12823), .A2(n13228), .B1(n1935), .B2(n12041), .ZN(
        n5841) );
  OAI22_X1 U3872 ( .A1(n12823), .A2(n13231), .B1(n1935), .B2(n12042), .ZN(
        n5842) );
  OAI22_X1 U3873 ( .A1(n12823), .A2(n13234), .B1(n1935), .B2(n12043), .ZN(
        n5843) );
  OAI22_X1 U3874 ( .A1(n12823), .A2(n13237), .B1(n1935), .B2(n12044), .ZN(
        n5844) );
  OAI22_X1 U3875 ( .A1(n12823), .A2(n13240), .B1(n1935), .B2(n12045), .ZN(
        n5845) );
  OAI22_X1 U3876 ( .A1(n13125), .A2(n13209), .B1(n13111), .B2(n12046), .ZN(
        n6795) );
  OAI22_X1 U3877 ( .A1(n13124), .A2(n13212), .B1(n13111), .B2(n12047), .ZN(
        n6796) );
  OAI22_X1 U3878 ( .A1(n13124), .A2(n13215), .B1(n13111), .B2(n12048), .ZN(
        n6797) );
  OAI22_X1 U3879 ( .A1(n13124), .A2(n13218), .B1(n13111), .B2(n12049), .ZN(
        n6798) );
  OAI22_X1 U3880 ( .A1(n13124), .A2(n13221), .B1(n13111), .B2(n12050), .ZN(
        n6799) );
  OAI22_X1 U3881 ( .A1(n13124), .A2(n13224), .B1(n13111), .B2(n12051), .ZN(
        n6800) );
  OAI22_X1 U3882 ( .A1(n13123), .A2(n13227), .B1(n13111), .B2(n12052), .ZN(
        n6801) );
  OAI22_X1 U3883 ( .A1(n13123), .A2(n13230), .B1(n13111), .B2(n12053), .ZN(
        n6802) );
  OAI22_X1 U3884 ( .A1(n13123), .A2(n13233), .B1(n13111), .B2(n12054), .ZN(
        n6803) );
  OAI22_X1 U3885 ( .A1(n13123), .A2(n13236), .B1(n13111), .B2(n12055), .ZN(
        n6804) );
  OAI22_X1 U3886 ( .A1(n13123), .A2(n13239), .B1(n13111), .B2(n12056), .ZN(
        n6805) );
  OAI22_X1 U3887 ( .A1(n13142), .A2(n13242), .B1(n13132), .B2(n11851), .ZN(
        n6870) );
  OAI22_X1 U3888 ( .A1(n13142), .A2(n13245), .B1(n13132), .B2(n11852), .ZN(
        n6871) );
  OAI22_X1 U3889 ( .A1(n13142), .A2(n13248), .B1(n13132), .B2(n11853), .ZN(
        n6872) );
  OAI22_X1 U3890 ( .A1(n13142), .A2(n13251), .B1(n13132), .B2(n11854), .ZN(
        n6873) );
  OAI22_X1 U3891 ( .A1(n13142), .A2(n13254), .B1(n13132), .B2(n11855), .ZN(
        n6874) );
  OAI22_X1 U3892 ( .A1(n13141), .A2(n13257), .B1(n13132), .B2(n11856), .ZN(
        n6875) );
  OAI22_X1 U3893 ( .A1(n13141), .A2(n13260), .B1(n13132), .B2(n11857), .ZN(
        n6876) );
  OAI22_X1 U3894 ( .A1(n13141), .A2(n13263), .B1(n13132), .B2(n11858), .ZN(
        n6877) );
  OAI22_X1 U3895 ( .A1(n13141), .A2(n13266), .B1(n13132), .B2(n11859), .ZN(
        n6878) );
  OAI22_X1 U3896 ( .A1(n13141), .A2(n13269), .B1(n13132), .B2(n11860), .ZN(
        n6879) );
  OAI22_X1 U3897 ( .A1(n13140), .A2(n13272), .B1(n13132), .B2(n11861), .ZN(
        n6880) );
  OAI22_X1 U3898 ( .A1(n13140), .A2(n13275), .B1(n13132), .B2(n11862), .ZN(
        n6881) );
  OAI22_X1 U3899 ( .A1(n13140), .A2(n13278), .B1(n13133), .B2(n11863), .ZN(
        n6882) );
  OAI22_X1 U3900 ( .A1(n13140), .A2(n13281), .B1(n13133), .B2(n11864), .ZN(
        n6883) );
  OAI22_X1 U3901 ( .A1(n13140), .A2(n13284), .B1(n13133), .B2(n11865), .ZN(
        n6884) );
  OAI22_X1 U3902 ( .A1(n13139), .A2(n13287), .B1(n13133), .B2(n11866), .ZN(
        n6885) );
  OAI22_X1 U3903 ( .A1(n13139), .A2(n13290), .B1(n13133), .B2(n11867), .ZN(
        n6886) );
  OAI22_X1 U3904 ( .A1(n13139), .A2(n13293), .B1(n13133), .B2(n11868), .ZN(
        n6887) );
  OAI22_X1 U3905 ( .A1(n13139), .A2(n13296), .B1(n13133), .B2(n11869), .ZN(
        n6888) );
  OAI22_X1 U3906 ( .A1(n13139), .A2(n13299), .B1(n13133), .B2(n11870), .ZN(
        n6889) );
  OAI22_X1 U3907 ( .A1(n13138), .A2(n13302), .B1(n13133), .B2(n11871), .ZN(
        n6890) );
  OAI22_X1 U3908 ( .A1(n13138), .A2(n13305), .B1(n13133), .B2(n11872), .ZN(
        n6891) );
  OAI22_X1 U3909 ( .A1(n13138), .A2(n13308), .B1(n13133), .B2(n11873), .ZN(
        n6892) );
  OAI22_X1 U3910 ( .A1(n13138), .A2(n13311), .B1(n13133), .B2(n11874), .ZN(
        n6893) );
  OAI22_X1 U3911 ( .A1(n13138), .A2(n13314), .B1(n13134), .B2(n11875), .ZN(
        n6894) );
  OAI22_X1 U3912 ( .A1(n13137), .A2(n13317), .B1(n13134), .B2(n11876), .ZN(
        n6895) );
  OAI22_X1 U3913 ( .A1(n13137), .A2(n13320), .B1(n13134), .B2(n11877), .ZN(
        n6896) );
  OAI22_X1 U3914 ( .A1(n13137), .A2(n13323), .B1(n13134), .B2(n11878), .ZN(
        n6897) );
  OAI22_X1 U3915 ( .A1(n13137), .A2(n13326), .B1(n13134), .B2(n11879), .ZN(
        n6898) );
  OAI22_X1 U3916 ( .A1(n13137), .A2(n13329), .B1(n13134), .B2(n11880), .ZN(
        n6899) );
  OAI22_X1 U3917 ( .A1(n13136), .A2(n13332), .B1(n13134), .B2(n11881), .ZN(
        n6900) );
  OAI22_X1 U3918 ( .A1(n13136), .A2(n13335), .B1(n13134), .B2(n11882), .ZN(
        n6901) );
  OAI22_X1 U3919 ( .A1(n13136), .A2(n13338), .B1(n13134), .B2(n11883), .ZN(
        n6902) );
  OAI22_X1 U3920 ( .A1(n13136), .A2(n13341), .B1(n13134), .B2(n11884), .ZN(
        n6903) );
  OAI22_X1 U3921 ( .A1(n13136), .A2(n13344), .B1(n13134), .B2(n11885), .ZN(
        n6904) );
  OAI22_X1 U3922 ( .A1(n13135), .A2(n13347), .B1(n13134), .B2(n11886), .ZN(
        n6905) );
  OAI22_X1 U3923 ( .A1(n12802), .A2(n13243), .B1(n12792), .B2(n11887), .ZN(
        n5782) );
  OAI22_X1 U3924 ( .A1(n12802), .A2(n13246), .B1(n12792), .B2(n11888), .ZN(
        n5783) );
  OAI22_X1 U3925 ( .A1(n12802), .A2(n13249), .B1(n12792), .B2(n11889), .ZN(
        n5784) );
  OAI22_X1 U3926 ( .A1(n12802), .A2(n13252), .B1(n12792), .B2(n11890), .ZN(
        n5785) );
  OAI22_X1 U3927 ( .A1(n12802), .A2(n13255), .B1(n12792), .B2(n11891), .ZN(
        n5786) );
  OAI22_X1 U3928 ( .A1(n12801), .A2(n13258), .B1(n12792), .B2(n11892), .ZN(
        n5787) );
  OAI22_X1 U3929 ( .A1(n12801), .A2(n13261), .B1(n12792), .B2(n11893), .ZN(
        n5788) );
  OAI22_X1 U3930 ( .A1(n12801), .A2(n13264), .B1(n12792), .B2(n11894), .ZN(
        n5789) );
  OAI22_X1 U3931 ( .A1(n12801), .A2(n13267), .B1(n12792), .B2(n11895), .ZN(
        n5790) );
  OAI22_X1 U3932 ( .A1(n12801), .A2(n13270), .B1(n12792), .B2(n11896), .ZN(
        n5791) );
  OAI22_X1 U3933 ( .A1(n12800), .A2(n13273), .B1(n12792), .B2(n11897), .ZN(
        n5792) );
  OAI22_X1 U3934 ( .A1(n12800), .A2(n13276), .B1(n12792), .B2(n11898), .ZN(
        n5793) );
  OAI22_X1 U3935 ( .A1(n12800), .A2(n13279), .B1(n12793), .B2(n11899), .ZN(
        n5794) );
  OAI22_X1 U3936 ( .A1(n12800), .A2(n13282), .B1(n12793), .B2(n11900), .ZN(
        n5795) );
  OAI22_X1 U3937 ( .A1(n12800), .A2(n13285), .B1(n12793), .B2(n11901), .ZN(
        n5796) );
  OAI22_X1 U3938 ( .A1(n12799), .A2(n13288), .B1(n12793), .B2(n11902), .ZN(
        n5797) );
  OAI22_X1 U3939 ( .A1(n12799), .A2(n13291), .B1(n12793), .B2(n11903), .ZN(
        n5798) );
  OAI22_X1 U3940 ( .A1(n12799), .A2(n13294), .B1(n12793), .B2(n11904), .ZN(
        n5799) );
  OAI22_X1 U3941 ( .A1(n12799), .A2(n13297), .B1(n12793), .B2(n11905), .ZN(
        n5800) );
  OAI22_X1 U3942 ( .A1(n12799), .A2(n13300), .B1(n12793), .B2(n11906), .ZN(
        n5801) );
  OAI22_X1 U3943 ( .A1(n12798), .A2(n13303), .B1(n12793), .B2(n11907), .ZN(
        n5802) );
  OAI22_X1 U3944 ( .A1(n12798), .A2(n13306), .B1(n12793), .B2(n11908), .ZN(
        n5803) );
  OAI22_X1 U3945 ( .A1(n12798), .A2(n13309), .B1(n12793), .B2(n11909), .ZN(
        n5804) );
  OAI22_X1 U3946 ( .A1(n12722), .A2(n13249), .B1(n12712), .B2(n11910), .ZN(
        n5528) );
  OAI22_X1 U3947 ( .A1(n12722), .A2(n13252), .B1(n12712), .B2(n11911), .ZN(
        n5529) );
  OAI22_X1 U3948 ( .A1(n12722), .A2(n13255), .B1(n12712), .B2(n11912), .ZN(
        n5530) );
  OAI22_X1 U3949 ( .A1(n12721), .A2(n13258), .B1(n12712), .B2(n11913), .ZN(
        n5531) );
  OAI22_X1 U3950 ( .A1(n12721), .A2(n13261), .B1(n12712), .B2(n11914), .ZN(
        n5532) );
  OAI22_X1 U3951 ( .A1(n12721), .A2(n13264), .B1(n12712), .B2(n11915), .ZN(
        n5533) );
  OAI22_X1 U3952 ( .A1(n12721), .A2(n13267), .B1(n12712), .B2(n11916), .ZN(
        n5534) );
  OAI22_X1 U3953 ( .A1(n12721), .A2(n13270), .B1(n12712), .B2(n11917), .ZN(
        n5535) );
  OAI22_X1 U3954 ( .A1(n12720), .A2(n13273), .B1(n12712), .B2(n11918), .ZN(
        n5536) );
  OAI22_X1 U3955 ( .A1(n12720), .A2(n13276), .B1(n12712), .B2(n11919), .ZN(
        n5537) );
  OAI22_X1 U3956 ( .A1(n12720), .A2(n13279), .B1(n12713), .B2(n11920), .ZN(
        n5538) );
  OAI22_X1 U3957 ( .A1(n12720), .A2(n13282), .B1(n12713), .B2(n11921), .ZN(
        n5539) );
  OAI22_X1 U3958 ( .A1(n12720), .A2(n13285), .B1(n12713), .B2(n11922), .ZN(
        n5540) );
  OAI22_X1 U3959 ( .A1(n12719), .A2(n13288), .B1(n12713), .B2(n11923), .ZN(
        n5541) );
  OAI22_X1 U3960 ( .A1(n12719), .A2(n13291), .B1(n12713), .B2(n11924), .ZN(
        n5542) );
  OAI22_X1 U3961 ( .A1(n12719), .A2(n13294), .B1(n12713), .B2(n11925), .ZN(
        n5543) );
  OAI22_X1 U3962 ( .A1(n12719), .A2(n13297), .B1(n12713), .B2(n11926), .ZN(
        n5544) );
  OAI22_X1 U3963 ( .A1(n12719), .A2(n13300), .B1(n12713), .B2(n11927), .ZN(
        n5545) );
  OAI22_X1 U3964 ( .A1(n12718), .A2(n13303), .B1(n12713), .B2(n11928), .ZN(
        n5546) );
  OAI22_X1 U3965 ( .A1(n12718), .A2(n13306), .B1(n12713), .B2(n11929), .ZN(
        n5547) );
  OAI22_X1 U3966 ( .A1(n12718), .A2(n13309), .B1(n12713), .B2(n11930), .ZN(
        n5548) );
  OAI22_X1 U3967 ( .A1(n12718), .A2(n13312), .B1(n12713), .B2(n11931), .ZN(
        n5549) );
  OAI22_X1 U3968 ( .A1(n12718), .A2(n13315), .B1(n12714), .B2(n11932), .ZN(
        n5550) );
  OAI22_X1 U3969 ( .A1(n12717), .A2(n13318), .B1(n12714), .B2(n11933), .ZN(
        n5551) );
  OAI22_X1 U3970 ( .A1(n12722), .A2(n13243), .B1(n12712), .B2(n11934), .ZN(
        n5526) );
  OAI22_X1 U3971 ( .A1(n12722), .A2(n13246), .B1(n12712), .B2(n11935), .ZN(
        n5527) );
  OAI22_X1 U3972 ( .A1(n12717), .A2(n13321), .B1(n12714), .B2(n11936), .ZN(
        n5552) );
  OAI22_X1 U3973 ( .A1(n12717), .A2(n13324), .B1(n12714), .B2(n11937), .ZN(
        n5553) );
  OAI22_X1 U3974 ( .A1(n12717), .A2(n13327), .B1(n12714), .B2(n11938), .ZN(
        n5554) );
  OAI22_X1 U3975 ( .A1(n12717), .A2(n13330), .B1(n12714), .B2(n11939), .ZN(
        n5555) );
  OAI22_X1 U3976 ( .A1(n12716), .A2(n13333), .B1(n12714), .B2(n11940), .ZN(
        n5556) );
  OAI22_X1 U3977 ( .A1(n12716), .A2(n13336), .B1(n12714), .B2(n11941), .ZN(
        n5557) );
  OAI22_X1 U3978 ( .A1(n12716), .A2(n13339), .B1(n12714), .B2(n11942), .ZN(
        n5558) );
  OAI22_X1 U3979 ( .A1(n12716), .A2(n13342), .B1(n12714), .B2(n11943), .ZN(
        n5559) );
  OAI22_X1 U3980 ( .A1(n12716), .A2(n13345), .B1(n12714), .B2(n11944), .ZN(
        n5560) );
  OAI22_X1 U3981 ( .A1(n12715), .A2(n13348), .B1(n12714), .B2(n11945), .ZN(
        n5561) );
  OAI22_X1 U3982 ( .A1(n12742), .A2(n13243), .B1(n12732), .B2(n12057), .ZN(
        n5590) );
  OAI22_X1 U3983 ( .A1(n12742), .A2(n13246), .B1(n12732), .B2(n12058), .ZN(
        n5591) );
  OAI22_X1 U3984 ( .A1(n12742), .A2(n13249), .B1(n12732), .B2(n12059), .ZN(
        n5592) );
  OAI22_X1 U3985 ( .A1(n12742), .A2(n13252), .B1(n12732), .B2(n12060), .ZN(
        n5593) );
  OAI22_X1 U3986 ( .A1(n12742), .A2(n13255), .B1(n12732), .B2(n12061), .ZN(
        n5594) );
  OAI22_X1 U3987 ( .A1(n12741), .A2(n13258), .B1(n12732), .B2(n12062), .ZN(
        n5595) );
  OAI22_X1 U3988 ( .A1(n12741), .A2(n13261), .B1(n12732), .B2(n12063), .ZN(
        n5596) );
  OAI22_X1 U3989 ( .A1(n12741), .A2(n13264), .B1(n12732), .B2(n12064), .ZN(
        n5597) );
  OAI22_X1 U3990 ( .A1(n12741), .A2(n13267), .B1(n12732), .B2(n12065), .ZN(
        n5598) );
  OAI22_X1 U3991 ( .A1(n12741), .A2(n13270), .B1(n12732), .B2(n12066), .ZN(
        n5599) );
  OAI22_X1 U3992 ( .A1(n12740), .A2(n13273), .B1(n12732), .B2(n12067), .ZN(
        n5600) );
  OAI22_X1 U3993 ( .A1(n12740), .A2(n13276), .B1(n12732), .B2(n12068), .ZN(
        n5601) );
  OAI22_X1 U3994 ( .A1(n12740), .A2(n13279), .B1(n12733), .B2(n12069), .ZN(
        n5602) );
  OAI22_X1 U3995 ( .A1(n12740), .A2(n13282), .B1(n12733), .B2(n12070), .ZN(
        n5603) );
  OAI22_X1 U3996 ( .A1(n12740), .A2(n13285), .B1(n12733), .B2(n12071), .ZN(
        n5604) );
  OAI22_X1 U3997 ( .A1(n12739), .A2(n13288), .B1(n12733), .B2(n12072), .ZN(
        n5605) );
  OAI22_X1 U3998 ( .A1(n12739), .A2(n13291), .B1(n12733), .B2(n12073), .ZN(
        n5606) );
  OAI22_X1 U3999 ( .A1(n12739), .A2(n13294), .B1(n12733), .B2(n12074), .ZN(
        n5607) );
  OAI22_X1 U4000 ( .A1(n12739), .A2(n13297), .B1(n12733), .B2(n12075), .ZN(
        n5608) );
  OAI22_X1 U4001 ( .A1(n12739), .A2(n13300), .B1(n12733), .B2(n12076), .ZN(
        n5609) );
  OAI22_X1 U4002 ( .A1(n12738), .A2(n13303), .B1(n12733), .B2(n12077), .ZN(
        n5610) );
  OAI22_X1 U4003 ( .A1(n12738), .A2(n13306), .B1(n12733), .B2(n12078), .ZN(
        n5611) );
  OAI22_X1 U4004 ( .A1(n12738), .A2(n13309), .B1(n12733), .B2(n12079), .ZN(
        n5612) );
  OAI22_X1 U4005 ( .A1(n12738), .A2(n13312), .B1(n12733), .B2(n12080), .ZN(
        n5613) );
  OAI22_X1 U4006 ( .A1(n12738), .A2(n13315), .B1(n12734), .B2(n12081), .ZN(
        n5614) );
  OAI22_X1 U4007 ( .A1(n12737), .A2(n13318), .B1(n12734), .B2(n12082), .ZN(
        n5615) );
  OAI22_X1 U4008 ( .A1(n12737), .A2(n13321), .B1(n12734), .B2(n12083), .ZN(
        n5616) );
  OAI22_X1 U4009 ( .A1(n12737), .A2(n13324), .B1(n12734), .B2(n12084), .ZN(
        n5617) );
  OAI22_X1 U4010 ( .A1(n12737), .A2(n13327), .B1(n12734), .B2(n12085), .ZN(
        n5618) );
  OAI22_X1 U4011 ( .A1(n12737), .A2(n13330), .B1(n12734), .B2(n12086), .ZN(
        n5619) );
  OAI22_X1 U4012 ( .A1(n12736), .A2(n13333), .B1(n12734), .B2(n12087), .ZN(
        n5620) );
  OAI22_X1 U4013 ( .A1(n12736), .A2(n13336), .B1(n12734), .B2(n12088), .ZN(
        n5621) );
  OAI22_X1 U4014 ( .A1(n12736), .A2(n13339), .B1(n12734), .B2(n12089), .ZN(
        n5622) );
  OAI22_X1 U4015 ( .A1(n12736), .A2(n13342), .B1(n12734), .B2(n12090), .ZN(
        n5623) );
  OAI22_X1 U4016 ( .A1(n12736), .A2(n13345), .B1(n12734), .B2(n12091), .ZN(
        n5624) );
  OAI22_X1 U4017 ( .A1(n12735), .A2(n13348), .B1(n12734), .B2(n12092), .ZN(
        n5625) );
  OAI22_X1 U4018 ( .A1(n12798), .A2(n13312), .B1(n12793), .B2(n11946), .ZN(
        n5805) );
  OAI22_X1 U4019 ( .A1(n12798), .A2(n13315), .B1(n12794), .B2(n11947), .ZN(
        n5806) );
  OAI22_X1 U4020 ( .A1(n12797), .A2(n13318), .B1(n12794), .B2(n11948), .ZN(
        n5807) );
  OAI22_X1 U4021 ( .A1(n12797), .A2(n13321), .B1(n12794), .B2(n11949), .ZN(
        n5808) );
  OAI22_X1 U4022 ( .A1(n12797), .A2(n13324), .B1(n12794), .B2(n11950), .ZN(
        n5809) );
  OAI22_X1 U4023 ( .A1(n12797), .A2(n13327), .B1(n12794), .B2(n11951), .ZN(
        n5810) );
  OAI22_X1 U4024 ( .A1(n12797), .A2(n13330), .B1(n12794), .B2(n11952), .ZN(
        n5811) );
  OAI22_X1 U4025 ( .A1(n12796), .A2(n13333), .B1(n12794), .B2(n11953), .ZN(
        n5812) );
  OAI22_X1 U4026 ( .A1(n12796), .A2(n13336), .B1(n12794), .B2(n11954), .ZN(
        n5813) );
  OAI22_X1 U4027 ( .A1(n12796), .A2(n13339), .B1(n12794), .B2(n11955), .ZN(
        n5814) );
  OAI22_X1 U4028 ( .A1(n12796), .A2(n13342), .B1(n12794), .B2(n11956), .ZN(
        n5815) );
  OAI22_X1 U4029 ( .A1(n12796), .A2(n13345), .B1(n12794), .B2(n11957), .ZN(
        n5816) );
  OAI22_X1 U4030 ( .A1(n12795), .A2(n13348), .B1(n12794), .B2(n11958), .ZN(
        n5817) );
  OAI22_X1 U4031 ( .A1(n12822), .A2(n13243), .B1(n12812), .B2(n12093), .ZN(
        n5846) );
  OAI22_X1 U4032 ( .A1(n12822), .A2(n13246), .B1(n12812), .B2(n12094), .ZN(
        n5847) );
  OAI22_X1 U4033 ( .A1(n12822), .A2(n13249), .B1(n12812), .B2(n12095), .ZN(
        n5848) );
  OAI22_X1 U4034 ( .A1(n12822), .A2(n13252), .B1(n12812), .B2(n12096), .ZN(
        n5849) );
  OAI22_X1 U4035 ( .A1(n12822), .A2(n13255), .B1(n12812), .B2(n12097), .ZN(
        n5850) );
  OAI22_X1 U4036 ( .A1(n12821), .A2(n13258), .B1(n12812), .B2(n12098), .ZN(
        n5851) );
  OAI22_X1 U4037 ( .A1(n12821), .A2(n13261), .B1(n12812), .B2(n12099), .ZN(
        n5852) );
  OAI22_X1 U4038 ( .A1(n12821), .A2(n13264), .B1(n12812), .B2(n12100), .ZN(
        n5853) );
  OAI22_X1 U4039 ( .A1(n12821), .A2(n13267), .B1(n12812), .B2(n12101), .ZN(
        n5854) );
  OAI22_X1 U4040 ( .A1(n12821), .A2(n13270), .B1(n12812), .B2(n12102), .ZN(
        n5855) );
  OAI22_X1 U4041 ( .A1(n12820), .A2(n13273), .B1(n12812), .B2(n12103), .ZN(
        n5856) );
  OAI22_X1 U4042 ( .A1(n12820), .A2(n13276), .B1(n12812), .B2(n12104), .ZN(
        n5857) );
  OAI22_X1 U4043 ( .A1(n12820), .A2(n13279), .B1(n12813), .B2(n12105), .ZN(
        n5858) );
  OAI22_X1 U4044 ( .A1(n12820), .A2(n13282), .B1(n12813), .B2(n12106), .ZN(
        n5859) );
  OAI22_X1 U4045 ( .A1(n12820), .A2(n13285), .B1(n12813), .B2(n12107), .ZN(
        n5860) );
  OAI22_X1 U4046 ( .A1(n12819), .A2(n13288), .B1(n12813), .B2(n12108), .ZN(
        n5861) );
  OAI22_X1 U4047 ( .A1(n12819), .A2(n13291), .B1(n12813), .B2(n12109), .ZN(
        n5862) );
  OAI22_X1 U4048 ( .A1(n12819), .A2(n13294), .B1(n12813), .B2(n12110), .ZN(
        n5863) );
  OAI22_X1 U4049 ( .A1(n12819), .A2(n13297), .B1(n12813), .B2(n12111), .ZN(
        n5864) );
  OAI22_X1 U4050 ( .A1(n12819), .A2(n13300), .B1(n12813), .B2(n12112), .ZN(
        n5865) );
  OAI22_X1 U4051 ( .A1(n12818), .A2(n13303), .B1(n12813), .B2(n12113), .ZN(
        n5866) );
  OAI22_X1 U4052 ( .A1(n12818), .A2(n13306), .B1(n12813), .B2(n12114), .ZN(
        n5867) );
  OAI22_X1 U4053 ( .A1(n12818), .A2(n13309), .B1(n12813), .B2(n12115), .ZN(
        n5868) );
  OAI22_X1 U4054 ( .A1(n12818), .A2(n13312), .B1(n12813), .B2(n12116), .ZN(
        n5869) );
  OAI22_X1 U4055 ( .A1(n12818), .A2(n13315), .B1(n12814), .B2(n12117), .ZN(
        n5870) );
  OAI22_X1 U4056 ( .A1(n12817), .A2(n13318), .B1(n12814), .B2(n12118), .ZN(
        n5871) );
  OAI22_X1 U4057 ( .A1(n12817), .A2(n13321), .B1(n12814), .B2(n12119), .ZN(
        n5872) );
  OAI22_X1 U4058 ( .A1(n12817), .A2(n13324), .B1(n12814), .B2(n12120), .ZN(
        n5873) );
  OAI22_X1 U4059 ( .A1(n12817), .A2(n13327), .B1(n12814), .B2(n12121), .ZN(
        n5874) );
  OAI22_X1 U4060 ( .A1(n12817), .A2(n13330), .B1(n12814), .B2(n12122), .ZN(
        n5875) );
  OAI22_X1 U4061 ( .A1(n12816), .A2(n13333), .B1(n12814), .B2(n12123), .ZN(
        n5876) );
  OAI22_X1 U4062 ( .A1(n12816), .A2(n13336), .B1(n12814), .B2(n12124), .ZN(
        n5877) );
  OAI22_X1 U4063 ( .A1(n12816), .A2(n13339), .B1(n12814), .B2(n12125), .ZN(
        n5878) );
  OAI22_X1 U4064 ( .A1(n12816), .A2(n13342), .B1(n12814), .B2(n12126), .ZN(
        n5879) );
  OAI22_X1 U4065 ( .A1(n12816), .A2(n13345), .B1(n12814), .B2(n12127), .ZN(
        n5880) );
  OAI22_X1 U4066 ( .A1(n12815), .A2(n13348), .B1(n12814), .B2(n12128), .ZN(
        n5881) );
  OAI22_X1 U4067 ( .A1(n8515), .A2(n12551), .B1(n12571), .B2(n13184), .ZN(
        n4994) );
  OAI22_X1 U4068 ( .A1(n8498), .A2(n12551), .B1(n12571), .B2(n13187), .ZN(
        n4995) );
  OAI22_X1 U4069 ( .A1(n8481), .A2(n12551), .B1(n12571), .B2(n13190), .ZN(
        n4996) );
  OAI22_X1 U4070 ( .A1(n8464), .A2(n12551), .B1(n12571), .B2(n13193), .ZN(
        n4997) );
  OAI22_X1 U4071 ( .A1(n8447), .A2(n12551), .B1(n12570), .B2(n13196), .ZN(
        n4998) );
  OAI22_X1 U4072 ( .A1(n8430), .A2(n12551), .B1(n12570), .B2(n13199), .ZN(
        n4999) );
  OAI22_X1 U4073 ( .A1(n8413), .A2(n12551), .B1(n12570), .B2(n13202), .ZN(
        n5000) );
  OAI22_X1 U4074 ( .A1(n8396), .A2(n12551), .B1(n12570), .B2(n13205), .ZN(
        n5001) );
  OAI22_X1 U4075 ( .A1(n8379), .A2(n12552), .B1(n12569), .B2(n13208), .ZN(
        n5002) );
  OAI22_X1 U4076 ( .A1(n8362), .A2(n12552), .B1(n12569), .B2(n13211), .ZN(
        n5003) );
  OAI22_X1 U4077 ( .A1(n8345), .A2(n12552), .B1(n12569), .B2(n13214), .ZN(
        n5004) );
  OAI22_X1 U4078 ( .A1(n8328), .A2(n12552), .B1(n12569), .B2(n13217), .ZN(
        n5005) );
  OAI22_X1 U4079 ( .A1(n8311), .A2(n12552), .B1(n12568), .B2(n13220), .ZN(
        n5006) );
  OAI22_X1 U4080 ( .A1(n8294), .A2(n12552), .B1(n12568), .B2(n13223), .ZN(
        n5007) );
  OAI22_X1 U4081 ( .A1(n8277), .A2(n12552), .B1(n12568), .B2(n13226), .ZN(
        n5008) );
  OAI22_X1 U4082 ( .A1(n8260), .A2(n12552), .B1(n12568), .B2(n13229), .ZN(
        n5009) );
  OAI22_X1 U4083 ( .A1(n8243), .A2(n12552), .B1(n12567), .B2(n13232), .ZN(
        n5010) );
  OAI22_X1 U4084 ( .A1(n8226), .A2(n12552), .B1(n12567), .B2(n13235), .ZN(
        n5011) );
  OAI22_X1 U4085 ( .A1(n8209), .A2(n12552), .B1(n12567), .B2(n13238), .ZN(
        n5012) );
  OAI22_X1 U4086 ( .A1(n8192), .A2(n12552), .B1(n12567), .B2(n13241), .ZN(
        n5013) );
  OAI22_X1 U4087 ( .A1(n8175), .A2(n12553), .B1(n12566), .B2(n13244), .ZN(
        n5014) );
  OAI22_X1 U4088 ( .A1(n8158), .A2(n12553), .B1(n12566), .B2(n13247), .ZN(
        n5015) );
  OAI22_X1 U4089 ( .A1(n8141), .A2(n12553), .B1(n12566), .B2(n13250), .ZN(
        n5016) );
  OAI22_X1 U4090 ( .A1(n8124), .A2(n12553), .B1(n12566), .B2(n13253), .ZN(
        n5017) );
  OAI22_X1 U4091 ( .A1(n8107), .A2(n12553), .B1(n12565), .B2(n13256), .ZN(
        n5018) );
  OAI22_X1 U4092 ( .A1(n8090), .A2(n12553), .B1(n12565), .B2(n13259), .ZN(
        n5019) );
  OAI22_X1 U4093 ( .A1(n8073), .A2(n12553), .B1(n12565), .B2(n13262), .ZN(
        n5020) );
  OAI22_X1 U4094 ( .A1(n8056), .A2(n12553), .B1(n12565), .B2(n13265), .ZN(
        n5021) );
  OAI22_X1 U4095 ( .A1(n8039), .A2(n12553), .B1(n12564), .B2(n13268), .ZN(
        n5022) );
  OAI22_X1 U4096 ( .A1(n8022), .A2(n12553), .B1(n12564), .B2(n13271), .ZN(
        n5023) );
  OAI22_X1 U4097 ( .A1(n8005), .A2(n12553), .B1(n12564), .B2(n13274), .ZN(
        n5024) );
  OAI22_X1 U4098 ( .A1(n7988), .A2(n12553), .B1(n12564), .B2(n13277), .ZN(
        n5025) );
  OAI22_X1 U4099 ( .A1(n7971), .A2(n12554), .B1(n12563), .B2(n13280), .ZN(
        n5026) );
  OAI22_X1 U4100 ( .A1(n7954), .A2(n12554), .B1(n12563), .B2(n13283), .ZN(
        n5027) );
  OAI22_X1 U4101 ( .A1(n7937), .A2(n12554), .B1(n12563), .B2(n13286), .ZN(
        n5028) );
  OAI22_X1 U4102 ( .A1(n7920), .A2(n12554), .B1(n12563), .B2(n13289), .ZN(
        n5029) );
  OAI22_X1 U4103 ( .A1(n7903), .A2(n12554), .B1(n12562), .B2(n13292), .ZN(
        n5030) );
  OAI22_X1 U4104 ( .A1(n7886), .A2(n12554), .B1(n12562), .B2(n13295), .ZN(
        n5031) );
  OAI22_X1 U4105 ( .A1(n7869), .A2(n12554), .B1(n12562), .B2(n13298), .ZN(
        n5032) );
  OAI22_X1 U4106 ( .A1(n7852), .A2(n12554), .B1(n12562), .B2(n13301), .ZN(
        n5033) );
  OAI22_X1 U4107 ( .A1(n7835), .A2(n12554), .B1(n12561), .B2(n13304), .ZN(
        n5034) );
  OAI22_X1 U4108 ( .A1(n7818), .A2(n12554), .B1(n12561), .B2(n13307), .ZN(
        n5035) );
  OAI22_X1 U4109 ( .A1(n7801), .A2(n12554), .B1(n12561), .B2(n13310), .ZN(
        n5036) );
  OAI22_X1 U4110 ( .A1(n7784), .A2(n12554), .B1(n12561), .B2(n13313), .ZN(
        n5037) );
  OAI22_X1 U4111 ( .A1(n7767), .A2(n12555), .B1(n12560), .B2(n13316), .ZN(
        n5038) );
  OAI22_X1 U4112 ( .A1(n7750), .A2(n12555), .B1(n12560), .B2(n13319), .ZN(
        n5039) );
  OAI22_X1 U4113 ( .A1(n7648), .A2(n12555), .B1(n12560), .B2(n13322), .ZN(
        n5040) );
  OAI22_X1 U4114 ( .A1(n7631), .A2(n12555), .B1(n12560), .B2(n13325), .ZN(
        n5041) );
  OAI22_X1 U4115 ( .A1(n7527), .A2(n12555), .B1(n12559), .B2(n13328), .ZN(
        n5042) );
  OAI22_X1 U4116 ( .A1(n7510), .A2(n12555), .B1(n12559), .B2(n13331), .ZN(
        n5043) );
  OAI22_X1 U4117 ( .A1(n7493), .A2(n12555), .B1(n12559), .B2(n13334), .ZN(
        n5044) );
  OAI22_X1 U4118 ( .A1(n7391), .A2(n12555), .B1(n12559), .B2(n13337), .ZN(
        n5045) );
  OAI22_X1 U4119 ( .A1(n7374), .A2(n12555), .B1(n12558), .B2(n13340), .ZN(
        n5046) );
  OAI22_X1 U4120 ( .A1(n7275), .A2(n12555), .B1(n12558), .B2(n13343), .ZN(
        n5047) );
  OAI22_X1 U4121 ( .A1(n7258), .A2(n12555), .B1(n12558), .B2(n13346), .ZN(
        n5048) );
  OAI22_X1 U4122 ( .A1(n7241), .A2(n12555), .B1(n12558), .B2(n13349), .ZN(
        n5049) );
  OAI22_X1 U4123 ( .A1(n7144), .A2(n12556), .B1(n12557), .B2(n13352), .ZN(
        n5050) );
  OAI22_X1 U4124 ( .A1(n7127), .A2(n12556), .B1(n12557), .B2(n13355), .ZN(
        n5051) );
  OAI22_X1 U4125 ( .A1(n7110), .A2(n12556), .B1(n12557), .B2(n13358), .ZN(
        n5052) );
  OAI22_X1 U4126 ( .A1(n4849), .A2(n12556), .B1(n12557), .B2(n13381), .ZN(
        n5053) );
  OAI22_X1 U4127 ( .A1(n8583), .A2(n12551), .B1(n12572), .B2(n13172), .ZN(
        n4990) );
  OAI22_X1 U4128 ( .A1(n8566), .A2(n12551), .B1(n12572), .B2(n13175), .ZN(
        n4991) );
  OAI22_X1 U4129 ( .A1(n8549), .A2(n12551), .B1(n12572), .B2(n13178), .ZN(
        n4992) );
  OAI22_X1 U4130 ( .A1(n8532), .A2(n12551), .B1(n12572), .B2(n13181), .ZN(
        n4993) );
  OAI22_X1 U4131 ( .A1(n12927), .A2(n13171), .B1(n8575), .B2(n12911), .ZN(
        n6142) );
  OAI22_X1 U4132 ( .A1(n12927), .A2(n13174), .B1(n8558), .B2(n12911), .ZN(
        n6143) );
  OAI22_X1 U4133 ( .A1(n12927), .A2(n13177), .B1(n8541), .B2(n12911), .ZN(
        n6144) );
  OAI22_X1 U4134 ( .A1(n12927), .A2(n13180), .B1(n8524), .B2(n12911), .ZN(
        n6145) );
  OAI22_X1 U4135 ( .A1(n12926), .A2(n13183), .B1(n8507), .B2(n12911), .ZN(
        n6146) );
  OAI22_X1 U4136 ( .A1(n12926), .A2(n13186), .B1(n8490), .B2(n12911), .ZN(
        n6147) );
  OAI22_X1 U4137 ( .A1(n12926), .A2(n13189), .B1(n8473), .B2(n12911), .ZN(
        n6148) );
  OAI22_X1 U4138 ( .A1(n12926), .A2(n13192), .B1(n8456), .B2(n12911), .ZN(
        n6149) );
  OAI22_X1 U4139 ( .A1(n12926), .A2(n13195), .B1(n8439), .B2(n12911), .ZN(
        n6150) );
  OAI22_X1 U4140 ( .A1(n12925), .A2(n13198), .B1(n8422), .B2(n12911), .ZN(
        n6151) );
  OAI22_X1 U4141 ( .A1(n12925), .A2(n13201), .B1(n8405), .B2(n12911), .ZN(
        n6152) );
  OAI22_X1 U4142 ( .A1(n12925), .A2(n13204), .B1(n8388), .B2(n12911), .ZN(
        n6153) );
  OAI22_X1 U4143 ( .A1(n12925), .A2(n13207), .B1(n8371), .B2(n12913), .ZN(
        n6154) );
  OAI22_X1 U4144 ( .A1(n12925), .A2(n13210), .B1(n8354), .B2(n12914), .ZN(
        n6155) );
  OAI22_X1 U4145 ( .A1(n12924), .A2(n13213), .B1(n8337), .B2(n12911), .ZN(
        n6156) );
  OAI22_X1 U4146 ( .A1(n12924), .A2(n13216), .B1(n8320), .B2(n12913), .ZN(
        n6157) );
  OAI22_X1 U4147 ( .A1(n12924), .A2(n13219), .B1(n8303), .B2(n12914), .ZN(
        n6158) );
  OAI22_X1 U4148 ( .A1(n12924), .A2(n13222), .B1(n8286), .B2(n12910), .ZN(
        n6159) );
  OAI22_X1 U4149 ( .A1(n12924), .A2(n13225), .B1(n8269), .B2(n1929), .ZN(n6160) );
  OAI22_X1 U4150 ( .A1(n12923), .A2(n13228), .B1(n8252), .B2(n1929), .ZN(n6161) );
  OAI22_X1 U4151 ( .A1(n12923), .A2(n13231), .B1(n8235), .B2(n1929), .ZN(n6162) );
  OAI22_X1 U4152 ( .A1(n12923), .A2(n13234), .B1(n8218), .B2(n1929), .ZN(n6163) );
  OAI22_X1 U4153 ( .A1(n12923), .A2(n13237), .B1(n8201), .B2(n1929), .ZN(n6164) );
  OAI22_X1 U4154 ( .A1(n12923), .A2(n13240), .B1(n8184), .B2(n1929), .ZN(n6165) );
  OAI22_X1 U4155 ( .A1(n12593), .A2(n13172), .B1(n8584), .B2(n12578), .ZN(
        n5054) );
  OAI22_X1 U4156 ( .A1(n12593), .A2(n13175), .B1(n8567), .B2(n12577), .ZN(
        n5055) );
  OAI22_X1 U4157 ( .A1(n12593), .A2(n13178), .B1(n8550), .B2(n12577), .ZN(
        n5056) );
  OAI22_X1 U4158 ( .A1(n12592), .A2(n13184), .B1(n8516), .B2(n1948), .ZN(n5058) );
  OAI22_X1 U4159 ( .A1(n12593), .A2(n13181), .B1(n8533), .B2(n1948), .ZN(n5057) );
  OAI22_X1 U4160 ( .A1(n12592), .A2(n13187), .B1(n8499), .B2(n1948), .ZN(n5059) );
  OAI22_X1 U4161 ( .A1(n12592), .A2(n13190), .B1(n8482), .B2(n1948), .ZN(n5060) );
  OAI22_X1 U4162 ( .A1(n12592), .A2(n13193), .B1(n8465), .B2(n1948), .ZN(n5061) );
  OAI22_X1 U4163 ( .A1(n12592), .A2(n13196), .B1(n8448), .B2(n12577), .ZN(
        n5062) );
  OAI22_X1 U4164 ( .A1(n12591), .A2(n13199), .B1(n8431), .B2(n12577), .ZN(
        n5063) );
  OAI22_X1 U4165 ( .A1(n12591), .A2(n13202), .B1(n8414), .B2(n12577), .ZN(
        n5064) );
  OAI22_X1 U4166 ( .A1(n12591), .A2(n13205), .B1(n8397), .B2(n12577), .ZN(
        n5065) );
  OAI22_X1 U4167 ( .A1(n12591), .A2(n13208), .B1(n8380), .B2(n12579), .ZN(
        n5066) );
  OAI22_X1 U4168 ( .A1(n12591), .A2(n13211), .B1(n8363), .B2(n12580), .ZN(
        n5067) );
  OAI22_X1 U4169 ( .A1(n12590), .A2(n13214), .B1(n8346), .B2(n12578), .ZN(
        n5068) );
  OAI22_X1 U4170 ( .A1(n12590), .A2(n13217), .B1(n8329), .B2(n12579), .ZN(
        n5069) );
  OAI22_X1 U4171 ( .A1(n12590), .A2(n13220), .B1(n8312), .B2(n12580), .ZN(
        n5070) );
  OAI22_X1 U4172 ( .A1(n12590), .A2(n13223), .B1(n8295), .B2(n12577), .ZN(
        n5071) );
  OAI22_X1 U4173 ( .A1(n12590), .A2(n13226), .B1(n8278), .B2(n1948), .ZN(n5072) );
  OAI22_X1 U4174 ( .A1(n12589), .A2(n13229), .B1(n8261), .B2(n1948), .ZN(n5073) );
  OAI22_X1 U4175 ( .A1(n12589), .A2(n13232), .B1(n8244), .B2(n1948), .ZN(n5074) );
  OAI22_X1 U4176 ( .A1(n12589), .A2(n13235), .B1(n8227), .B2(n1948), .ZN(n5075) );
  OAI22_X1 U4177 ( .A1(n12589), .A2(n13238), .B1(n8210), .B2(n1948), .ZN(n5076) );
  OAI22_X1 U4178 ( .A1(n12589), .A2(n13241), .B1(n8193), .B2(n1948), .ZN(n5077) );
  OAI22_X1 U4179 ( .A1(n13007), .A2(n13170), .B1(n8573), .B2(n12991), .ZN(
        n6398) );
  OAI22_X1 U4180 ( .A1(n13007), .A2(n13173), .B1(n8556), .B2(n12991), .ZN(
        n6399) );
  OAI22_X1 U4181 ( .A1(n13007), .A2(n13176), .B1(n8539), .B2(n12991), .ZN(
        n6400) );
  OAI22_X1 U4182 ( .A1(n13007), .A2(n13179), .B1(n8522), .B2(n12991), .ZN(
        n6401) );
  OAI22_X1 U4183 ( .A1(n13006), .A2(n13182), .B1(n8505), .B2(n12991), .ZN(
        n6402) );
  OAI22_X1 U4184 ( .A1(n13006), .A2(n13185), .B1(n8488), .B2(n12991), .ZN(
        n6403) );
  OAI22_X1 U4185 ( .A1(n13006), .A2(n13188), .B1(n8471), .B2(n12991), .ZN(
        n6404) );
  OAI22_X1 U4186 ( .A1(n13006), .A2(n13191), .B1(n8454), .B2(n12991), .ZN(
        n6405) );
  OAI22_X1 U4187 ( .A1(n13006), .A2(n13194), .B1(n8437), .B2(n12991), .ZN(
        n6406) );
  OAI22_X1 U4188 ( .A1(n13005), .A2(n13197), .B1(n8420), .B2(n12991), .ZN(
        n6407) );
  OAI22_X1 U4189 ( .A1(n13005), .A2(n13200), .B1(n8403), .B2(n12991), .ZN(
        n6408) );
  OAI22_X1 U4190 ( .A1(n13005), .A2(n13203), .B1(n8386), .B2(n12991), .ZN(
        n6409) );
  OAI22_X1 U4191 ( .A1(n13005), .A2(n13206), .B1(n8369), .B2(n12993), .ZN(
        n6410) );
  OAI22_X1 U4192 ( .A1(n13005), .A2(n13209), .B1(n8352), .B2(n12994), .ZN(
        n6411) );
  OAI22_X1 U4193 ( .A1(n13004), .A2(n13212), .B1(n8335), .B2(n12991), .ZN(
        n6412) );
  OAI22_X1 U4194 ( .A1(n13004), .A2(n13215), .B1(n8318), .B2(n12993), .ZN(
        n6413) );
  OAI22_X1 U4195 ( .A1(n13004), .A2(n13218), .B1(n8301), .B2(n12994), .ZN(
        n6414) );
  OAI22_X1 U4196 ( .A1(n13004), .A2(n13221), .B1(n8284), .B2(n12990), .ZN(
        n6415) );
  OAI22_X1 U4197 ( .A1(n13004), .A2(n13224), .B1(n8267), .B2(n1925), .ZN(n6416) );
  OAI22_X1 U4198 ( .A1(n13003), .A2(n13227), .B1(n8250), .B2(n1925), .ZN(n6417) );
  OAI22_X1 U4199 ( .A1(n13003), .A2(n13230), .B1(n8233), .B2(n1925), .ZN(n6418) );
  OAI22_X1 U4200 ( .A1(n13003), .A2(n13233), .B1(n8216), .B2(n1925), .ZN(n6419) );
  OAI22_X1 U4201 ( .A1(n13003), .A2(n13236), .B1(n8199), .B2(n1925), .ZN(n6420) );
  OAI22_X1 U4202 ( .A1(n13003), .A2(n13239), .B1(n8182), .B2(n1925), .ZN(n6421) );
  OAI22_X1 U4203 ( .A1(n12847), .A2(n13171), .B1(n8577), .B2(n12831), .ZN(
        n5886) );
  OAI22_X1 U4204 ( .A1(n12847), .A2(n13174), .B1(n8560), .B2(n12831), .ZN(
        n5887) );
  OAI22_X1 U4205 ( .A1(n12847), .A2(n13177), .B1(n8543), .B2(n12831), .ZN(
        n5888) );
  OAI22_X1 U4206 ( .A1(n12847), .A2(n13180), .B1(n8526), .B2(n12831), .ZN(
        n5889) );
  OAI22_X1 U4207 ( .A1(n12846), .A2(n13183), .B1(n8509), .B2(n12831), .ZN(
        n5890) );
  OAI22_X1 U4208 ( .A1(n12846), .A2(n13186), .B1(n8492), .B2(n12831), .ZN(
        n5891) );
  OAI22_X1 U4209 ( .A1(n12846), .A2(n13189), .B1(n8475), .B2(n12831), .ZN(
        n5892) );
  OAI22_X1 U4210 ( .A1(n12846), .A2(n13192), .B1(n8458), .B2(n12831), .ZN(
        n5893) );
  OAI22_X1 U4211 ( .A1(n12846), .A2(n13195), .B1(n8441), .B2(n12831), .ZN(
        n5894) );
  OAI22_X1 U4212 ( .A1(n12845), .A2(n13198), .B1(n8424), .B2(n12831), .ZN(
        n5895) );
  OAI22_X1 U4213 ( .A1(n12845), .A2(n13201), .B1(n8407), .B2(n12831), .ZN(
        n5896) );
  OAI22_X1 U4214 ( .A1(n12845), .A2(n13204), .B1(n8390), .B2(n12831), .ZN(
        n5897) );
  OAI22_X1 U4215 ( .A1(n12845), .A2(n13207), .B1(n8373), .B2(n12833), .ZN(
        n5898) );
  OAI22_X1 U4216 ( .A1(n12845), .A2(n13210), .B1(n8356), .B2(n12834), .ZN(
        n5899) );
  OAI22_X1 U4217 ( .A1(n12844), .A2(n13213), .B1(n8339), .B2(n12831), .ZN(
        n5900) );
  OAI22_X1 U4218 ( .A1(n12844), .A2(n13216), .B1(n8322), .B2(n12833), .ZN(
        n5901) );
  OAI22_X1 U4219 ( .A1(n12844), .A2(n13219), .B1(n8305), .B2(n12834), .ZN(
        n5902) );
  OAI22_X1 U4220 ( .A1(n12844), .A2(n13222), .B1(n8288), .B2(n12830), .ZN(
        n5903) );
  OAI22_X1 U4221 ( .A1(n12844), .A2(n13225), .B1(n8271), .B2(n1934), .ZN(n5904) );
  OAI22_X1 U4222 ( .A1(n12843), .A2(n13228), .B1(n8254), .B2(n1934), .ZN(n5905) );
  OAI22_X1 U4223 ( .A1(n12843), .A2(n13231), .B1(n8237), .B2(n1934), .ZN(n5906) );
  OAI22_X1 U4224 ( .A1(n12843), .A2(n13234), .B1(n8220), .B2(n1934), .ZN(n5907) );
  OAI22_X1 U4225 ( .A1(n12843), .A2(n13237), .B1(n8203), .B2(n1934), .ZN(n5908) );
  OAI22_X1 U4226 ( .A1(n12843), .A2(n13240), .B1(n8186), .B2(n1934), .ZN(n5909) );
  OAI22_X1 U4227 ( .A1(n12787), .A2(n13171), .B1(n8580), .B2(n12771), .ZN(
        n5694) );
  OAI22_X1 U4228 ( .A1(n12787), .A2(n13174), .B1(n8563), .B2(n12771), .ZN(
        n5695) );
  OAI22_X1 U4229 ( .A1(n12787), .A2(n13177), .B1(n8546), .B2(n12771), .ZN(
        n5696) );
  OAI22_X1 U4230 ( .A1(n12787), .A2(n13180), .B1(n8529), .B2(n12771), .ZN(
        n5697) );
  OAI22_X1 U4231 ( .A1(n12786), .A2(n13183), .B1(n8512), .B2(n12771), .ZN(
        n5698) );
  OAI22_X1 U4232 ( .A1(n12786), .A2(n13186), .B1(n8495), .B2(n12771), .ZN(
        n5699) );
  OAI22_X1 U4233 ( .A1(n12786), .A2(n13189), .B1(n8478), .B2(n12771), .ZN(
        n5700) );
  OAI22_X1 U4234 ( .A1(n12786), .A2(n13192), .B1(n8461), .B2(n12771), .ZN(
        n5701) );
  OAI22_X1 U4235 ( .A1(n12786), .A2(n13195), .B1(n8444), .B2(n12771), .ZN(
        n5702) );
  OAI22_X1 U4236 ( .A1(n12785), .A2(n13198), .B1(n8427), .B2(n12771), .ZN(
        n5703) );
  OAI22_X1 U4237 ( .A1(n12785), .A2(n13201), .B1(n8410), .B2(n12771), .ZN(
        n5704) );
  OAI22_X1 U4238 ( .A1(n12785), .A2(n13204), .B1(n8393), .B2(n12771), .ZN(
        n5705) );
  OAI22_X1 U4239 ( .A1(n12785), .A2(n13207), .B1(n8376), .B2(n12773), .ZN(
        n5706) );
  OAI22_X1 U4240 ( .A1(n12785), .A2(n13210), .B1(n8359), .B2(n12774), .ZN(
        n5707) );
  OAI22_X1 U4241 ( .A1(n12784), .A2(n13213), .B1(n8342), .B2(n12771), .ZN(
        n5708) );
  OAI22_X1 U4242 ( .A1(n12784), .A2(n13216), .B1(n8325), .B2(n12773), .ZN(
        n5709) );
  OAI22_X1 U4243 ( .A1(n12784), .A2(n13219), .B1(n8308), .B2(n12774), .ZN(
        n5710) );
  OAI22_X1 U4244 ( .A1(n12784), .A2(n13222), .B1(n8291), .B2(n12770), .ZN(
        n5711) );
  OAI22_X1 U4245 ( .A1(n12784), .A2(n13225), .B1(n8274), .B2(n1937), .ZN(n5712) );
  OAI22_X1 U4246 ( .A1(n12783), .A2(n13228), .B1(n8257), .B2(n1937), .ZN(n5713) );
  OAI22_X1 U4247 ( .A1(n12783), .A2(n13231), .B1(n8240), .B2(n1937), .ZN(n5714) );
  OAI22_X1 U4248 ( .A1(n12783), .A2(n13234), .B1(n8223), .B2(n1937), .ZN(n5715) );
  OAI22_X1 U4249 ( .A1(n12783), .A2(n13237), .B1(n8206), .B2(n1937), .ZN(n5716) );
  OAI22_X1 U4250 ( .A1(n12783), .A2(n13240), .B1(n8189), .B2(n1937), .ZN(n5717) );
  OAI22_X1 U4251 ( .A1(n12767), .A2(n13171), .B1(n8579), .B2(n12751), .ZN(
        n5630) );
  OAI22_X1 U4252 ( .A1(n12767), .A2(n13174), .B1(n8562), .B2(n12751), .ZN(
        n5631) );
  OAI22_X1 U4253 ( .A1(n12767), .A2(n13177), .B1(n8545), .B2(n12751), .ZN(
        n5632) );
  OAI22_X1 U4254 ( .A1(n12767), .A2(n13180), .B1(n8528), .B2(n12751), .ZN(
        n5633) );
  OAI22_X1 U4255 ( .A1(n12766), .A2(n13183), .B1(n8511), .B2(n12751), .ZN(
        n5634) );
  OAI22_X1 U4256 ( .A1(n12766), .A2(n13186), .B1(n8494), .B2(n12751), .ZN(
        n5635) );
  OAI22_X1 U4257 ( .A1(n12766), .A2(n13189), .B1(n8477), .B2(n12751), .ZN(
        n5636) );
  OAI22_X1 U4258 ( .A1(n12766), .A2(n13192), .B1(n8460), .B2(n12751), .ZN(
        n5637) );
  OAI22_X1 U4259 ( .A1(n12766), .A2(n13195), .B1(n8443), .B2(n12751), .ZN(
        n5638) );
  OAI22_X1 U4260 ( .A1(n12765), .A2(n13198), .B1(n8426), .B2(n12751), .ZN(
        n5639) );
  OAI22_X1 U4261 ( .A1(n12765), .A2(n13201), .B1(n8409), .B2(n12751), .ZN(
        n5640) );
  OAI22_X1 U4262 ( .A1(n12765), .A2(n13204), .B1(n8392), .B2(n12751), .ZN(
        n5641) );
  OAI22_X1 U4263 ( .A1(n12765), .A2(n13207), .B1(n8375), .B2(n12753), .ZN(
        n5642) );
  OAI22_X1 U4264 ( .A1(n12765), .A2(n13210), .B1(n8358), .B2(n12754), .ZN(
        n5643) );
  OAI22_X1 U4265 ( .A1(n12764), .A2(n13213), .B1(n8341), .B2(n12751), .ZN(
        n5644) );
  OAI22_X1 U4266 ( .A1(n12764), .A2(n13216), .B1(n8324), .B2(n12753), .ZN(
        n5645) );
  OAI22_X1 U4267 ( .A1(n12764), .A2(n13219), .B1(n8307), .B2(n12754), .ZN(
        n5646) );
  OAI22_X1 U4268 ( .A1(n12764), .A2(n13222), .B1(n8290), .B2(n12750), .ZN(
        n5647) );
  OAI22_X1 U4269 ( .A1(n12764), .A2(n13225), .B1(n8273), .B2(n1938), .ZN(n5648) );
  OAI22_X1 U4270 ( .A1(n12763), .A2(n13228), .B1(n8256), .B2(n1938), .ZN(n5649) );
  OAI22_X1 U4271 ( .A1(n12763), .A2(n13231), .B1(n8239), .B2(n1938), .ZN(n5650) );
  OAI22_X1 U4272 ( .A1(n12763), .A2(n13234), .B1(n8222), .B2(n1938), .ZN(n5651) );
  OAI22_X1 U4273 ( .A1(n12763), .A2(n13237), .B1(n8205), .B2(n1938), .ZN(n5652) );
  OAI22_X1 U4274 ( .A1(n12763), .A2(n13240), .B1(n8188), .B2(n1938), .ZN(n5653) );
  OAI22_X1 U4275 ( .A1(n12650), .A2(n13172), .B1(n8581), .B2(n12635), .ZN(
        n5246) );
  OAI22_X1 U4276 ( .A1(n12669), .A2(n13172), .B1(n8582), .B2(n12654), .ZN(
        n5310) );
  OAI22_X1 U4277 ( .A1(n12650), .A2(n13175), .B1(n8564), .B2(n12634), .ZN(
        n5247) );
  OAI22_X1 U4278 ( .A1(n12650), .A2(n13178), .B1(n8547), .B2(n12634), .ZN(
        n5248) );
  OAI22_X1 U4279 ( .A1(n12649), .A2(n13184), .B1(n8513), .B2(n1945), .ZN(n5250) );
  OAI22_X1 U4280 ( .A1(n12650), .A2(n13181), .B1(n8530), .B2(n1945), .ZN(n5249) );
  OAI22_X1 U4281 ( .A1(n12649), .A2(n13187), .B1(n8496), .B2(n1945), .ZN(n5251) );
  OAI22_X1 U4282 ( .A1(n12649), .A2(n13190), .B1(n8479), .B2(n1945), .ZN(n5252) );
  OAI22_X1 U4283 ( .A1(n12649), .A2(n13193), .B1(n8462), .B2(n1945), .ZN(n5253) );
  OAI22_X1 U4284 ( .A1(n12649), .A2(n13196), .B1(n8445), .B2(n12634), .ZN(
        n5254) );
  OAI22_X1 U4285 ( .A1(n12648), .A2(n13199), .B1(n8428), .B2(n12634), .ZN(
        n5255) );
  OAI22_X1 U4286 ( .A1(n12648), .A2(n13202), .B1(n8411), .B2(n12634), .ZN(
        n5256) );
  OAI22_X1 U4287 ( .A1(n12648), .A2(n13205), .B1(n8394), .B2(n12634), .ZN(
        n5257) );
  OAI22_X1 U4288 ( .A1(n12648), .A2(n13208), .B1(n8377), .B2(n12636), .ZN(
        n5258) );
  OAI22_X1 U4289 ( .A1(n12648), .A2(n13211), .B1(n8360), .B2(n12637), .ZN(
        n5259) );
  OAI22_X1 U4290 ( .A1(n12647), .A2(n13214), .B1(n8343), .B2(n12635), .ZN(
        n5260) );
  OAI22_X1 U4291 ( .A1(n12647), .A2(n13217), .B1(n8326), .B2(n12636), .ZN(
        n5261) );
  OAI22_X1 U4292 ( .A1(n12647), .A2(n13220), .B1(n8309), .B2(n12637), .ZN(
        n5262) );
  OAI22_X1 U4293 ( .A1(n12647), .A2(n13223), .B1(n8292), .B2(n12634), .ZN(
        n5263) );
  OAI22_X1 U4294 ( .A1(n12647), .A2(n13226), .B1(n8275), .B2(n1945), .ZN(n5264) );
  OAI22_X1 U4295 ( .A1(n12646), .A2(n13229), .B1(n8258), .B2(n1945), .ZN(n5265) );
  OAI22_X1 U4296 ( .A1(n12646), .A2(n13232), .B1(n8241), .B2(n1945), .ZN(n5266) );
  OAI22_X1 U4297 ( .A1(n12646), .A2(n13235), .B1(n8224), .B2(n1945), .ZN(n5267) );
  OAI22_X1 U4298 ( .A1(n12646), .A2(n13238), .B1(n8207), .B2(n1945), .ZN(n5268) );
  OAI22_X1 U4299 ( .A1(n12646), .A2(n13241), .B1(n8190), .B2(n1945), .ZN(n5269) );
  OAI22_X1 U4300 ( .A1(n12669), .A2(n13175), .B1(n8565), .B2(n12653), .ZN(
        n5311) );
  OAI22_X1 U4301 ( .A1(n12669), .A2(n13178), .B1(n8548), .B2(n12653), .ZN(
        n5312) );
  OAI22_X1 U4302 ( .A1(n12668), .A2(n13184), .B1(n8514), .B2(n1944), .ZN(n5314) );
  OAI22_X1 U4303 ( .A1(n12669), .A2(n13181), .B1(n8531), .B2(n1944), .ZN(n5313) );
  OAI22_X1 U4304 ( .A1(n12668), .A2(n13187), .B1(n8497), .B2(n1944), .ZN(n5315) );
  OAI22_X1 U4305 ( .A1(n12668), .A2(n13190), .B1(n8480), .B2(n1944), .ZN(n5316) );
  OAI22_X1 U4306 ( .A1(n12668), .A2(n13193), .B1(n8463), .B2(n1944), .ZN(n5317) );
  OAI22_X1 U4307 ( .A1(n12668), .A2(n13196), .B1(n8446), .B2(n12653), .ZN(
        n5318) );
  OAI22_X1 U4308 ( .A1(n12667), .A2(n13199), .B1(n8429), .B2(n12653), .ZN(
        n5319) );
  OAI22_X1 U4309 ( .A1(n12667), .A2(n13202), .B1(n8412), .B2(n12653), .ZN(
        n5320) );
  OAI22_X1 U4310 ( .A1(n12667), .A2(n13205), .B1(n8395), .B2(n12653), .ZN(
        n5321) );
  OAI22_X1 U4311 ( .A1(n12667), .A2(n13208), .B1(n8378), .B2(n12655), .ZN(
        n5322) );
  OAI22_X1 U4312 ( .A1(n12667), .A2(n13211), .B1(n8361), .B2(n12656), .ZN(
        n5323) );
  OAI22_X1 U4313 ( .A1(n12666), .A2(n13214), .B1(n8344), .B2(n12654), .ZN(
        n5324) );
  OAI22_X1 U4314 ( .A1(n12666), .A2(n13217), .B1(n8327), .B2(n12655), .ZN(
        n5325) );
  OAI22_X1 U4315 ( .A1(n12666), .A2(n13220), .B1(n8310), .B2(n12656), .ZN(
        n5326) );
  OAI22_X1 U4316 ( .A1(n12666), .A2(n13223), .B1(n8293), .B2(n12653), .ZN(
        n5327) );
  OAI22_X1 U4317 ( .A1(n12666), .A2(n13226), .B1(n8276), .B2(n1944), .ZN(n5328) );
  OAI22_X1 U4318 ( .A1(n12665), .A2(n13229), .B1(n8259), .B2(n1944), .ZN(n5329) );
  OAI22_X1 U4319 ( .A1(n12665), .A2(n13232), .B1(n8242), .B2(n1944), .ZN(n5330) );
  OAI22_X1 U4320 ( .A1(n12665), .A2(n13235), .B1(n8225), .B2(n1944), .ZN(n5331) );
  OAI22_X1 U4321 ( .A1(n12665), .A2(n13238), .B1(n8208), .B2(n1944), .ZN(n5332) );
  OAI22_X1 U4322 ( .A1(n12665), .A2(n13241), .B1(n8191), .B2(n1944), .ZN(n5333) );
  OAI22_X1 U4323 ( .A1(n13025), .A2(n13206), .B1(n8370), .B2(n13011), .ZN(
        n6474) );
  OAI22_X1 U4324 ( .A1(n13025), .A2(n13209), .B1(n8353), .B2(n13011), .ZN(
        n6475) );
  OAI22_X1 U4325 ( .A1(n13024), .A2(n13212), .B1(n8336), .B2(n13011), .ZN(
        n6476) );
  OAI22_X1 U4326 ( .A1(n13024), .A2(n13215), .B1(n8319), .B2(n13011), .ZN(
        n6477) );
  OAI22_X1 U4327 ( .A1(n13024), .A2(n13218), .B1(n8302), .B2(n13011), .ZN(
        n6478) );
  OAI22_X1 U4328 ( .A1(n13024), .A2(n13221), .B1(n8285), .B2(n13011), .ZN(
        n6479) );
  OAI22_X1 U4329 ( .A1(n13024), .A2(n13224), .B1(n8268), .B2(n13011), .ZN(
        n6480) );
  OAI22_X1 U4330 ( .A1(n13023), .A2(n13227), .B1(n8251), .B2(n13011), .ZN(
        n6481) );
  OAI22_X1 U4331 ( .A1(n13023), .A2(n13230), .B1(n8234), .B2(n13011), .ZN(
        n6482) );
  OAI22_X1 U4332 ( .A1(n13023), .A2(n13233), .B1(n8217), .B2(n13011), .ZN(
        n6483) );
  OAI22_X1 U4333 ( .A1(n13023), .A2(n13236), .B1(n8200), .B2(n13011), .ZN(
        n6484) );
  OAI22_X1 U4334 ( .A1(n13023), .A2(n13239), .B1(n8183), .B2(n13011), .ZN(
        n6485) );
  OAI22_X1 U4335 ( .A1(n13065), .A2(n13206), .B1(n8367), .B2(n13051), .ZN(
        n6602) );
  OAI22_X1 U4336 ( .A1(n13065), .A2(n13209), .B1(n8350), .B2(n13051), .ZN(
        n6603) );
  OAI22_X1 U4337 ( .A1(n13064), .A2(n13212), .B1(n8333), .B2(n13051), .ZN(
        n6604) );
  OAI22_X1 U4338 ( .A1(n13064), .A2(n13215), .B1(n8316), .B2(n13051), .ZN(
        n6605) );
  OAI22_X1 U4339 ( .A1(n13064), .A2(n13218), .B1(n8299), .B2(n13051), .ZN(
        n6606) );
  OAI22_X1 U4340 ( .A1(n13064), .A2(n13221), .B1(n8282), .B2(n13051), .ZN(
        n6607) );
  OAI22_X1 U4341 ( .A1(n13064), .A2(n13224), .B1(n8265), .B2(n13051), .ZN(
        n6608) );
  OAI22_X1 U4342 ( .A1(n13063), .A2(n13227), .B1(n8248), .B2(n13051), .ZN(
        n6609) );
  OAI22_X1 U4343 ( .A1(n13063), .A2(n13230), .B1(n8231), .B2(n13051), .ZN(
        n6610) );
  OAI22_X1 U4344 ( .A1(n13063), .A2(n13233), .B1(n8214), .B2(n13051), .ZN(
        n6611) );
  OAI22_X1 U4345 ( .A1(n13063), .A2(n13236), .B1(n8197), .B2(n13051), .ZN(
        n6612) );
  OAI22_X1 U4346 ( .A1(n13063), .A2(n13239), .B1(n8180), .B2(n13051), .ZN(
        n6613) );
  OAI22_X1 U4347 ( .A1(n13045), .A2(n13206), .B1(n8368), .B2(n13031), .ZN(
        n6538) );
  OAI22_X1 U4348 ( .A1(n13045), .A2(n13209), .B1(n8351), .B2(n13031), .ZN(
        n6539) );
  OAI22_X1 U4349 ( .A1(n13044), .A2(n13212), .B1(n8334), .B2(n13031), .ZN(
        n6540) );
  OAI22_X1 U4350 ( .A1(n13044), .A2(n13215), .B1(n8317), .B2(n13031), .ZN(
        n6541) );
  OAI22_X1 U4351 ( .A1(n13044), .A2(n13218), .B1(n8300), .B2(n13031), .ZN(
        n6542) );
  OAI22_X1 U4352 ( .A1(n13044), .A2(n13221), .B1(n8283), .B2(n13031), .ZN(
        n6543) );
  OAI22_X1 U4353 ( .A1(n13044), .A2(n13224), .B1(n8266), .B2(n13031), .ZN(
        n6544) );
  OAI22_X1 U4354 ( .A1(n13043), .A2(n13227), .B1(n8249), .B2(n13031), .ZN(
        n6545) );
  OAI22_X1 U4355 ( .A1(n13043), .A2(n13230), .B1(n8232), .B2(n13031), .ZN(
        n6546) );
  OAI22_X1 U4356 ( .A1(n13043), .A2(n13233), .B1(n8215), .B2(n13031), .ZN(
        n6547) );
  OAI22_X1 U4357 ( .A1(n13043), .A2(n13236), .B1(n8198), .B2(n13031), .ZN(
        n6548) );
  OAI22_X1 U4358 ( .A1(n13043), .A2(n13239), .B1(n8181), .B2(n13031), .ZN(
        n6549) );
  OAI22_X1 U4359 ( .A1(n12922), .A2(n13243), .B1(n8167), .B2(n12912), .ZN(
        n6166) );
  OAI22_X1 U4360 ( .A1(n12922), .A2(n13246), .B1(n8150), .B2(n12912), .ZN(
        n6167) );
  OAI22_X1 U4361 ( .A1(n12922), .A2(n13249), .B1(n8133), .B2(n12912), .ZN(
        n6168) );
  OAI22_X1 U4362 ( .A1(n12922), .A2(n13252), .B1(n8116), .B2(n12912), .ZN(
        n6169) );
  OAI22_X1 U4363 ( .A1(n12922), .A2(n13255), .B1(n8099), .B2(n12912), .ZN(
        n6170) );
  OAI22_X1 U4364 ( .A1(n12921), .A2(n13258), .B1(n8082), .B2(n12912), .ZN(
        n6171) );
  OAI22_X1 U4365 ( .A1(n12921), .A2(n13261), .B1(n8065), .B2(n12912), .ZN(
        n6172) );
  OAI22_X1 U4366 ( .A1(n12921), .A2(n13264), .B1(n8048), .B2(n12912), .ZN(
        n6173) );
  OAI22_X1 U4367 ( .A1(n12921), .A2(n13267), .B1(n8031), .B2(n12912), .ZN(
        n6174) );
  OAI22_X1 U4368 ( .A1(n12921), .A2(n13270), .B1(n8014), .B2(n12912), .ZN(
        n6175) );
  OAI22_X1 U4369 ( .A1(n12920), .A2(n13273), .B1(n7997), .B2(n12912), .ZN(
        n6176) );
  OAI22_X1 U4370 ( .A1(n12920), .A2(n13276), .B1(n7980), .B2(n12912), .ZN(
        n6177) );
  OAI22_X1 U4371 ( .A1(n12920), .A2(n13279), .B1(n7963), .B2(n12913), .ZN(
        n6178) );
  OAI22_X1 U4372 ( .A1(n12920), .A2(n13282), .B1(n7946), .B2(n12913), .ZN(
        n6179) );
  OAI22_X1 U4373 ( .A1(n12920), .A2(n13285), .B1(n7929), .B2(n12913), .ZN(
        n6180) );
  OAI22_X1 U4374 ( .A1(n12919), .A2(n13288), .B1(n7912), .B2(n12913), .ZN(
        n6181) );
  OAI22_X1 U4375 ( .A1(n12919), .A2(n13291), .B1(n7895), .B2(n12913), .ZN(
        n6182) );
  OAI22_X1 U4376 ( .A1(n12919), .A2(n13294), .B1(n7878), .B2(n12913), .ZN(
        n6183) );
  OAI22_X1 U4377 ( .A1(n12919), .A2(n13297), .B1(n7861), .B2(n12913), .ZN(
        n6184) );
  OAI22_X1 U4378 ( .A1(n12919), .A2(n13300), .B1(n7844), .B2(n12913), .ZN(
        n6185) );
  OAI22_X1 U4379 ( .A1(n12918), .A2(n13303), .B1(n7827), .B2(n12913), .ZN(
        n6186) );
  OAI22_X1 U4380 ( .A1(n12918), .A2(n13306), .B1(n7810), .B2(n12913), .ZN(
        n6187) );
  OAI22_X1 U4381 ( .A1(n12918), .A2(n13309), .B1(n7793), .B2(n12913), .ZN(
        n6188) );
  OAI22_X1 U4382 ( .A1(n12918), .A2(n13312), .B1(n7776), .B2(n12913), .ZN(
        n6189) );
  OAI22_X1 U4383 ( .A1(n12918), .A2(n13315), .B1(n7759), .B2(n12914), .ZN(
        n6190) );
  OAI22_X1 U4384 ( .A1(n12917), .A2(n13318), .B1(n7742), .B2(n12914), .ZN(
        n6191) );
  OAI22_X1 U4385 ( .A1(n12917), .A2(n13321), .B1(n7640), .B2(n12914), .ZN(
        n6192) );
  OAI22_X1 U4386 ( .A1(n12917), .A2(n13324), .B1(n7623), .B2(n12914), .ZN(
        n6193) );
  OAI22_X1 U4387 ( .A1(n12917), .A2(n13327), .B1(n7519), .B2(n12914), .ZN(
        n6194) );
  OAI22_X1 U4388 ( .A1(n12917), .A2(n13330), .B1(n7502), .B2(n12914), .ZN(
        n6195) );
  OAI22_X1 U4389 ( .A1(n12916), .A2(n13333), .B1(n7400), .B2(n12914), .ZN(
        n6196) );
  OAI22_X1 U4390 ( .A1(n12916), .A2(n13336), .B1(n7383), .B2(n12914), .ZN(
        n6197) );
  OAI22_X1 U4391 ( .A1(n12916), .A2(n13339), .B1(n7366), .B2(n12914), .ZN(
        n6198) );
  OAI22_X1 U4392 ( .A1(n12916), .A2(n13342), .B1(n7267), .B2(n12914), .ZN(
        n6199) );
  OAI22_X1 U4393 ( .A1(n12916), .A2(n13345), .B1(n7250), .B2(n12914), .ZN(
        n6200) );
  OAI22_X1 U4394 ( .A1(n12915), .A2(n13348), .B1(n7153), .B2(n12914), .ZN(
        n6201) );
  OAI22_X1 U4395 ( .A1(n12942), .A2(n13243), .B1(n8168), .B2(n12932), .ZN(
        n6230) );
  OAI22_X1 U4396 ( .A1(n12942), .A2(n13246), .B1(n8151), .B2(n12932), .ZN(
        n6231) );
  OAI22_X1 U4397 ( .A1(n12942), .A2(n13249), .B1(n8134), .B2(n12932), .ZN(
        n6232) );
  OAI22_X1 U4398 ( .A1(n12942), .A2(n13252), .B1(n8117), .B2(n12932), .ZN(
        n6233) );
  OAI22_X1 U4399 ( .A1(n12942), .A2(n13255), .B1(n8100), .B2(n12932), .ZN(
        n6234) );
  OAI22_X1 U4400 ( .A1(n12941), .A2(n13258), .B1(n8083), .B2(n12932), .ZN(
        n6235) );
  OAI22_X1 U4401 ( .A1(n12941), .A2(n13261), .B1(n8066), .B2(n12932), .ZN(
        n6236) );
  OAI22_X1 U4402 ( .A1(n12941), .A2(n13264), .B1(n8049), .B2(n12932), .ZN(
        n6237) );
  OAI22_X1 U4403 ( .A1(n12941), .A2(n13267), .B1(n8032), .B2(n12932), .ZN(
        n6238) );
  OAI22_X1 U4404 ( .A1(n12941), .A2(n13270), .B1(n8015), .B2(n12932), .ZN(
        n6239) );
  OAI22_X1 U4405 ( .A1(n12940), .A2(n13273), .B1(n7998), .B2(n12932), .ZN(
        n6240) );
  OAI22_X1 U4406 ( .A1(n12940), .A2(n13276), .B1(n7981), .B2(n12932), .ZN(
        n6241) );
  OAI22_X1 U4407 ( .A1(n12940), .A2(n13279), .B1(n7964), .B2(n12933), .ZN(
        n6242) );
  OAI22_X1 U4408 ( .A1(n12940), .A2(n13282), .B1(n7947), .B2(n12933), .ZN(
        n6243) );
  OAI22_X1 U4409 ( .A1(n12940), .A2(n13285), .B1(n7930), .B2(n12933), .ZN(
        n6244) );
  OAI22_X1 U4410 ( .A1(n12939), .A2(n13288), .B1(n7913), .B2(n12933), .ZN(
        n6245) );
  OAI22_X1 U4411 ( .A1(n12939), .A2(n13291), .B1(n7896), .B2(n12933), .ZN(
        n6246) );
  OAI22_X1 U4412 ( .A1(n12939), .A2(n13294), .B1(n7879), .B2(n12933), .ZN(
        n6247) );
  OAI22_X1 U4413 ( .A1(n12939), .A2(n13297), .B1(n7862), .B2(n12933), .ZN(
        n6248) );
  OAI22_X1 U4414 ( .A1(n12939), .A2(n13300), .B1(n7845), .B2(n12933), .ZN(
        n6249) );
  OAI22_X1 U4415 ( .A1(n12938), .A2(n13303), .B1(n7828), .B2(n12933), .ZN(
        n6250) );
  OAI22_X1 U4416 ( .A1(n12938), .A2(n13306), .B1(n7811), .B2(n12933), .ZN(
        n6251) );
  OAI22_X1 U4417 ( .A1(n12938), .A2(n13309), .B1(n7794), .B2(n12933), .ZN(
        n6252) );
  OAI22_X1 U4418 ( .A1(n12938), .A2(n13312), .B1(n7777), .B2(n12933), .ZN(
        n6253) );
  OAI22_X1 U4419 ( .A1(n12938), .A2(n13315), .B1(n7760), .B2(n12934), .ZN(
        n6254) );
  OAI22_X1 U4420 ( .A1(n12937), .A2(n13318), .B1(n7743), .B2(n12934), .ZN(
        n6255) );
  OAI22_X1 U4421 ( .A1(n12937), .A2(n13321), .B1(n7641), .B2(n12934), .ZN(
        n6256) );
  OAI22_X1 U4422 ( .A1(n12937), .A2(n13324), .B1(n7624), .B2(n12934), .ZN(
        n6257) );
  OAI22_X1 U4423 ( .A1(n12937), .A2(n13327), .B1(n7520), .B2(n12934), .ZN(
        n6258) );
  OAI22_X1 U4424 ( .A1(n12937), .A2(n13330), .B1(n7503), .B2(n12934), .ZN(
        n6259) );
  OAI22_X1 U4425 ( .A1(n12936), .A2(n13333), .B1(n7401), .B2(n12934), .ZN(
        n6260) );
  OAI22_X1 U4426 ( .A1(n12936), .A2(n13336), .B1(n7384), .B2(n12934), .ZN(
        n6261) );
  OAI22_X1 U4427 ( .A1(n12936), .A2(n13339), .B1(n7367), .B2(n12934), .ZN(
        n6262) );
  OAI22_X1 U4428 ( .A1(n12936), .A2(n13342), .B1(n7268), .B2(n12934), .ZN(
        n6263) );
  OAI22_X1 U4429 ( .A1(n12936), .A2(n13345), .B1(n7251), .B2(n12934), .ZN(
        n6264) );
  OAI22_X1 U4430 ( .A1(n12935), .A2(n13348), .B1(n7234), .B2(n12934), .ZN(
        n6265) );
  OAI22_X1 U4431 ( .A1(n13022), .A2(n13242), .B1(n8166), .B2(n13012), .ZN(
        n6486) );
  OAI22_X1 U4432 ( .A1(n13022), .A2(n13245), .B1(n8149), .B2(n13012), .ZN(
        n6487) );
  OAI22_X1 U4433 ( .A1(n13022), .A2(n13248), .B1(n8132), .B2(n13012), .ZN(
        n6488) );
  OAI22_X1 U4434 ( .A1(n13022), .A2(n13251), .B1(n8115), .B2(n13012), .ZN(
        n6489) );
  OAI22_X1 U4435 ( .A1(n13022), .A2(n13254), .B1(n8098), .B2(n13012), .ZN(
        n6490) );
  OAI22_X1 U4436 ( .A1(n13021), .A2(n13257), .B1(n8081), .B2(n13012), .ZN(
        n6491) );
  OAI22_X1 U4437 ( .A1(n13021), .A2(n13260), .B1(n8064), .B2(n13012), .ZN(
        n6492) );
  OAI22_X1 U4438 ( .A1(n13021), .A2(n13263), .B1(n8047), .B2(n13012), .ZN(
        n6493) );
  OAI22_X1 U4439 ( .A1(n13021), .A2(n13266), .B1(n8030), .B2(n13012), .ZN(
        n6494) );
  OAI22_X1 U4440 ( .A1(n13021), .A2(n13269), .B1(n8013), .B2(n13012), .ZN(
        n6495) );
  OAI22_X1 U4441 ( .A1(n13020), .A2(n13272), .B1(n7996), .B2(n13012), .ZN(
        n6496) );
  OAI22_X1 U4442 ( .A1(n13020), .A2(n13275), .B1(n7979), .B2(n13012), .ZN(
        n6497) );
  OAI22_X1 U4443 ( .A1(n13020), .A2(n13278), .B1(n7962), .B2(n13013), .ZN(
        n6498) );
  OAI22_X1 U4444 ( .A1(n13020), .A2(n13281), .B1(n7945), .B2(n13013), .ZN(
        n6499) );
  OAI22_X1 U4445 ( .A1(n13020), .A2(n13284), .B1(n7928), .B2(n13013), .ZN(
        n6500) );
  OAI22_X1 U4446 ( .A1(n13019), .A2(n13287), .B1(n7911), .B2(n13013), .ZN(
        n6501) );
  OAI22_X1 U4447 ( .A1(n13019), .A2(n13290), .B1(n7894), .B2(n13013), .ZN(
        n6502) );
  OAI22_X1 U4448 ( .A1(n13019), .A2(n13293), .B1(n7877), .B2(n13013), .ZN(
        n6503) );
  OAI22_X1 U4449 ( .A1(n13019), .A2(n13296), .B1(n7860), .B2(n13013), .ZN(
        n6504) );
  OAI22_X1 U4450 ( .A1(n13019), .A2(n13299), .B1(n7843), .B2(n13013), .ZN(
        n6505) );
  OAI22_X1 U4451 ( .A1(n13018), .A2(n13302), .B1(n7826), .B2(n13013), .ZN(
        n6506) );
  OAI22_X1 U4452 ( .A1(n13018), .A2(n13305), .B1(n7809), .B2(n13013), .ZN(
        n6507) );
  OAI22_X1 U4453 ( .A1(n13018), .A2(n13308), .B1(n7792), .B2(n13013), .ZN(
        n6508) );
  OAI22_X1 U4454 ( .A1(n13018), .A2(n13311), .B1(n7775), .B2(n13013), .ZN(
        n6509) );
  OAI22_X1 U4455 ( .A1(n13018), .A2(n13314), .B1(n7758), .B2(n13014), .ZN(
        n6510) );
  OAI22_X1 U4456 ( .A1(n13017), .A2(n13317), .B1(n7656), .B2(n13014), .ZN(
        n6511) );
  OAI22_X1 U4457 ( .A1(n13017), .A2(n13320), .B1(n7639), .B2(n13014), .ZN(
        n6512) );
  OAI22_X1 U4458 ( .A1(n13017), .A2(n13323), .B1(n7622), .B2(n13014), .ZN(
        n6513) );
  OAI22_X1 U4459 ( .A1(n13017), .A2(n13326), .B1(n7518), .B2(n13014), .ZN(
        n6514) );
  OAI22_X1 U4460 ( .A1(n13017), .A2(n13329), .B1(n7501), .B2(n13014), .ZN(
        n6515) );
  OAI22_X1 U4461 ( .A1(n13016), .A2(n13332), .B1(n7399), .B2(n13014), .ZN(
        n6516) );
  OAI22_X1 U4462 ( .A1(n13016), .A2(n13335), .B1(n7382), .B2(n13014), .ZN(
        n6517) );
  OAI22_X1 U4463 ( .A1(n13016), .A2(n13338), .B1(n7365), .B2(n13014), .ZN(
        n6518) );
  OAI22_X1 U4464 ( .A1(n13016), .A2(n13341), .B1(n7266), .B2(n13014), .ZN(
        n6519) );
  OAI22_X1 U4465 ( .A1(n13016), .A2(n13344), .B1(n7249), .B2(n13014), .ZN(
        n6520) );
  OAI22_X1 U4466 ( .A1(n13015), .A2(n13347), .B1(n7152), .B2(n13014), .ZN(
        n6521) );
  OAI22_X1 U4467 ( .A1(n13002), .A2(n13242), .B1(n8165), .B2(n12992), .ZN(
        n6422) );
  OAI22_X1 U4468 ( .A1(n13002), .A2(n13245), .B1(n8148), .B2(n12992), .ZN(
        n6423) );
  OAI22_X1 U4469 ( .A1(n13002), .A2(n13248), .B1(n8131), .B2(n12992), .ZN(
        n6424) );
  OAI22_X1 U4470 ( .A1(n13002), .A2(n13251), .B1(n8114), .B2(n12992), .ZN(
        n6425) );
  OAI22_X1 U4471 ( .A1(n13002), .A2(n13254), .B1(n8097), .B2(n12992), .ZN(
        n6426) );
  OAI22_X1 U4472 ( .A1(n13001), .A2(n13257), .B1(n8080), .B2(n12992), .ZN(
        n6427) );
  OAI22_X1 U4473 ( .A1(n13001), .A2(n13260), .B1(n8063), .B2(n12992), .ZN(
        n6428) );
  OAI22_X1 U4474 ( .A1(n13001), .A2(n13263), .B1(n8046), .B2(n12992), .ZN(
        n6429) );
  OAI22_X1 U4475 ( .A1(n13001), .A2(n13266), .B1(n8029), .B2(n12992), .ZN(
        n6430) );
  OAI22_X1 U4476 ( .A1(n13001), .A2(n13269), .B1(n8012), .B2(n12992), .ZN(
        n6431) );
  OAI22_X1 U4477 ( .A1(n13000), .A2(n13272), .B1(n7995), .B2(n12992), .ZN(
        n6432) );
  OAI22_X1 U4478 ( .A1(n13000), .A2(n13275), .B1(n7978), .B2(n12992), .ZN(
        n6433) );
  OAI22_X1 U4479 ( .A1(n13000), .A2(n13278), .B1(n7961), .B2(n12993), .ZN(
        n6434) );
  OAI22_X1 U4480 ( .A1(n13000), .A2(n13281), .B1(n7944), .B2(n12993), .ZN(
        n6435) );
  OAI22_X1 U4481 ( .A1(n13000), .A2(n13284), .B1(n7927), .B2(n12993), .ZN(
        n6436) );
  OAI22_X1 U4482 ( .A1(n12999), .A2(n13287), .B1(n7910), .B2(n12993), .ZN(
        n6437) );
  OAI22_X1 U4483 ( .A1(n12999), .A2(n13290), .B1(n7893), .B2(n12993), .ZN(
        n6438) );
  OAI22_X1 U4484 ( .A1(n12999), .A2(n13293), .B1(n7876), .B2(n12993), .ZN(
        n6439) );
  OAI22_X1 U4485 ( .A1(n12999), .A2(n13296), .B1(n7859), .B2(n12993), .ZN(
        n6440) );
  OAI22_X1 U4486 ( .A1(n12999), .A2(n13299), .B1(n7842), .B2(n12993), .ZN(
        n6441) );
  OAI22_X1 U4487 ( .A1(n12998), .A2(n13302), .B1(n7825), .B2(n12993), .ZN(
        n6442) );
  OAI22_X1 U4488 ( .A1(n12998), .A2(n13305), .B1(n7808), .B2(n12993), .ZN(
        n6443) );
  OAI22_X1 U4489 ( .A1(n12998), .A2(n13308), .B1(n7791), .B2(n12993), .ZN(
        n6444) );
  OAI22_X1 U4490 ( .A1(n12998), .A2(n13311), .B1(n7774), .B2(n12993), .ZN(
        n6445) );
  OAI22_X1 U4491 ( .A1(n12998), .A2(n13314), .B1(n7757), .B2(n12994), .ZN(
        n6446) );
  OAI22_X1 U4492 ( .A1(n12997), .A2(n13317), .B1(n7655), .B2(n12994), .ZN(
        n6447) );
  OAI22_X1 U4493 ( .A1(n12997), .A2(n13320), .B1(n7638), .B2(n12994), .ZN(
        n6448) );
  OAI22_X1 U4494 ( .A1(n12997), .A2(n13323), .B1(n7621), .B2(n12994), .ZN(
        n6449) );
  OAI22_X1 U4495 ( .A1(n12997), .A2(n13326), .B1(n7517), .B2(n12994), .ZN(
        n6450) );
  OAI22_X1 U4496 ( .A1(n12997), .A2(n13329), .B1(n7500), .B2(n12994), .ZN(
        n6451) );
  OAI22_X1 U4497 ( .A1(n12996), .A2(n13332), .B1(n7398), .B2(n12994), .ZN(
        n6452) );
  OAI22_X1 U4498 ( .A1(n12996), .A2(n13335), .B1(n7381), .B2(n12994), .ZN(
        n6453) );
  OAI22_X1 U4499 ( .A1(n12996), .A2(n13338), .B1(n7364), .B2(n12994), .ZN(
        n6454) );
  OAI22_X1 U4500 ( .A1(n12996), .A2(n13341), .B1(n7265), .B2(n12994), .ZN(
        n6455) );
  OAI22_X1 U4501 ( .A1(n12996), .A2(n13344), .B1(n7248), .B2(n12994), .ZN(
        n6456) );
  OAI22_X1 U4502 ( .A1(n12995), .A2(n13347), .B1(n7151), .B2(n12994), .ZN(
        n6457) );
  OAI22_X1 U4503 ( .A1(n13062), .A2(n13242), .B1(n8163), .B2(n13052), .ZN(
        n6614) );
  OAI22_X1 U4504 ( .A1(n13062), .A2(n13245), .B1(n8146), .B2(n13052), .ZN(
        n6615) );
  OAI22_X1 U4505 ( .A1(n13062), .A2(n13248), .B1(n8129), .B2(n13052), .ZN(
        n6616) );
  OAI22_X1 U4506 ( .A1(n13062), .A2(n13251), .B1(n8112), .B2(n13052), .ZN(
        n6617) );
  OAI22_X1 U4507 ( .A1(n13062), .A2(n13254), .B1(n8095), .B2(n13052), .ZN(
        n6618) );
  OAI22_X1 U4508 ( .A1(n13061), .A2(n13257), .B1(n8078), .B2(n13052), .ZN(
        n6619) );
  OAI22_X1 U4509 ( .A1(n13061), .A2(n13260), .B1(n8061), .B2(n13052), .ZN(
        n6620) );
  OAI22_X1 U4510 ( .A1(n13061), .A2(n13263), .B1(n8044), .B2(n13052), .ZN(
        n6621) );
  OAI22_X1 U4511 ( .A1(n13061), .A2(n13266), .B1(n8027), .B2(n13052), .ZN(
        n6622) );
  OAI22_X1 U4512 ( .A1(n13061), .A2(n13269), .B1(n8010), .B2(n13052), .ZN(
        n6623) );
  OAI22_X1 U4513 ( .A1(n13060), .A2(n13272), .B1(n7993), .B2(n13052), .ZN(
        n6624) );
  OAI22_X1 U4514 ( .A1(n13060), .A2(n13275), .B1(n7976), .B2(n13052), .ZN(
        n6625) );
  OAI22_X1 U4515 ( .A1(n13060), .A2(n13278), .B1(n7959), .B2(n13053), .ZN(
        n6626) );
  OAI22_X1 U4516 ( .A1(n13060), .A2(n13281), .B1(n7942), .B2(n13053), .ZN(
        n6627) );
  OAI22_X1 U4517 ( .A1(n13060), .A2(n13284), .B1(n7925), .B2(n13053), .ZN(
        n6628) );
  OAI22_X1 U4518 ( .A1(n13059), .A2(n13287), .B1(n7908), .B2(n13053), .ZN(
        n6629) );
  OAI22_X1 U4519 ( .A1(n13059), .A2(n13290), .B1(n7891), .B2(n13053), .ZN(
        n6630) );
  OAI22_X1 U4520 ( .A1(n13059), .A2(n13293), .B1(n7874), .B2(n13053), .ZN(
        n6631) );
  OAI22_X1 U4521 ( .A1(n13059), .A2(n13296), .B1(n7857), .B2(n13053), .ZN(
        n6632) );
  OAI22_X1 U4522 ( .A1(n13059), .A2(n13299), .B1(n7840), .B2(n13053), .ZN(
        n6633) );
  OAI22_X1 U4523 ( .A1(n13058), .A2(n13302), .B1(n7823), .B2(n13053), .ZN(
        n6634) );
  OAI22_X1 U4524 ( .A1(n13058), .A2(n13305), .B1(n7806), .B2(n13053), .ZN(
        n6635) );
  OAI22_X1 U4525 ( .A1(n13058), .A2(n13308), .B1(n7789), .B2(n13053), .ZN(
        n6636) );
  OAI22_X1 U4526 ( .A1(n13058), .A2(n13311), .B1(n7772), .B2(n13053), .ZN(
        n6637) );
  OAI22_X1 U4527 ( .A1(n13058), .A2(n13314), .B1(n7755), .B2(n13054), .ZN(
        n6638) );
  OAI22_X1 U4528 ( .A1(n13057), .A2(n13317), .B1(n7653), .B2(n13054), .ZN(
        n6639) );
  OAI22_X1 U4529 ( .A1(n13057), .A2(n13320), .B1(n7636), .B2(n13054), .ZN(
        n6640) );
  OAI22_X1 U4530 ( .A1(n13057), .A2(n13323), .B1(n7619), .B2(n13054), .ZN(
        n6641) );
  OAI22_X1 U4531 ( .A1(n13057), .A2(n13326), .B1(n7515), .B2(n13054), .ZN(
        n6642) );
  OAI22_X1 U4532 ( .A1(n13057), .A2(n13329), .B1(n7498), .B2(n13054), .ZN(
        n6643) );
  OAI22_X1 U4533 ( .A1(n13056), .A2(n13332), .B1(n7396), .B2(n13054), .ZN(
        n6644) );
  OAI22_X1 U4534 ( .A1(n13056), .A2(n13335), .B1(n7379), .B2(n13054), .ZN(
        n6645) );
  OAI22_X1 U4535 ( .A1(n13056), .A2(n13338), .B1(n7362), .B2(n13054), .ZN(
        n6646) );
  OAI22_X1 U4536 ( .A1(n13056), .A2(n13341), .B1(n7263), .B2(n13054), .ZN(
        n6647) );
  OAI22_X1 U4537 ( .A1(n13056), .A2(n13344), .B1(n7246), .B2(n13054), .ZN(
        n6648) );
  OAI22_X1 U4538 ( .A1(n13055), .A2(n13347), .B1(n7149), .B2(n13054), .ZN(
        n6649) );
  OAI22_X1 U4539 ( .A1(n13042), .A2(n13242), .B1(n8164), .B2(n13032), .ZN(
        n6550) );
  OAI22_X1 U4540 ( .A1(n13042), .A2(n13245), .B1(n8147), .B2(n13032), .ZN(
        n6551) );
  OAI22_X1 U4541 ( .A1(n13042), .A2(n13248), .B1(n8130), .B2(n13032), .ZN(
        n6552) );
  OAI22_X1 U4542 ( .A1(n13042), .A2(n13251), .B1(n8113), .B2(n13032), .ZN(
        n6553) );
  OAI22_X1 U4543 ( .A1(n13042), .A2(n13254), .B1(n8096), .B2(n13032), .ZN(
        n6554) );
  OAI22_X1 U4544 ( .A1(n13041), .A2(n13257), .B1(n8079), .B2(n13032), .ZN(
        n6555) );
  OAI22_X1 U4545 ( .A1(n13041), .A2(n13260), .B1(n8062), .B2(n13032), .ZN(
        n6556) );
  OAI22_X1 U4546 ( .A1(n13041), .A2(n13263), .B1(n8045), .B2(n13032), .ZN(
        n6557) );
  OAI22_X1 U4547 ( .A1(n13041), .A2(n13266), .B1(n8028), .B2(n13032), .ZN(
        n6558) );
  OAI22_X1 U4548 ( .A1(n13041), .A2(n13269), .B1(n8011), .B2(n13032), .ZN(
        n6559) );
  OAI22_X1 U4549 ( .A1(n13040), .A2(n13272), .B1(n7994), .B2(n13032), .ZN(
        n6560) );
  OAI22_X1 U4550 ( .A1(n13040), .A2(n13275), .B1(n7977), .B2(n13032), .ZN(
        n6561) );
  OAI22_X1 U4551 ( .A1(n13040), .A2(n13278), .B1(n7960), .B2(n13033), .ZN(
        n6562) );
  OAI22_X1 U4552 ( .A1(n13040), .A2(n13281), .B1(n7943), .B2(n13033), .ZN(
        n6563) );
  OAI22_X1 U4553 ( .A1(n13040), .A2(n13284), .B1(n7926), .B2(n13033), .ZN(
        n6564) );
  OAI22_X1 U4554 ( .A1(n13039), .A2(n13287), .B1(n7909), .B2(n13033), .ZN(
        n6565) );
  OAI22_X1 U4555 ( .A1(n13039), .A2(n13290), .B1(n7892), .B2(n13033), .ZN(
        n6566) );
  OAI22_X1 U4556 ( .A1(n13039), .A2(n13293), .B1(n7875), .B2(n13033), .ZN(
        n6567) );
  OAI22_X1 U4557 ( .A1(n13039), .A2(n13296), .B1(n7858), .B2(n13033), .ZN(
        n6568) );
  OAI22_X1 U4558 ( .A1(n13039), .A2(n13299), .B1(n7841), .B2(n13033), .ZN(
        n6569) );
  OAI22_X1 U4559 ( .A1(n13038), .A2(n13302), .B1(n7824), .B2(n13033), .ZN(
        n6570) );
  OAI22_X1 U4560 ( .A1(n13038), .A2(n13305), .B1(n7807), .B2(n13033), .ZN(
        n6571) );
  OAI22_X1 U4561 ( .A1(n13038), .A2(n13308), .B1(n7790), .B2(n13033), .ZN(
        n6572) );
  OAI22_X1 U4562 ( .A1(n13038), .A2(n13311), .B1(n7773), .B2(n13033), .ZN(
        n6573) );
  OAI22_X1 U4563 ( .A1(n13038), .A2(n13314), .B1(n7756), .B2(n13034), .ZN(
        n6574) );
  OAI22_X1 U4564 ( .A1(n13037), .A2(n13317), .B1(n7654), .B2(n13034), .ZN(
        n6575) );
  OAI22_X1 U4565 ( .A1(n13037), .A2(n13320), .B1(n7637), .B2(n13034), .ZN(
        n6576) );
  OAI22_X1 U4566 ( .A1(n13037), .A2(n13323), .B1(n7620), .B2(n13034), .ZN(
        n6577) );
  OAI22_X1 U4567 ( .A1(n13037), .A2(n13326), .B1(n7516), .B2(n13034), .ZN(
        n6578) );
  OAI22_X1 U4568 ( .A1(n13037), .A2(n13329), .B1(n7499), .B2(n13034), .ZN(
        n6579) );
  OAI22_X1 U4569 ( .A1(n13036), .A2(n13332), .B1(n7397), .B2(n13034), .ZN(
        n6580) );
  OAI22_X1 U4570 ( .A1(n13036), .A2(n13335), .B1(n7380), .B2(n13034), .ZN(
        n6581) );
  OAI22_X1 U4571 ( .A1(n13036), .A2(n13338), .B1(n7363), .B2(n13034), .ZN(
        n6582) );
  OAI22_X1 U4572 ( .A1(n13036), .A2(n13341), .B1(n7264), .B2(n13034), .ZN(
        n6583) );
  OAI22_X1 U4573 ( .A1(n13036), .A2(n13344), .B1(n7247), .B2(n13034), .ZN(
        n6584) );
  OAI22_X1 U4574 ( .A1(n13035), .A2(n13347), .B1(n7150), .B2(n13034), .ZN(
        n6585) );
  OAI22_X1 U4575 ( .A1(n12865), .A2(n13207), .B1(n8374), .B2(n12851), .ZN(
        n5962) );
  OAI22_X1 U4576 ( .A1(n12865), .A2(n13210), .B1(n8357), .B2(n12851), .ZN(
        n5963) );
  OAI22_X1 U4577 ( .A1(n12864), .A2(n13213), .B1(n8340), .B2(n12851), .ZN(
        n5964) );
  OAI22_X1 U4578 ( .A1(n12864), .A2(n13216), .B1(n8323), .B2(n12851), .ZN(
        n5965) );
  OAI22_X1 U4579 ( .A1(n12864), .A2(n13219), .B1(n8306), .B2(n12851), .ZN(
        n5966) );
  OAI22_X1 U4580 ( .A1(n12864), .A2(n13222), .B1(n8289), .B2(n12851), .ZN(
        n5967) );
  OAI22_X1 U4581 ( .A1(n12864), .A2(n13225), .B1(n8272), .B2(n12851), .ZN(
        n5968) );
  OAI22_X1 U4582 ( .A1(n12863), .A2(n13228), .B1(n8255), .B2(n12851), .ZN(
        n5969) );
  OAI22_X1 U4583 ( .A1(n12863), .A2(n13231), .B1(n8238), .B2(n12851), .ZN(
        n5970) );
  OAI22_X1 U4584 ( .A1(n12863), .A2(n13234), .B1(n8221), .B2(n12851), .ZN(
        n5971) );
  OAI22_X1 U4585 ( .A1(n12863), .A2(n13237), .B1(n8204), .B2(n12851), .ZN(
        n5972) );
  OAI22_X1 U4586 ( .A1(n12863), .A2(n13240), .B1(n8187), .B2(n12851), .ZN(
        n5973) );
  OAI22_X1 U4587 ( .A1(n12862), .A2(n13243), .B1(n8170), .B2(n12852), .ZN(
        n5974) );
  OAI22_X1 U4588 ( .A1(n12862), .A2(n13246), .B1(n8153), .B2(n12852), .ZN(
        n5975) );
  OAI22_X1 U4589 ( .A1(n12862), .A2(n13249), .B1(n8136), .B2(n12852), .ZN(
        n5976) );
  OAI22_X1 U4590 ( .A1(n12862), .A2(n13252), .B1(n8119), .B2(n12852), .ZN(
        n5977) );
  OAI22_X1 U4591 ( .A1(n12862), .A2(n13255), .B1(n8102), .B2(n12852), .ZN(
        n5978) );
  OAI22_X1 U4592 ( .A1(n12861), .A2(n13258), .B1(n8085), .B2(n12852), .ZN(
        n5979) );
  OAI22_X1 U4593 ( .A1(n12861), .A2(n13261), .B1(n8068), .B2(n12852), .ZN(
        n5980) );
  OAI22_X1 U4594 ( .A1(n12861), .A2(n13264), .B1(n8051), .B2(n12852), .ZN(
        n5981) );
  OAI22_X1 U4595 ( .A1(n12861), .A2(n13267), .B1(n8034), .B2(n12852), .ZN(
        n5982) );
  OAI22_X1 U4596 ( .A1(n12861), .A2(n13270), .B1(n8017), .B2(n12852), .ZN(
        n5983) );
  OAI22_X1 U4597 ( .A1(n12860), .A2(n13273), .B1(n8000), .B2(n12852), .ZN(
        n5984) );
  OAI22_X1 U4598 ( .A1(n12860), .A2(n13276), .B1(n7983), .B2(n12852), .ZN(
        n5985) );
  OAI22_X1 U4599 ( .A1(n12860), .A2(n13279), .B1(n7966), .B2(n12853), .ZN(
        n5986) );
  OAI22_X1 U4600 ( .A1(n12860), .A2(n13282), .B1(n7949), .B2(n12853), .ZN(
        n5987) );
  OAI22_X1 U4601 ( .A1(n12860), .A2(n13285), .B1(n7932), .B2(n12853), .ZN(
        n5988) );
  OAI22_X1 U4602 ( .A1(n12859), .A2(n13288), .B1(n7915), .B2(n12853), .ZN(
        n5989) );
  OAI22_X1 U4603 ( .A1(n12859), .A2(n13291), .B1(n7898), .B2(n12853), .ZN(
        n5990) );
  OAI22_X1 U4604 ( .A1(n12859), .A2(n13294), .B1(n7881), .B2(n12853), .ZN(
        n5991) );
  OAI22_X1 U4605 ( .A1(n12859), .A2(n13297), .B1(n7864), .B2(n12853), .ZN(
        n5992) );
  OAI22_X1 U4606 ( .A1(n12859), .A2(n13300), .B1(n7847), .B2(n12853), .ZN(
        n5993) );
  OAI22_X1 U4607 ( .A1(n12858), .A2(n13303), .B1(n7830), .B2(n12853), .ZN(
        n5994) );
  OAI22_X1 U4608 ( .A1(n12858), .A2(n13306), .B1(n7813), .B2(n12853), .ZN(
        n5995) );
  OAI22_X1 U4609 ( .A1(n12858), .A2(n13309), .B1(n7796), .B2(n12853), .ZN(
        n5996) );
  OAI22_X1 U4610 ( .A1(n12858), .A2(n13312), .B1(n7779), .B2(n12853), .ZN(
        n5997) );
  OAI22_X1 U4611 ( .A1(n12858), .A2(n13315), .B1(n7762), .B2(n12854), .ZN(
        n5998) );
  OAI22_X1 U4612 ( .A1(n12857), .A2(n13318), .B1(n7745), .B2(n12854), .ZN(
        n5999) );
  OAI22_X1 U4613 ( .A1(n12857), .A2(n13321), .B1(n7643), .B2(n12854), .ZN(
        n6000) );
  OAI22_X1 U4614 ( .A1(n12857), .A2(n13324), .B1(n7626), .B2(n12854), .ZN(
        n6001) );
  OAI22_X1 U4615 ( .A1(n12857), .A2(n13327), .B1(n7522), .B2(n12854), .ZN(
        n6002) );
  OAI22_X1 U4616 ( .A1(n12857), .A2(n13330), .B1(n7505), .B2(n12854), .ZN(
        n6003) );
  OAI22_X1 U4617 ( .A1(n12856), .A2(n13333), .B1(n7403), .B2(n12854), .ZN(
        n6004) );
  OAI22_X1 U4618 ( .A1(n12856), .A2(n13336), .B1(n7386), .B2(n12854), .ZN(
        n6005) );
  OAI22_X1 U4619 ( .A1(n12856), .A2(n13339), .B1(n7369), .B2(n12854), .ZN(
        n6006) );
  OAI22_X1 U4620 ( .A1(n12856), .A2(n13342), .B1(n7270), .B2(n12854), .ZN(
        n6007) );
  OAI22_X1 U4621 ( .A1(n12856), .A2(n13345), .B1(n7253), .B2(n12854), .ZN(
        n6008) );
  OAI22_X1 U4622 ( .A1(n12855), .A2(n13348), .B1(n7236), .B2(n12854), .ZN(
        n6009) );
  OAI22_X1 U4623 ( .A1(n12842), .A2(n13243), .B1(n8169), .B2(n12832), .ZN(
        n5910) );
  OAI22_X1 U4624 ( .A1(n12842), .A2(n13246), .B1(n8152), .B2(n12832), .ZN(
        n5911) );
  OAI22_X1 U4625 ( .A1(n12842), .A2(n13249), .B1(n8135), .B2(n12832), .ZN(
        n5912) );
  OAI22_X1 U4626 ( .A1(n12842), .A2(n13252), .B1(n8118), .B2(n12832), .ZN(
        n5913) );
  OAI22_X1 U4627 ( .A1(n12842), .A2(n13255), .B1(n8101), .B2(n12832), .ZN(
        n5914) );
  OAI22_X1 U4628 ( .A1(n12841), .A2(n13258), .B1(n8084), .B2(n12832), .ZN(
        n5915) );
  OAI22_X1 U4629 ( .A1(n12841), .A2(n13261), .B1(n8067), .B2(n12832), .ZN(
        n5916) );
  OAI22_X1 U4630 ( .A1(n12841), .A2(n13264), .B1(n8050), .B2(n12832), .ZN(
        n5917) );
  OAI22_X1 U4631 ( .A1(n12841), .A2(n13267), .B1(n8033), .B2(n12832), .ZN(
        n5918) );
  OAI22_X1 U4632 ( .A1(n12841), .A2(n13270), .B1(n8016), .B2(n12832), .ZN(
        n5919) );
  OAI22_X1 U4633 ( .A1(n12840), .A2(n13273), .B1(n7999), .B2(n12832), .ZN(
        n5920) );
  OAI22_X1 U4634 ( .A1(n12840), .A2(n13276), .B1(n7982), .B2(n12832), .ZN(
        n5921) );
  OAI22_X1 U4635 ( .A1(n12840), .A2(n13279), .B1(n7965), .B2(n12833), .ZN(
        n5922) );
  OAI22_X1 U4636 ( .A1(n12840), .A2(n13282), .B1(n7948), .B2(n12833), .ZN(
        n5923) );
  OAI22_X1 U4637 ( .A1(n12840), .A2(n13285), .B1(n7931), .B2(n12833), .ZN(
        n5924) );
  OAI22_X1 U4638 ( .A1(n12839), .A2(n13288), .B1(n7914), .B2(n12833), .ZN(
        n5925) );
  OAI22_X1 U4639 ( .A1(n12839), .A2(n13291), .B1(n7897), .B2(n12833), .ZN(
        n5926) );
  OAI22_X1 U4640 ( .A1(n12839), .A2(n13294), .B1(n7880), .B2(n12833), .ZN(
        n5927) );
  OAI22_X1 U4641 ( .A1(n12839), .A2(n13297), .B1(n7863), .B2(n12833), .ZN(
        n5928) );
  OAI22_X1 U4642 ( .A1(n12839), .A2(n13300), .B1(n7846), .B2(n12833), .ZN(
        n5929) );
  OAI22_X1 U4643 ( .A1(n12838), .A2(n13303), .B1(n7829), .B2(n12833), .ZN(
        n5930) );
  OAI22_X1 U4644 ( .A1(n12838), .A2(n13306), .B1(n7812), .B2(n12833), .ZN(
        n5931) );
  OAI22_X1 U4645 ( .A1(n12838), .A2(n13309), .B1(n7795), .B2(n12833), .ZN(
        n5932) );
  OAI22_X1 U4646 ( .A1(n12838), .A2(n13312), .B1(n7778), .B2(n12833), .ZN(
        n5933) );
  OAI22_X1 U4647 ( .A1(n12838), .A2(n13315), .B1(n7761), .B2(n12834), .ZN(
        n5934) );
  OAI22_X1 U4648 ( .A1(n12837), .A2(n13318), .B1(n7744), .B2(n12834), .ZN(
        n5935) );
  OAI22_X1 U4649 ( .A1(n12837), .A2(n13321), .B1(n7642), .B2(n12834), .ZN(
        n5936) );
  OAI22_X1 U4650 ( .A1(n12837), .A2(n13324), .B1(n7625), .B2(n12834), .ZN(
        n5937) );
  OAI22_X1 U4651 ( .A1(n12837), .A2(n13327), .B1(n7521), .B2(n12834), .ZN(
        n5938) );
  OAI22_X1 U4652 ( .A1(n12837), .A2(n13330), .B1(n7504), .B2(n12834), .ZN(
        n5939) );
  OAI22_X1 U4653 ( .A1(n12836), .A2(n13333), .B1(n7402), .B2(n12834), .ZN(
        n5940) );
  OAI22_X1 U4654 ( .A1(n12836), .A2(n13336), .B1(n7385), .B2(n12834), .ZN(
        n5941) );
  OAI22_X1 U4655 ( .A1(n12836), .A2(n13339), .B1(n7368), .B2(n12834), .ZN(
        n5942) );
  OAI22_X1 U4656 ( .A1(n12836), .A2(n13342), .B1(n7269), .B2(n12834), .ZN(
        n5943) );
  OAI22_X1 U4657 ( .A1(n12836), .A2(n13345), .B1(n7252), .B2(n12834), .ZN(
        n5944) );
  OAI22_X1 U4658 ( .A1(n12835), .A2(n13348), .B1(n7235), .B2(n12834), .ZN(
        n5945) );
  OAI22_X1 U4659 ( .A1(n12782), .A2(n13243), .B1(n8172), .B2(n12772), .ZN(
        n5718) );
  OAI22_X1 U4660 ( .A1(n12782), .A2(n13246), .B1(n8155), .B2(n12772), .ZN(
        n5719) );
  OAI22_X1 U4661 ( .A1(n12782), .A2(n13249), .B1(n8138), .B2(n12772), .ZN(
        n5720) );
  OAI22_X1 U4662 ( .A1(n12782), .A2(n13252), .B1(n8121), .B2(n12772), .ZN(
        n5721) );
  OAI22_X1 U4663 ( .A1(n12782), .A2(n13255), .B1(n8104), .B2(n12772), .ZN(
        n5722) );
  OAI22_X1 U4664 ( .A1(n12781), .A2(n13258), .B1(n8087), .B2(n12772), .ZN(
        n5723) );
  OAI22_X1 U4665 ( .A1(n12781), .A2(n13261), .B1(n8070), .B2(n12772), .ZN(
        n5724) );
  OAI22_X1 U4666 ( .A1(n12781), .A2(n13264), .B1(n8053), .B2(n12772), .ZN(
        n5725) );
  OAI22_X1 U4667 ( .A1(n12781), .A2(n13267), .B1(n8036), .B2(n12772), .ZN(
        n5726) );
  OAI22_X1 U4668 ( .A1(n12781), .A2(n13270), .B1(n8019), .B2(n12772), .ZN(
        n5727) );
  OAI22_X1 U4669 ( .A1(n12780), .A2(n13273), .B1(n8002), .B2(n12772), .ZN(
        n5728) );
  OAI22_X1 U4670 ( .A1(n12780), .A2(n13276), .B1(n7985), .B2(n12772), .ZN(
        n5729) );
  OAI22_X1 U4671 ( .A1(n12780), .A2(n13279), .B1(n7968), .B2(n12773), .ZN(
        n5730) );
  OAI22_X1 U4672 ( .A1(n12780), .A2(n13282), .B1(n7951), .B2(n12773), .ZN(
        n5731) );
  OAI22_X1 U4673 ( .A1(n12780), .A2(n13285), .B1(n7934), .B2(n12773), .ZN(
        n5732) );
  OAI22_X1 U4674 ( .A1(n12779), .A2(n13288), .B1(n7917), .B2(n12773), .ZN(
        n5733) );
  OAI22_X1 U4675 ( .A1(n12779), .A2(n13291), .B1(n7900), .B2(n12773), .ZN(
        n5734) );
  OAI22_X1 U4676 ( .A1(n12779), .A2(n13294), .B1(n7883), .B2(n12773), .ZN(
        n5735) );
  OAI22_X1 U4677 ( .A1(n12779), .A2(n13297), .B1(n7866), .B2(n12773), .ZN(
        n5736) );
  OAI22_X1 U4678 ( .A1(n12779), .A2(n13300), .B1(n7849), .B2(n12773), .ZN(
        n5737) );
  OAI22_X1 U4679 ( .A1(n12778), .A2(n13303), .B1(n7832), .B2(n12773), .ZN(
        n5738) );
  OAI22_X1 U4680 ( .A1(n12778), .A2(n13306), .B1(n7815), .B2(n12773), .ZN(
        n5739) );
  OAI22_X1 U4681 ( .A1(n12778), .A2(n13309), .B1(n7798), .B2(n12773), .ZN(
        n5740) );
  OAI22_X1 U4682 ( .A1(n12778), .A2(n13312), .B1(n7781), .B2(n12773), .ZN(
        n5741) );
  OAI22_X1 U4683 ( .A1(n12778), .A2(n13315), .B1(n7764), .B2(n12774), .ZN(
        n5742) );
  OAI22_X1 U4684 ( .A1(n12777), .A2(n13318), .B1(n7747), .B2(n12774), .ZN(
        n5743) );
  OAI22_X1 U4685 ( .A1(n12777), .A2(n13321), .B1(n7645), .B2(n12774), .ZN(
        n5744) );
  OAI22_X1 U4686 ( .A1(n12777), .A2(n13324), .B1(n7628), .B2(n12774), .ZN(
        n5745) );
  OAI22_X1 U4687 ( .A1(n12777), .A2(n13327), .B1(n7524), .B2(n12774), .ZN(
        n5746) );
  OAI22_X1 U4688 ( .A1(n12777), .A2(n13330), .B1(n7507), .B2(n12774), .ZN(
        n5747) );
  OAI22_X1 U4689 ( .A1(n12776), .A2(n13333), .B1(n7490), .B2(n12774), .ZN(
        n5748) );
  OAI22_X1 U4690 ( .A1(n12776), .A2(n13336), .B1(n7388), .B2(n12774), .ZN(
        n5749) );
  OAI22_X1 U4691 ( .A1(n12776), .A2(n13339), .B1(n7371), .B2(n12774), .ZN(
        n5750) );
  OAI22_X1 U4692 ( .A1(n12776), .A2(n13342), .B1(n7272), .B2(n12774), .ZN(
        n5751) );
  OAI22_X1 U4693 ( .A1(n12776), .A2(n13345), .B1(n7255), .B2(n12774), .ZN(
        n5752) );
  OAI22_X1 U4694 ( .A1(n12775), .A2(n13348), .B1(n7238), .B2(n12774), .ZN(
        n5753) );
  OAI22_X1 U4695 ( .A1(n12762), .A2(n13243), .B1(n8171), .B2(n12752), .ZN(
        n5654) );
  OAI22_X1 U4696 ( .A1(n12762), .A2(n13246), .B1(n8154), .B2(n12752), .ZN(
        n5655) );
  OAI22_X1 U4697 ( .A1(n12762), .A2(n13249), .B1(n8137), .B2(n12752), .ZN(
        n5656) );
  OAI22_X1 U4698 ( .A1(n12762), .A2(n13252), .B1(n8120), .B2(n12752), .ZN(
        n5657) );
  OAI22_X1 U4699 ( .A1(n12762), .A2(n13255), .B1(n8103), .B2(n12752), .ZN(
        n5658) );
  OAI22_X1 U4700 ( .A1(n12761), .A2(n13258), .B1(n8086), .B2(n12752), .ZN(
        n5659) );
  OAI22_X1 U4701 ( .A1(n12761), .A2(n13261), .B1(n8069), .B2(n12752), .ZN(
        n5660) );
  OAI22_X1 U4702 ( .A1(n12761), .A2(n13264), .B1(n8052), .B2(n12752), .ZN(
        n5661) );
  OAI22_X1 U4703 ( .A1(n12761), .A2(n13267), .B1(n8035), .B2(n12752), .ZN(
        n5662) );
  OAI22_X1 U4704 ( .A1(n12761), .A2(n13270), .B1(n8018), .B2(n12752), .ZN(
        n5663) );
  OAI22_X1 U4705 ( .A1(n12760), .A2(n13273), .B1(n8001), .B2(n12752), .ZN(
        n5664) );
  OAI22_X1 U4706 ( .A1(n12760), .A2(n13276), .B1(n7984), .B2(n12752), .ZN(
        n5665) );
  OAI22_X1 U4707 ( .A1(n12760), .A2(n13279), .B1(n7967), .B2(n12753), .ZN(
        n5666) );
  OAI22_X1 U4708 ( .A1(n12760), .A2(n13282), .B1(n7950), .B2(n12753), .ZN(
        n5667) );
  OAI22_X1 U4709 ( .A1(n12760), .A2(n13285), .B1(n7933), .B2(n12753), .ZN(
        n5668) );
  OAI22_X1 U4710 ( .A1(n12759), .A2(n13288), .B1(n7916), .B2(n12753), .ZN(
        n5669) );
  OAI22_X1 U4711 ( .A1(n12759), .A2(n13291), .B1(n7899), .B2(n12753), .ZN(
        n5670) );
  OAI22_X1 U4712 ( .A1(n12759), .A2(n13294), .B1(n7882), .B2(n12753), .ZN(
        n5671) );
  OAI22_X1 U4713 ( .A1(n12759), .A2(n13297), .B1(n7865), .B2(n12753), .ZN(
        n5672) );
  OAI22_X1 U4714 ( .A1(n12759), .A2(n13300), .B1(n7848), .B2(n12753), .ZN(
        n5673) );
  OAI22_X1 U4715 ( .A1(n12758), .A2(n13303), .B1(n7831), .B2(n12753), .ZN(
        n5674) );
  OAI22_X1 U4716 ( .A1(n12758), .A2(n13306), .B1(n7814), .B2(n12753), .ZN(
        n5675) );
  OAI22_X1 U4717 ( .A1(n12758), .A2(n13309), .B1(n7797), .B2(n12753), .ZN(
        n5676) );
  OAI22_X1 U4718 ( .A1(n12758), .A2(n13312), .B1(n7780), .B2(n12753), .ZN(
        n5677) );
  OAI22_X1 U4719 ( .A1(n12758), .A2(n13315), .B1(n7763), .B2(n12754), .ZN(
        n5678) );
  OAI22_X1 U4720 ( .A1(n12757), .A2(n13318), .B1(n7746), .B2(n12754), .ZN(
        n5679) );
  OAI22_X1 U4721 ( .A1(n12757), .A2(n13321), .B1(n7644), .B2(n12754), .ZN(
        n5680) );
  OAI22_X1 U4722 ( .A1(n12757), .A2(n13324), .B1(n7627), .B2(n12754), .ZN(
        n5681) );
  OAI22_X1 U4723 ( .A1(n12757), .A2(n13327), .B1(n7523), .B2(n12754), .ZN(
        n5682) );
  OAI22_X1 U4724 ( .A1(n12757), .A2(n13330), .B1(n7506), .B2(n12754), .ZN(
        n5683) );
  OAI22_X1 U4725 ( .A1(n12756), .A2(n13333), .B1(n7404), .B2(n12754), .ZN(
        n5684) );
  OAI22_X1 U4726 ( .A1(n12756), .A2(n13336), .B1(n7387), .B2(n12754), .ZN(
        n5685) );
  OAI22_X1 U4727 ( .A1(n12756), .A2(n13339), .B1(n7370), .B2(n12754), .ZN(
        n5686) );
  OAI22_X1 U4728 ( .A1(n12756), .A2(n13342), .B1(n7271), .B2(n12754), .ZN(
        n5687) );
  OAI22_X1 U4729 ( .A1(n12756), .A2(n13345), .B1(n7254), .B2(n12754), .ZN(
        n5688) );
  OAI22_X1 U4730 ( .A1(n12755), .A2(n13348), .B1(n7237), .B2(n12754), .ZN(
        n5689) );
  OAI22_X1 U4731 ( .A1(n12588), .A2(n13244), .B1(n8176), .B2(n12578), .ZN(
        n5078) );
  OAI22_X1 U4732 ( .A1(n12588), .A2(n13247), .B1(n8159), .B2(n12578), .ZN(
        n5079) );
  OAI22_X1 U4733 ( .A1(n12588), .A2(n13250), .B1(n8142), .B2(n12578), .ZN(
        n5080) );
  OAI22_X1 U4734 ( .A1(n12588), .A2(n13253), .B1(n8125), .B2(n12578), .ZN(
        n5081) );
  OAI22_X1 U4735 ( .A1(n12588), .A2(n13256), .B1(n8108), .B2(n12578), .ZN(
        n5082) );
  OAI22_X1 U4736 ( .A1(n12587), .A2(n13259), .B1(n8091), .B2(n12578), .ZN(
        n5083) );
  OAI22_X1 U4737 ( .A1(n12587), .A2(n13262), .B1(n8074), .B2(n12578), .ZN(
        n5084) );
  OAI22_X1 U4738 ( .A1(n12587), .A2(n13265), .B1(n8057), .B2(n12578), .ZN(
        n5085) );
  OAI22_X1 U4739 ( .A1(n12587), .A2(n13268), .B1(n8040), .B2(n12578), .ZN(
        n5086) );
  OAI22_X1 U4740 ( .A1(n12587), .A2(n13271), .B1(n8023), .B2(n12578), .ZN(
        n5087) );
  OAI22_X1 U4741 ( .A1(n12586), .A2(n13274), .B1(n8006), .B2(n12578), .ZN(
        n5088) );
  OAI22_X1 U4742 ( .A1(n12586), .A2(n13277), .B1(n7989), .B2(n12578), .ZN(
        n5089) );
  OAI22_X1 U4743 ( .A1(n12586), .A2(n13280), .B1(n7972), .B2(n12579), .ZN(
        n5090) );
  OAI22_X1 U4744 ( .A1(n12586), .A2(n13283), .B1(n7955), .B2(n12579), .ZN(
        n5091) );
  OAI22_X1 U4745 ( .A1(n12586), .A2(n13286), .B1(n7938), .B2(n12579), .ZN(
        n5092) );
  OAI22_X1 U4746 ( .A1(n12585), .A2(n13289), .B1(n7921), .B2(n12579), .ZN(
        n5093) );
  OAI22_X1 U4747 ( .A1(n12585), .A2(n13292), .B1(n7904), .B2(n12579), .ZN(
        n5094) );
  OAI22_X1 U4748 ( .A1(n12585), .A2(n13295), .B1(n7887), .B2(n12579), .ZN(
        n5095) );
  OAI22_X1 U4749 ( .A1(n12585), .A2(n13298), .B1(n7870), .B2(n12579), .ZN(
        n5096) );
  OAI22_X1 U4750 ( .A1(n12585), .A2(n13301), .B1(n7853), .B2(n12579), .ZN(
        n5097) );
  OAI22_X1 U4751 ( .A1(n12584), .A2(n13304), .B1(n7836), .B2(n12579), .ZN(
        n5098) );
  OAI22_X1 U4752 ( .A1(n12584), .A2(n13307), .B1(n7819), .B2(n12579), .ZN(
        n5099) );
  OAI22_X1 U4753 ( .A1(n12584), .A2(n13310), .B1(n7802), .B2(n12579), .ZN(
        n5100) );
  OAI22_X1 U4754 ( .A1(n12584), .A2(n13313), .B1(n7785), .B2(n12579), .ZN(
        n5101) );
  OAI22_X1 U4755 ( .A1(n12584), .A2(n13316), .B1(n7768), .B2(n12580), .ZN(
        n5102) );
  OAI22_X1 U4756 ( .A1(n12583), .A2(n13319), .B1(n7751), .B2(n12580), .ZN(
        n5103) );
  OAI22_X1 U4757 ( .A1(n12583), .A2(n13322), .B1(n7649), .B2(n12580), .ZN(
        n5104) );
  OAI22_X1 U4758 ( .A1(n12583), .A2(n13325), .B1(n7632), .B2(n12580), .ZN(
        n5105) );
  OAI22_X1 U4759 ( .A1(n12583), .A2(n13328), .B1(n7528), .B2(n12580), .ZN(
        n5106) );
  OAI22_X1 U4760 ( .A1(n12583), .A2(n13331), .B1(n7511), .B2(n12580), .ZN(
        n5107) );
  OAI22_X1 U4761 ( .A1(n12582), .A2(n13334), .B1(n7494), .B2(n12580), .ZN(
        n5108) );
  OAI22_X1 U4762 ( .A1(n12582), .A2(n13337), .B1(n7392), .B2(n12580), .ZN(
        n5109) );
  OAI22_X1 U4763 ( .A1(n12582), .A2(n13340), .B1(n7375), .B2(n12580), .ZN(
        n5110) );
  OAI22_X1 U4764 ( .A1(n12582), .A2(n13343), .B1(n7276), .B2(n12580), .ZN(
        n5111) );
  OAI22_X1 U4765 ( .A1(n12582), .A2(n13346), .B1(n7259), .B2(n12580), .ZN(
        n5112) );
  OAI22_X1 U4766 ( .A1(n12581), .A2(n13349), .B1(n7242), .B2(n12580), .ZN(
        n5113) );
  OAI22_X1 U4767 ( .A1(n12645), .A2(n13244), .B1(n8173), .B2(n12635), .ZN(
        n5270) );
  OAI22_X1 U4768 ( .A1(n12645), .A2(n13247), .B1(n8156), .B2(n12635), .ZN(
        n5271) );
  OAI22_X1 U4769 ( .A1(n12645), .A2(n13250), .B1(n8139), .B2(n12635), .ZN(
        n5272) );
  OAI22_X1 U4770 ( .A1(n12645), .A2(n13253), .B1(n8122), .B2(n12635), .ZN(
        n5273) );
  OAI22_X1 U4771 ( .A1(n12645), .A2(n13256), .B1(n8105), .B2(n12635), .ZN(
        n5274) );
  OAI22_X1 U4772 ( .A1(n12644), .A2(n13259), .B1(n8088), .B2(n12635), .ZN(
        n5275) );
  OAI22_X1 U4773 ( .A1(n12644), .A2(n13262), .B1(n8071), .B2(n12635), .ZN(
        n5276) );
  OAI22_X1 U4774 ( .A1(n12644), .A2(n13265), .B1(n8054), .B2(n12635), .ZN(
        n5277) );
  OAI22_X1 U4775 ( .A1(n12644), .A2(n13268), .B1(n8037), .B2(n12635), .ZN(
        n5278) );
  OAI22_X1 U4776 ( .A1(n12644), .A2(n13271), .B1(n8020), .B2(n12635), .ZN(
        n5279) );
  OAI22_X1 U4777 ( .A1(n12643), .A2(n13274), .B1(n8003), .B2(n12635), .ZN(
        n5280) );
  OAI22_X1 U4778 ( .A1(n12643), .A2(n13277), .B1(n7986), .B2(n12635), .ZN(
        n5281) );
  OAI22_X1 U4779 ( .A1(n12643), .A2(n13280), .B1(n7969), .B2(n12636), .ZN(
        n5282) );
  OAI22_X1 U4780 ( .A1(n12643), .A2(n13283), .B1(n7952), .B2(n12636), .ZN(
        n5283) );
  OAI22_X1 U4781 ( .A1(n12643), .A2(n13286), .B1(n7935), .B2(n12636), .ZN(
        n5284) );
  OAI22_X1 U4782 ( .A1(n12642), .A2(n13289), .B1(n7918), .B2(n12636), .ZN(
        n5285) );
  OAI22_X1 U4783 ( .A1(n12642), .A2(n13292), .B1(n7901), .B2(n12636), .ZN(
        n5286) );
  OAI22_X1 U4784 ( .A1(n12642), .A2(n13295), .B1(n7884), .B2(n12636), .ZN(
        n5287) );
  OAI22_X1 U4785 ( .A1(n12642), .A2(n13298), .B1(n7867), .B2(n12636), .ZN(
        n5288) );
  OAI22_X1 U4786 ( .A1(n12642), .A2(n13301), .B1(n7850), .B2(n12636), .ZN(
        n5289) );
  OAI22_X1 U4787 ( .A1(n12641), .A2(n13304), .B1(n7833), .B2(n12636), .ZN(
        n5290) );
  OAI22_X1 U4788 ( .A1(n12641), .A2(n13307), .B1(n7816), .B2(n12636), .ZN(
        n5291) );
  OAI22_X1 U4789 ( .A1(n12641), .A2(n13310), .B1(n7799), .B2(n12636), .ZN(
        n5292) );
  OAI22_X1 U4790 ( .A1(n12641), .A2(n13313), .B1(n7782), .B2(n12636), .ZN(
        n5293) );
  OAI22_X1 U4791 ( .A1(n12641), .A2(n13316), .B1(n7765), .B2(n12637), .ZN(
        n5294) );
  OAI22_X1 U4792 ( .A1(n12640), .A2(n13319), .B1(n7748), .B2(n12637), .ZN(
        n5295) );
  OAI22_X1 U4793 ( .A1(n12640), .A2(n13322), .B1(n7646), .B2(n12637), .ZN(
        n5296) );
  OAI22_X1 U4794 ( .A1(n12640), .A2(n13325), .B1(n7629), .B2(n12637), .ZN(
        n5297) );
  OAI22_X1 U4795 ( .A1(n12640), .A2(n13328), .B1(n7525), .B2(n12637), .ZN(
        n5298) );
  OAI22_X1 U4796 ( .A1(n12640), .A2(n13331), .B1(n7508), .B2(n12637), .ZN(
        n5299) );
  OAI22_X1 U4797 ( .A1(n12639), .A2(n13334), .B1(n7491), .B2(n12637), .ZN(
        n5300) );
  OAI22_X1 U4798 ( .A1(n12639), .A2(n13337), .B1(n7389), .B2(n12637), .ZN(
        n5301) );
  OAI22_X1 U4799 ( .A1(n12639), .A2(n13340), .B1(n7372), .B2(n12637), .ZN(
        n5302) );
  OAI22_X1 U4800 ( .A1(n12639), .A2(n13343), .B1(n7273), .B2(n12637), .ZN(
        n5303) );
  OAI22_X1 U4801 ( .A1(n12639), .A2(n13346), .B1(n7256), .B2(n12637), .ZN(
        n5304) );
  OAI22_X1 U4802 ( .A1(n12638), .A2(n13349), .B1(n7239), .B2(n12637), .ZN(
        n5305) );
  OAI22_X1 U4803 ( .A1(n12664), .A2(n13244), .B1(n8174), .B2(n12654), .ZN(
        n5334) );
  OAI22_X1 U4804 ( .A1(n12664), .A2(n13247), .B1(n8157), .B2(n12654), .ZN(
        n5335) );
  OAI22_X1 U4805 ( .A1(n12664), .A2(n13250), .B1(n8140), .B2(n12654), .ZN(
        n5336) );
  OAI22_X1 U4806 ( .A1(n12664), .A2(n13253), .B1(n8123), .B2(n12654), .ZN(
        n5337) );
  OAI22_X1 U4807 ( .A1(n12664), .A2(n13256), .B1(n8106), .B2(n12654), .ZN(
        n5338) );
  OAI22_X1 U4808 ( .A1(n12663), .A2(n13259), .B1(n8089), .B2(n12654), .ZN(
        n5339) );
  OAI22_X1 U4809 ( .A1(n12663), .A2(n13262), .B1(n8072), .B2(n12654), .ZN(
        n5340) );
  OAI22_X1 U4810 ( .A1(n12663), .A2(n13265), .B1(n8055), .B2(n12654), .ZN(
        n5341) );
  OAI22_X1 U4811 ( .A1(n12663), .A2(n13268), .B1(n8038), .B2(n12654), .ZN(
        n5342) );
  OAI22_X1 U4812 ( .A1(n12663), .A2(n13271), .B1(n8021), .B2(n12654), .ZN(
        n5343) );
  OAI22_X1 U4813 ( .A1(n12662), .A2(n13274), .B1(n8004), .B2(n12654), .ZN(
        n5344) );
  OAI22_X1 U4814 ( .A1(n12662), .A2(n13277), .B1(n7987), .B2(n12654), .ZN(
        n5345) );
  OAI22_X1 U4815 ( .A1(n12662), .A2(n13280), .B1(n7970), .B2(n12655), .ZN(
        n5346) );
  OAI22_X1 U4816 ( .A1(n12662), .A2(n13283), .B1(n7953), .B2(n12655), .ZN(
        n5347) );
  OAI22_X1 U4817 ( .A1(n12662), .A2(n13286), .B1(n7936), .B2(n12655), .ZN(
        n5348) );
  OAI22_X1 U4818 ( .A1(n12661), .A2(n13289), .B1(n7919), .B2(n12655), .ZN(
        n5349) );
  OAI22_X1 U4819 ( .A1(n12661), .A2(n13292), .B1(n7902), .B2(n12655), .ZN(
        n5350) );
  OAI22_X1 U4820 ( .A1(n12661), .A2(n13295), .B1(n7885), .B2(n12655), .ZN(
        n5351) );
  OAI22_X1 U4821 ( .A1(n12661), .A2(n13298), .B1(n7868), .B2(n12655), .ZN(
        n5352) );
  OAI22_X1 U4822 ( .A1(n12661), .A2(n13301), .B1(n7851), .B2(n12655), .ZN(
        n5353) );
  OAI22_X1 U4823 ( .A1(n12660), .A2(n13304), .B1(n7834), .B2(n12655), .ZN(
        n5354) );
  OAI22_X1 U4824 ( .A1(n12660), .A2(n13307), .B1(n7817), .B2(n12655), .ZN(
        n5355) );
  OAI22_X1 U4825 ( .A1(n12660), .A2(n13310), .B1(n7800), .B2(n12655), .ZN(
        n5356) );
  OAI22_X1 U4826 ( .A1(n12660), .A2(n13313), .B1(n7783), .B2(n12655), .ZN(
        n5357) );
  OAI22_X1 U4827 ( .A1(n12660), .A2(n13316), .B1(n7766), .B2(n12656), .ZN(
        n5358) );
  OAI22_X1 U4828 ( .A1(n12659), .A2(n13319), .B1(n7749), .B2(n12656), .ZN(
        n5359) );
  OAI22_X1 U4829 ( .A1(n12659), .A2(n13322), .B1(n7647), .B2(n12656), .ZN(
        n5360) );
  OAI22_X1 U4830 ( .A1(n12659), .A2(n13325), .B1(n7630), .B2(n12656), .ZN(
        n5361) );
  OAI22_X1 U4831 ( .A1(n12659), .A2(n13328), .B1(n7526), .B2(n12656), .ZN(
        n5362) );
  OAI22_X1 U4832 ( .A1(n12659), .A2(n13331), .B1(n7509), .B2(n12656), .ZN(
        n5363) );
  OAI22_X1 U4833 ( .A1(n12658), .A2(n13334), .B1(n7492), .B2(n12656), .ZN(
        n5364) );
  OAI22_X1 U4834 ( .A1(n12658), .A2(n13337), .B1(n7390), .B2(n12656), .ZN(
        n5365) );
  OAI22_X1 U4835 ( .A1(n12658), .A2(n13340), .B1(n7373), .B2(n12656), .ZN(
        n5366) );
  OAI22_X1 U4836 ( .A1(n12658), .A2(n13343), .B1(n7274), .B2(n12656), .ZN(
        n5367) );
  OAI22_X1 U4837 ( .A1(n12658), .A2(n13346), .B1(n7257), .B2(n12656), .ZN(
        n5368) );
  OAI22_X1 U4838 ( .A1(n12657), .A2(n13349), .B1(n7240), .B2(n12656), .ZN(
        n5369) );
  OAI22_X1 U4839 ( .A1(n12855), .A2(n13351), .B1(n7139), .B2(n12852), .ZN(
        n6010) );
  OAI22_X1 U4840 ( .A1(n12855), .A2(n13354), .B1(n7122), .B2(n12853), .ZN(
        n6011) );
  OAI22_X1 U4841 ( .A1(n12855), .A2(n13357), .B1(n4861), .B2(n12854), .ZN(
        n6012) );
  OAI22_X1 U4842 ( .A1(n12855), .A2(n13380), .B1(n4844), .B2(n12852), .ZN(
        n6013) );
  OAI22_X1 U4843 ( .A1(n12775), .A2(n13351), .B1(n7141), .B2(n12772), .ZN(
        n5754) );
  OAI22_X1 U4844 ( .A1(n12775), .A2(n13354), .B1(n7124), .B2(n12773), .ZN(
        n5755) );
  OAI22_X1 U4845 ( .A1(n12775), .A2(n13357), .B1(n7107), .B2(n12774), .ZN(
        n5756) );
  OAI22_X1 U4846 ( .A1(n12775), .A2(n13380), .B1(n4846), .B2(n12772), .ZN(
        n5757) );
  OAI22_X1 U4847 ( .A1(n12835), .A2(n13351), .B1(n7138), .B2(n12832), .ZN(
        n5946) );
  OAI22_X1 U4848 ( .A1(n12835), .A2(n13354), .B1(n7121), .B2(n12833), .ZN(
        n5947) );
  OAI22_X1 U4849 ( .A1(n12835), .A2(n13357), .B1(n4860), .B2(n12834), .ZN(
        n5948) );
  OAI22_X1 U4850 ( .A1(n12835), .A2(n13380), .B1(n4843), .B2(n12832), .ZN(
        n5949) );
  OAI22_X1 U4851 ( .A1(n12755), .A2(n13351), .B1(n7140), .B2(n12752), .ZN(
        n5690) );
  OAI22_X1 U4852 ( .A1(n12755), .A2(n13354), .B1(n7123), .B2(n12753), .ZN(
        n5691) );
  OAI22_X1 U4853 ( .A1(n12755), .A2(n13357), .B1(n7106), .B2(n12754), .ZN(
        n5692) );
  OAI22_X1 U4854 ( .A1(n12755), .A2(n13380), .B1(n4845), .B2(n12752), .ZN(
        n5693) );
  OAI22_X1 U4855 ( .A1(n13125), .A2(n13206), .B1(n8366), .B2(n13111), .ZN(
        n6794) );
  OAI22_X1 U4856 ( .A1(n12947), .A2(n13171), .B1(n8576), .B2(n12933), .ZN(
        n6206) );
  OAI22_X1 U4857 ( .A1(n12947), .A2(n13174), .B1(n8559), .B2(n12934), .ZN(
        n6207) );
  OAI22_X1 U4858 ( .A1(n12947), .A2(n13177), .B1(n8542), .B2(n12931), .ZN(
        n6208) );
  OAI22_X1 U4859 ( .A1(n12947), .A2(n13180), .B1(n8525), .B2(n12933), .ZN(
        n6209) );
  OAI22_X1 U4860 ( .A1(n12946), .A2(n13183), .B1(n8508), .B2(n12934), .ZN(
        n6210) );
  OAI22_X1 U4861 ( .A1(n12946), .A2(n13186), .B1(n8491), .B2(n12930), .ZN(
        n6211) );
  OAI22_X1 U4862 ( .A1(n12945), .A2(n13210), .B1(n8355), .B2(n12931), .ZN(
        n6219) );
  OAI22_X1 U4863 ( .A1(n12944), .A2(n13213), .B1(n8338), .B2(n12931), .ZN(
        n6220) );
  OAI22_X1 U4864 ( .A1(n12944), .A2(n13216), .B1(n8321), .B2(n12931), .ZN(
        n6221) );
  OAI22_X1 U4865 ( .A1(n12944), .A2(n13219), .B1(n8304), .B2(n12931), .ZN(
        n6222) );
  OAI22_X1 U4866 ( .A1(n12944), .A2(n13222), .B1(n8287), .B2(n12931), .ZN(
        n6223) );
  OAI22_X1 U4867 ( .A1(n12944), .A2(n13225), .B1(n8270), .B2(n12931), .ZN(
        n6224) );
  OAI22_X1 U4868 ( .A1(n12915), .A2(n13351), .B1(n7136), .B2(n12912), .ZN(
        n6202) );
  OAI22_X1 U4869 ( .A1(n12915), .A2(n13354), .B1(n7119), .B2(n12913), .ZN(
        n6203) );
  OAI22_X1 U4870 ( .A1(n12915), .A2(n13357), .B1(n4858), .B2(n12914), .ZN(
        n6204) );
  OAI22_X1 U4871 ( .A1(n12915), .A2(n13380), .B1(n4841), .B2(n12912), .ZN(
        n6205) );
  OAI22_X1 U4872 ( .A1(n12935), .A2(n13351), .B1(n7137), .B2(n12932), .ZN(
        n6266) );
  OAI22_X1 U4873 ( .A1(n12935), .A2(n13354), .B1(n7120), .B2(n12933), .ZN(
        n6267) );
  OAI22_X1 U4874 ( .A1(n12935), .A2(n13357), .B1(n4859), .B2(n12934), .ZN(
        n6268) );
  OAI22_X1 U4875 ( .A1(n12935), .A2(n13380), .B1(n4842), .B2(n12932), .ZN(
        n6269) );
  OAI22_X1 U4876 ( .A1(n13015), .A2(n13350), .B1(n7135), .B2(n13012), .ZN(
        n6522) );
  OAI22_X1 U4877 ( .A1(n13015), .A2(n13353), .B1(n7118), .B2(n13013), .ZN(
        n6523) );
  OAI22_X1 U4878 ( .A1(n13015), .A2(n13356), .B1(n4857), .B2(n13014), .ZN(
        n6524) );
  OAI22_X1 U4879 ( .A1(n13015), .A2(n13379), .B1(n4840), .B2(n13012), .ZN(
        n6525) );
  OAI22_X1 U4880 ( .A1(n12995), .A2(n13350), .B1(n7134), .B2(n12992), .ZN(
        n6458) );
  OAI22_X1 U4881 ( .A1(n12995), .A2(n13353), .B1(n7117), .B2(n12993), .ZN(
        n6459) );
  OAI22_X1 U4882 ( .A1(n12995), .A2(n13356), .B1(n4856), .B2(n12994), .ZN(
        n6460) );
  OAI22_X1 U4883 ( .A1(n12995), .A2(n13379), .B1(n4839), .B2(n12992), .ZN(
        n6461) );
  OAI22_X1 U4884 ( .A1(n13055), .A2(n13350), .B1(n7132), .B2(n13052), .ZN(
        n6650) );
  OAI22_X1 U4885 ( .A1(n13055), .A2(n13353), .B1(n7115), .B2(n13053), .ZN(
        n6651) );
  OAI22_X1 U4886 ( .A1(n13055), .A2(n13356), .B1(n4854), .B2(n13054), .ZN(
        n6652) );
  OAI22_X1 U4887 ( .A1(n13055), .A2(n13379), .B1(n4837), .B2(n13052), .ZN(
        n6653) );
  OAI22_X1 U4888 ( .A1(n13035), .A2(n13350), .B1(n7133), .B2(n13032), .ZN(
        n6586) );
  OAI22_X1 U4889 ( .A1(n13035), .A2(n13353), .B1(n7116), .B2(n13033), .ZN(
        n6587) );
  OAI22_X1 U4890 ( .A1(n13035), .A2(n13356), .B1(n4855), .B2(n13034), .ZN(
        n6588) );
  OAI22_X1 U4891 ( .A1(n13035), .A2(n13379), .B1(n4838), .B2(n13032), .ZN(
        n6589) );
  OAI22_X1 U4892 ( .A1(n12581), .A2(n13352), .B1(n7145), .B2(n12578), .ZN(
        n5114) );
  OAI22_X1 U4893 ( .A1(n12581), .A2(n13355), .B1(n7128), .B2(n12579), .ZN(
        n5115) );
  OAI22_X1 U4894 ( .A1(n12581), .A2(n13358), .B1(n7111), .B2(n12580), .ZN(
        n5116) );
  OAI22_X1 U4895 ( .A1(n12581), .A2(n13381), .B1(n4850), .B2(n12578), .ZN(
        n5117) );
  OAI22_X1 U4896 ( .A1(n12638), .A2(n13352), .B1(n7142), .B2(n12635), .ZN(
        n5306) );
  OAI22_X1 U4897 ( .A1(n12638), .A2(n13355), .B1(n7125), .B2(n12636), .ZN(
        n5307) );
  OAI22_X1 U4898 ( .A1(n12638), .A2(n13358), .B1(n7108), .B2(n12637), .ZN(
        n5308) );
  OAI22_X1 U4899 ( .A1(n12638), .A2(n13381), .B1(n4847), .B2(n12635), .ZN(
        n5309) );
  OAI22_X1 U4900 ( .A1(n12657), .A2(n13352), .B1(n7143), .B2(n12654), .ZN(
        n5370) );
  OAI22_X1 U4901 ( .A1(n12657), .A2(n13355), .B1(n7126), .B2(n12655), .ZN(
        n5371) );
  OAI22_X1 U4902 ( .A1(n12657), .A2(n13358), .B1(n7109), .B2(n12656), .ZN(
        n5372) );
  OAI22_X1 U4903 ( .A1(n12657), .A2(n13381), .B1(n4848), .B2(n12654), .ZN(
        n5373) );
  OAI22_X1 U4904 ( .A1(n13115), .A2(n13379), .B1(n13112), .B2(n13848), .ZN(
        n6845) );
  OAI22_X1 U4905 ( .A1(n13135), .A2(n13350), .B1(n13132), .B2(n13852), .ZN(
        n6906) );
  OAI22_X1 U4906 ( .A1(n13135), .A2(n13353), .B1(n13133), .B2(n13851), .ZN(
        n6907) );
  OAI22_X1 U4907 ( .A1(n13135), .A2(n13356), .B1(n13134), .B2(n13850), .ZN(
        n6908) );
  OAI22_X1 U4908 ( .A1(n13135), .A2(n13379), .B1(n13132), .B2(n13849), .ZN(
        n6909) );
  OAI22_X1 U4909 ( .A1(n12715), .A2(n13351), .B1(n12713), .B2(n13666), .ZN(
        n5562) );
  OAI22_X1 U4910 ( .A1(n12715), .A2(n13354), .B1(n12712), .B2(n13665), .ZN(
        n5563) );
  OAI22_X1 U4911 ( .A1(n12715), .A2(n13357), .B1(n12714), .B2(n13664), .ZN(
        n5564) );
  OAI22_X1 U4912 ( .A1(n12715), .A2(n13380), .B1(n12713), .B2(n13663), .ZN(
        n5565) );
  OAI22_X1 U4913 ( .A1(n12735), .A2(n13351), .B1(n12732), .B2(n13662), .ZN(
        n5626) );
  OAI22_X1 U4914 ( .A1(n12735), .A2(n13354), .B1(n12733), .B2(n13661), .ZN(
        n5627) );
  OAI22_X1 U4915 ( .A1(n12735), .A2(n13357), .B1(n12734), .B2(n13660), .ZN(
        n5628) );
  OAI22_X1 U4916 ( .A1(n12735), .A2(n13380), .B1(n12732), .B2(n13659), .ZN(
        n5629) );
  OAI22_X1 U4917 ( .A1(n12795), .A2(n13351), .B1(n12792), .B2(n13658), .ZN(
        n5818) );
  OAI22_X1 U4918 ( .A1(n12795), .A2(n13354), .B1(n12793), .B2(n13657), .ZN(
        n5819) );
  OAI22_X1 U4919 ( .A1(n12795), .A2(n13357), .B1(n12794), .B2(n13656), .ZN(
        n5820) );
  OAI22_X1 U4920 ( .A1(n12795), .A2(n13380), .B1(n12792), .B2(n13655), .ZN(
        n5821) );
  OAI22_X1 U4921 ( .A1(n12815), .A2(n13351), .B1(n12812), .B2(n13654), .ZN(
        n5882) );
  OAI22_X1 U4922 ( .A1(n12815), .A2(n13354), .B1(n12813), .B2(n13653), .ZN(
        n5883) );
  OAI22_X1 U4923 ( .A1(n12815), .A2(n13357), .B1(n12814), .B2(n13652), .ZN(
        n5884) );
  OAI22_X1 U4924 ( .A1(n12815), .A2(n13380), .B1(n12812), .B2(n13651), .ZN(
        n5885) );
  OAI21_X1 U4925 ( .B1(n4833), .B2(n12544), .A(n3180), .ZN(n4926) );
  OAI21_X1 U4926 ( .B1(n3181), .B2(n3182), .A(n12549), .ZN(n3180) );
  NAND4_X1 U4927 ( .A1(n3183), .A2(n3184), .A3(n3185), .A4(n3186), .ZN(n3182)
         );
  NAND4_X1 U4928 ( .A1(n3199), .A2(n3200), .A3(n3201), .A4(n3202), .ZN(n3181)
         );
  OAI21_X1 U4929 ( .B1(n4832), .B2(n12543), .A(n3161), .ZN(n4927) );
  OAI21_X1 U4930 ( .B1(n3162), .B2(n3163), .A(n12549), .ZN(n3161) );
  NAND4_X1 U4931 ( .A1(n3164), .A2(n3165), .A3(n3166), .A4(n3167), .ZN(n3163)
         );
  NAND4_X1 U4932 ( .A1(n3172), .A2(n3173), .A3(n3174), .A4(n3175), .ZN(n3162)
         );
  OAI21_X1 U4933 ( .B1(n4831), .B2(n12544), .A(n3142), .ZN(n4928) );
  OAI21_X1 U4934 ( .B1(n3143), .B2(n3144), .A(n12549), .ZN(n3142) );
  NAND4_X1 U4935 ( .A1(n3145), .A2(n3146), .A3(n3147), .A4(n3148), .ZN(n3144)
         );
  NAND4_X1 U4936 ( .A1(n3153), .A2(n3154), .A3(n3155), .A4(n3156), .ZN(n3143)
         );
  OAI21_X1 U4937 ( .B1(n4830), .B2(n12543), .A(n3123), .ZN(n4929) );
  OAI21_X1 U4938 ( .B1(n3124), .B2(n3125), .A(n12548), .ZN(n3123) );
  NAND4_X1 U4939 ( .A1(n3126), .A2(n3127), .A3(n3128), .A4(n3129), .ZN(n3125)
         );
  NAND4_X1 U4940 ( .A1(n3134), .A2(n3135), .A3(n3136), .A4(n3137), .ZN(n3124)
         );
  OAI21_X1 U4941 ( .B1(n4829), .B2(n12543), .A(n3104), .ZN(n4930) );
  OAI21_X1 U4942 ( .B1(n3105), .B2(n3106), .A(n12548), .ZN(n3104) );
  NAND4_X1 U4943 ( .A1(n3107), .A2(n3108), .A3(n3109), .A4(n3110), .ZN(n3106)
         );
  NAND4_X1 U4944 ( .A1(n3115), .A2(n3116), .A3(n3117), .A4(n3118), .ZN(n3105)
         );
  OAI21_X1 U4945 ( .B1(n4828), .B2(n12544), .A(n3085), .ZN(n4931) );
  OAI21_X1 U4946 ( .B1(n3086), .B2(n3087), .A(n12548), .ZN(n3085) );
  NAND4_X1 U4947 ( .A1(n3088), .A2(n3089), .A3(n3090), .A4(n3091), .ZN(n3087)
         );
  NAND4_X1 U4948 ( .A1(n3096), .A2(n3097), .A3(n3098), .A4(n3099), .ZN(n3086)
         );
  OAI21_X1 U4949 ( .B1(n4827), .B2(n12544), .A(n3066), .ZN(n4932) );
  OAI21_X1 U4950 ( .B1(n3067), .B2(n3068), .A(n12548), .ZN(n3066) );
  NAND4_X1 U4951 ( .A1(n3069), .A2(n3070), .A3(n3071), .A4(n3072), .ZN(n3068)
         );
  NAND4_X1 U4952 ( .A1(n3077), .A2(n3078), .A3(n3079), .A4(n3080), .ZN(n3067)
         );
  OAI21_X1 U4953 ( .B1(n4826), .B2(n12543), .A(n3047), .ZN(n4933) );
  OAI21_X1 U4954 ( .B1(n3048), .B2(n3049), .A(n12548), .ZN(n3047) );
  NAND4_X1 U4955 ( .A1(n3050), .A2(n3051), .A3(n3052), .A4(n3053), .ZN(n3049)
         );
  NAND4_X1 U4956 ( .A1(n3058), .A2(n3059), .A3(n3060), .A4(n3061), .ZN(n3048)
         );
  OAI21_X1 U4957 ( .B1(n4825), .B2(n12543), .A(n3028), .ZN(n4934) );
  OAI21_X1 U4958 ( .B1(n3029), .B2(n3030), .A(n12547), .ZN(n3028) );
  NAND4_X1 U4959 ( .A1(n3031), .A2(n3032), .A3(n3033), .A4(n3034), .ZN(n3030)
         );
  NAND4_X1 U4960 ( .A1(n3039), .A2(n3040), .A3(n3041), .A4(n3042), .ZN(n3029)
         );
  OAI21_X1 U4961 ( .B1(n4824), .B2(n12543), .A(n3009), .ZN(n4935) );
  OAI21_X1 U4962 ( .B1(n3010), .B2(n3011), .A(n12547), .ZN(n3009) );
  NAND4_X1 U4963 ( .A1(n3012), .A2(n3013), .A3(n3014), .A4(n3015), .ZN(n3011)
         );
  NAND4_X1 U4964 ( .A1(n3020), .A2(n3021), .A3(n3022), .A4(n3023), .ZN(n3010)
         );
  OAI21_X1 U4965 ( .B1(n4823), .B2(n12542), .A(n2990), .ZN(n4936) );
  OAI21_X1 U4966 ( .B1(n2991), .B2(n2992), .A(n12546), .ZN(n2990) );
  NAND4_X1 U4967 ( .A1(n2993), .A2(n2994), .A3(n2995), .A4(n2996), .ZN(n2992)
         );
  NAND4_X1 U4968 ( .A1(n3001), .A2(n3002), .A3(n3003), .A4(n3004), .ZN(n2991)
         );
  OAI21_X1 U4969 ( .B1(n4822), .B2(n12543), .A(n2971), .ZN(n4937) );
  OAI21_X1 U4970 ( .B1(n2972), .B2(n2973), .A(n12546), .ZN(n2971) );
  NAND4_X1 U4971 ( .A1(n2974), .A2(n2975), .A3(n2976), .A4(n2977), .ZN(n2973)
         );
  NAND4_X1 U4972 ( .A1(n2982), .A2(n2983), .A3(n2984), .A4(n2985), .ZN(n2972)
         );
  OAI21_X1 U4973 ( .B1(n4821), .B2(n12543), .A(n2952), .ZN(n4938) );
  OAI21_X1 U4974 ( .B1(n2953), .B2(n2954), .A(n12546), .ZN(n2952) );
  NAND4_X1 U4975 ( .A1(n2955), .A2(n2956), .A3(n2957), .A4(n2958), .ZN(n2954)
         );
  NAND4_X1 U4976 ( .A1(n2963), .A2(n2964), .A3(n2965), .A4(n2966), .ZN(n2953)
         );
  OAI21_X1 U4977 ( .B1(n4820), .B2(n12543), .A(n2933), .ZN(n4939) );
  OAI21_X1 U4978 ( .B1(n2934), .B2(n2935), .A(n12545), .ZN(n2933) );
  NAND4_X1 U4979 ( .A1(n2936), .A2(n2937), .A3(n2938), .A4(n2939), .ZN(n2935)
         );
  NAND4_X1 U4980 ( .A1(n2944), .A2(n2945), .A3(n2946), .A4(n2947), .ZN(n2934)
         );
  OAI21_X1 U4981 ( .B1(n4819), .B2(n12543), .A(n2914), .ZN(n4940) );
  OAI21_X1 U4982 ( .B1(n2915), .B2(n2916), .A(n12547), .ZN(n2914) );
  NAND4_X1 U4983 ( .A1(n2917), .A2(n2918), .A3(n2919), .A4(n2920), .ZN(n2916)
         );
  NAND4_X1 U4984 ( .A1(n2925), .A2(n2926), .A3(n2927), .A4(n2928), .ZN(n2915)
         );
  OAI21_X1 U4985 ( .B1(n4818), .B2(n12543), .A(n2895), .ZN(n4941) );
  OAI21_X1 U4986 ( .B1(n2896), .B2(n2897), .A(n12546), .ZN(n2895) );
  NAND4_X1 U4987 ( .A1(n2898), .A2(n2899), .A3(n2900), .A4(n2901), .ZN(n2897)
         );
  NAND4_X1 U4988 ( .A1(n2906), .A2(n2907), .A3(n2908), .A4(n2909), .ZN(n2896)
         );
  OAI21_X1 U4989 ( .B1(n4817), .B2(n12542), .A(n2876), .ZN(n4942) );
  OAI21_X1 U4990 ( .B1(n2877), .B2(n2878), .A(n12544), .ZN(n2876) );
  NAND4_X1 U4991 ( .A1(n2879), .A2(n2880), .A3(n2881), .A4(n2882), .ZN(n2878)
         );
  NAND4_X1 U4992 ( .A1(n2887), .A2(n2888), .A3(n2889), .A4(n2890), .ZN(n2877)
         );
  OAI21_X1 U4993 ( .B1(n4816), .B2(n12542), .A(n2857), .ZN(n4943) );
  OAI21_X1 U4994 ( .B1(n2858), .B2(n2859), .A(n12546), .ZN(n2857) );
  NAND4_X1 U4995 ( .A1(n2860), .A2(n2861), .A3(n2862), .A4(n2863), .ZN(n2859)
         );
  NAND4_X1 U4996 ( .A1(n2868), .A2(n2869), .A3(n2870), .A4(n2871), .ZN(n2858)
         );
  OAI21_X1 U4997 ( .B1(n4815), .B2(n12543), .A(n2838), .ZN(n4944) );
  OAI21_X1 U4998 ( .B1(n2839), .B2(n2840), .A(n12545), .ZN(n2838) );
  NAND4_X1 U4999 ( .A1(n2841), .A2(n2842), .A3(n2843), .A4(n2844), .ZN(n2840)
         );
  NAND4_X1 U5000 ( .A1(n2849), .A2(n2850), .A3(n2851), .A4(n2852), .ZN(n2839)
         );
  OAI21_X1 U5001 ( .B1(n4814), .B2(n12542), .A(n2819), .ZN(n4945) );
  OAI21_X1 U5002 ( .B1(n2820), .B2(n2821), .A(n12546), .ZN(n2819) );
  NAND4_X1 U5003 ( .A1(n2822), .A2(n2823), .A3(n2824), .A4(n2825), .ZN(n2821)
         );
  NAND4_X1 U5004 ( .A1(n2830), .A2(n2831), .A3(n2832), .A4(n2833), .ZN(n2820)
         );
  OAI21_X1 U5005 ( .B1(n4813), .B2(n12542), .A(n2800), .ZN(n4946) );
  OAI21_X1 U5006 ( .B1(n2801), .B2(n2802), .A(n12544), .ZN(n2800) );
  NAND4_X1 U5007 ( .A1(n2803), .A2(n2804), .A3(n2805), .A4(n2806), .ZN(n2802)
         );
  NAND4_X1 U5008 ( .A1(n2811), .A2(n2812), .A3(n2813), .A4(n2814), .ZN(n2801)
         );
  OAI21_X1 U5009 ( .B1(n4812), .B2(n12542), .A(n2781), .ZN(n4947) );
  OAI21_X1 U5010 ( .B1(n2782), .B2(n2783), .A(n12545), .ZN(n2781) );
  NAND4_X1 U5011 ( .A1(n2784), .A2(n2785), .A3(n2786), .A4(n2787), .ZN(n2783)
         );
  NAND4_X1 U5012 ( .A1(n2792), .A2(n2793), .A3(n2794), .A4(n2795), .ZN(n2782)
         );
  OAI21_X1 U5013 ( .B1(n4811), .B2(n12542), .A(n2762), .ZN(n4948) );
  OAI21_X1 U5014 ( .B1(n2763), .B2(n2764), .A(n12544), .ZN(n2762) );
  NAND4_X1 U5015 ( .A1(n2765), .A2(n2766), .A3(n2767), .A4(n2768), .ZN(n2764)
         );
  NAND4_X1 U5016 ( .A1(n2773), .A2(n2774), .A3(n2775), .A4(n2776), .ZN(n2763)
         );
  OAI21_X1 U5017 ( .B1(n4810), .B2(n12542), .A(n2743), .ZN(n4949) );
  OAI21_X1 U5018 ( .B1(n2744), .B2(n2745), .A(n12545), .ZN(n2743) );
  NAND4_X1 U5019 ( .A1(n2746), .A2(n2747), .A3(n2748), .A4(n2749), .ZN(n2745)
         );
  NAND4_X1 U5020 ( .A1(n2754), .A2(n2755), .A3(n2756), .A4(n2757), .ZN(n2744)
         );
  OAI21_X1 U5021 ( .B1(n4809), .B2(n12542), .A(n2724), .ZN(n4950) );
  OAI21_X1 U5022 ( .B1(n2725), .B2(n2726), .A(n12544), .ZN(n2724) );
  NAND4_X1 U5023 ( .A1(n2727), .A2(n2728), .A3(n2729), .A4(n2730), .ZN(n2726)
         );
  NAND4_X1 U5024 ( .A1(n2735), .A2(n2736), .A3(n2737), .A4(n2738), .ZN(n2725)
         );
  OAI21_X1 U5025 ( .B1(n4808), .B2(n12542), .A(n2705), .ZN(n4951) );
  OAI21_X1 U5026 ( .B1(n2706), .B2(n2707), .A(n12545), .ZN(n2705) );
  NAND4_X1 U5027 ( .A1(n2708), .A2(n2709), .A3(n2710), .A4(n2711), .ZN(n2707)
         );
  NAND4_X1 U5028 ( .A1(n2716), .A2(n2717), .A3(n2718), .A4(n2719), .ZN(n2706)
         );
  OAI21_X1 U5029 ( .B1(n4807), .B2(n12542), .A(n2686), .ZN(n4952) );
  OAI21_X1 U5030 ( .B1(n2687), .B2(n2688), .A(n12545), .ZN(n2686) );
  NAND4_X1 U5031 ( .A1(n2689), .A2(n2690), .A3(n2691), .A4(n2692), .ZN(n2688)
         );
  NAND4_X1 U5032 ( .A1(n2697), .A2(n2698), .A3(n2699), .A4(n2700), .ZN(n2687)
         );
  OAI21_X1 U5033 ( .B1(n4806), .B2(n12541), .A(n2667), .ZN(n4953) );
  OAI21_X1 U5034 ( .B1(n2668), .B2(n2669), .A(n12544), .ZN(n2667) );
  NAND4_X1 U5035 ( .A1(n2670), .A2(n2671), .A3(n2672), .A4(n2673), .ZN(n2669)
         );
  NAND4_X1 U5036 ( .A1(n2678), .A2(n2679), .A3(n2680), .A4(n2681), .ZN(n2668)
         );
  OAI21_X1 U5037 ( .B1(n4805), .B2(n12541), .A(n2648), .ZN(n4954) );
  OAI21_X1 U5038 ( .B1(n2649), .B2(n2650), .A(n12544), .ZN(n2648) );
  NAND4_X1 U5039 ( .A1(n2651), .A2(n2652), .A3(n2653), .A4(n2654), .ZN(n2650)
         );
  NAND4_X1 U5040 ( .A1(n2659), .A2(n2660), .A3(n2661), .A4(n2662), .ZN(n2649)
         );
  OAI21_X1 U5041 ( .B1(n4804), .B2(n12541), .A(n2629), .ZN(n4955) );
  OAI21_X1 U5042 ( .B1(n2630), .B2(n2631), .A(n12545), .ZN(n2629) );
  NAND4_X1 U5043 ( .A1(n2632), .A2(n2633), .A3(n2634), .A4(n2635), .ZN(n2631)
         );
  NAND4_X1 U5044 ( .A1(n2640), .A2(n2641), .A3(n2642), .A4(n2643), .ZN(n2630)
         );
  OAI21_X1 U5045 ( .B1(n4803), .B2(n12541), .A(n2610), .ZN(n4956) );
  OAI21_X1 U5046 ( .B1(n2611), .B2(n2612), .A(n12544), .ZN(n2610) );
  NAND4_X1 U5047 ( .A1(n2613), .A2(n2614), .A3(n2615), .A4(n2616), .ZN(n2612)
         );
  NAND4_X1 U5048 ( .A1(n2621), .A2(n2622), .A3(n2623), .A4(n2624), .ZN(n2611)
         );
  OAI21_X1 U5049 ( .B1(n4797), .B2(n12542), .A(n2591), .ZN(n4957) );
  OAI21_X1 U5050 ( .B1(n2592), .B2(n2593), .A(n12544), .ZN(n2591) );
  NAND4_X1 U5051 ( .A1(n2594), .A2(n2595), .A3(n2596), .A4(n2597), .ZN(n2593)
         );
  NAND4_X1 U5052 ( .A1(n2602), .A2(n2603), .A3(n2604), .A4(n2605), .ZN(n2592)
         );
  OAI21_X1 U5053 ( .B1(n4796), .B2(n12541), .A(n2572), .ZN(n4958) );
  OAI21_X1 U5054 ( .B1(n2573), .B2(n2574), .A(n12545), .ZN(n2572) );
  NAND4_X1 U5055 ( .A1(n2575), .A2(n2576), .A3(n2577), .A4(n2578), .ZN(n2574)
         );
  NAND4_X1 U5056 ( .A1(n2583), .A2(n2584), .A3(n2585), .A4(n2586), .ZN(n2573)
         );
  OAI21_X1 U5057 ( .B1(n4795), .B2(n12541), .A(n2553), .ZN(n4959) );
  OAI21_X1 U5058 ( .B1(n2554), .B2(n2555), .A(n12545), .ZN(n2553) );
  NAND4_X1 U5059 ( .A1(n2556), .A2(n2557), .A3(n2558), .A4(n2559), .ZN(n2555)
         );
  NAND4_X1 U5060 ( .A1(n2564), .A2(n2565), .A3(n2566), .A4(n2567), .ZN(n2554)
         );
  OAI21_X1 U5061 ( .B1(n4794), .B2(n12541), .A(n2534), .ZN(n4960) );
  OAI21_X1 U5062 ( .B1(n2535), .B2(n2536), .A(n12545), .ZN(n2534) );
  NAND4_X1 U5063 ( .A1(n2537), .A2(n2538), .A3(n2539), .A4(n2540), .ZN(n2536)
         );
  NAND4_X1 U5064 ( .A1(n2545), .A2(n2546), .A3(n2547), .A4(n2548), .ZN(n2535)
         );
  OAI21_X1 U5065 ( .B1(n4793), .B2(n12541), .A(n2515), .ZN(n4961) );
  OAI21_X1 U5066 ( .B1(n2516), .B2(n2517), .A(n12546), .ZN(n2515) );
  NAND4_X1 U5067 ( .A1(n2518), .A2(n2519), .A3(n2520), .A4(n2521), .ZN(n2517)
         );
  NAND4_X1 U5068 ( .A1(n2526), .A2(n2527), .A3(n2528), .A4(n2529), .ZN(n2516)
         );
  OAI21_X1 U5069 ( .B1(n4792), .B2(n12541), .A(n2496), .ZN(n4962) );
  OAI21_X1 U5070 ( .B1(n2497), .B2(n2498), .A(n12545), .ZN(n2496) );
  NAND4_X1 U5071 ( .A1(n2499), .A2(n2500), .A3(n2501), .A4(n2502), .ZN(n2498)
         );
  NAND4_X1 U5072 ( .A1(n2507), .A2(n2508), .A3(n2509), .A4(n2510), .ZN(n2497)
         );
  OAI21_X1 U5073 ( .B1(n4791), .B2(n12541), .A(n2477), .ZN(n4963) );
  OAI21_X1 U5074 ( .B1(n2478), .B2(n2479), .A(n12545), .ZN(n2477) );
  NAND4_X1 U5075 ( .A1(n2480), .A2(n2481), .A3(n2482), .A4(n2483), .ZN(n2479)
         );
  NAND4_X1 U5076 ( .A1(n2488), .A2(n2489), .A3(n2490), .A4(n2491), .ZN(n2478)
         );
  OAI21_X1 U5077 ( .B1(n4790), .B2(n12541), .A(n2458), .ZN(n4964) );
  OAI21_X1 U5078 ( .B1(n2459), .B2(n2460), .A(n12547), .ZN(n2458) );
  NAND4_X1 U5079 ( .A1(n2461), .A2(n2462), .A3(n2463), .A4(n2464), .ZN(n2460)
         );
  NAND4_X1 U5080 ( .A1(n2469), .A2(n2470), .A3(n2471), .A4(n2472), .ZN(n2459)
         );
  OAI21_X1 U5081 ( .B1(n4789), .B2(n12540), .A(n2439), .ZN(n4965) );
  OAI21_X1 U5082 ( .B1(n2440), .B2(n2441), .A(n12547), .ZN(n2439) );
  NAND4_X1 U5083 ( .A1(n2442), .A2(n2443), .A3(n2444), .A4(n2445), .ZN(n2441)
         );
  NAND4_X1 U5084 ( .A1(n2450), .A2(n2451), .A3(n2452), .A4(n2453), .ZN(n2440)
         );
  OAI21_X1 U5085 ( .B1(n4788), .B2(n12540), .A(n2420), .ZN(n4966) );
  OAI21_X1 U5086 ( .B1(n2421), .B2(n2422), .A(n12546), .ZN(n2420) );
  NAND4_X1 U5087 ( .A1(n2423), .A2(n2424), .A3(n2425), .A4(n2426), .ZN(n2422)
         );
  NAND4_X1 U5088 ( .A1(n2431), .A2(n2432), .A3(n2433), .A4(n2434), .ZN(n2421)
         );
  OAI21_X1 U5089 ( .B1(n4787), .B2(n12540), .A(n2401), .ZN(n4967) );
  OAI21_X1 U5090 ( .B1(n2402), .B2(n2403), .A(n12546), .ZN(n2401) );
  NAND4_X1 U5091 ( .A1(n2404), .A2(n2405), .A3(n2406), .A4(n2407), .ZN(n2403)
         );
  NAND4_X1 U5092 ( .A1(n2412), .A2(n2413), .A3(n2414), .A4(n2415), .ZN(n2402)
         );
  OAI21_X1 U5093 ( .B1(n4786), .B2(n12540), .A(n2382), .ZN(n4968) );
  OAI21_X1 U5094 ( .B1(n2383), .B2(n2384), .A(n12546), .ZN(n2382) );
  NAND4_X1 U5095 ( .A1(n2385), .A2(n2386), .A3(n2387), .A4(n2388), .ZN(n2384)
         );
  NAND4_X1 U5096 ( .A1(n2393), .A2(n2394), .A3(n2395), .A4(n2396), .ZN(n2383)
         );
  OAI21_X1 U5097 ( .B1(n4785), .B2(n12540), .A(n2363), .ZN(n4969) );
  OAI21_X1 U5098 ( .B1(n2364), .B2(n2365), .A(n12546), .ZN(n2363) );
  NAND4_X1 U5099 ( .A1(n2366), .A2(n2367), .A3(n2368), .A4(n2369), .ZN(n2365)
         );
  NAND4_X1 U5100 ( .A1(n2374), .A2(n2375), .A3(n2376), .A4(n2377), .ZN(n2364)
         );
  OAI21_X1 U5101 ( .B1(n4784), .B2(n12540), .A(n2344), .ZN(n4970) );
  OAI21_X1 U5102 ( .B1(n2345), .B2(n2346), .A(n12547), .ZN(n2344) );
  NAND4_X1 U5103 ( .A1(n2347), .A2(n2348), .A3(n2349), .A4(n2350), .ZN(n2346)
         );
  NAND4_X1 U5104 ( .A1(n2355), .A2(n2356), .A3(n2357), .A4(n2358), .ZN(n2345)
         );
  OAI21_X1 U5105 ( .B1(n4783), .B2(n12540), .A(n2325), .ZN(n4971) );
  OAI21_X1 U5106 ( .B1(n2326), .B2(n2327), .A(n12546), .ZN(n2325) );
  NAND4_X1 U5107 ( .A1(n2328), .A2(n2329), .A3(n2330), .A4(n2331), .ZN(n2327)
         );
  NAND4_X1 U5108 ( .A1(n2336), .A2(n2337), .A3(n2338), .A4(n2339), .ZN(n2326)
         );
  OAI21_X1 U5109 ( .B1(n4782), .B2(n12540), .A(n2306), .ZN(n4972) );
  OAI21_X1 U5110 ( .B1(n2307), .B2(n2308), .A(n12547), .ZN(n2306) );
  NAND4_X1 U5111 ( .A1(n2309), .A2(n2310), .A3(n2311), .A4(n2312), .ZN(n2308)
         );
  NAND4_X1 U5112 ( .A1(n2317), .A2(n2318), .A3(n2319), .A4(n2320), .ZN(n2307)
         );
  OAI21_X1 U5113 ( .B1(n4781), .B2(n12540), .A(n2287), .ZN(n4973) );
  OAI21_X1 U5114 ( .B1(n2288), .B2(n2289), .A(n12547), .ZN(n2287) );
  NAND4_X1 U5115 ( .A1(n2290), .A2(n2291), .A3(n2292), .A4(n2293), .ZN(n2289)
         );
  NAND4_X1 U5116 ( .A1(n2298), .A2(n2299), .A3(n2300), .A4(n2301), .ZN(n2288)
         );
  OAI21_X1 U5117 ( .B1(n4780), .B2(n12540), .A(n2268), .ZN(n4974) );
  OAI21_X1 U5118 ( .B1(n2269), .B2(n2270), .A(n12547), .ZN(n2268) );
  NAND4_X1 U5119 ( .A1(n2271), .A2(n2272), .A3(n2273), .A4(n2274), .ZN(n2270)
         );
  NAND4_X1 U5120 ( .A1(n2279), .A2(n2280), .A3(n2281), .A4(n2282), .ZN(n2269)
         );
  OAI21_X1 U5121 ( .B1(n4779), .B2(n12540), .A(n2249), .ZN(n4975) );
  OAI21_X1 U5122 ( .B1(n2250), .B2(n2251), .A(n12547), .ZN(n2249) );
  NAND4_X1 U5123 ( .A1(n2252), .A2(n2253), .A3(n2254), .A4(n2255), .ZN(n2251)
         );
  NAND4_X1 U5124 ( .A1(n2260), .A2(n2261), .A3(n2262), .A4(n2263), .ZN(n2250)
         );
  OAI21_X1 U5125 ( .B1(n4778), .B2(n12540), .A(n2230), .ZN(n4976) );
  OAI21_X1 U5126 ( .B1(n2231), .B2(n2232), .A(n12548), .ZN(n2230) );
  NAND4_X1 U5127 ( .A1(n2233), .A2(n2234), .A3(n2235), .A4(n2236), .ZN(n2232)
         );
  NAND4_X1 U5128 ( .A1(n2241), .A2(n2242), .A3(n2243), .A4(n2244), .ZN(n2231)
         );
  OAI21_X1 U5129 ( .B1(n4777), .B2(n12539), .A(n2211), .ZN(n4977) );
  OAI21_X1 U5130 ( .B1(n2212), .B2(n2213), .A(n12547), .ZN(n2211) );
  NAND4_X1 U5131 ( .A1(n2214), .A2(n2215), .A3(n2216), .A4(n2217), .ZN(n2213)
         );
  NAND4_X1 U5132 ( .A1(n2222), .A2(n2223), .A3(n2224), .A4(n2225), .ZN(n2212)
         );
  OAI21_X1 U5133 ( .B1(n4776), .B2(n12539), .A(n2192), .ZN(n4978) );
  OAI21_X1 U5134 ( .B1(n2193), .B2(n2194), .A(n12547), .ZN(n2192) );
  NAND4_X1 U5135 ( .A1(n2195), .A2(n2196), .A3(n2197), .A4(n2198), .ZN(n2194)
         );
  NAND4_X1 U5136 ( .A1(n2203), .A2(n2204), .A3(n2205), .A4(n2206), .ZN(n2193)
         );
  OAI21_X1 U5137 ( .B1(n4775), .B2(n12539), .A(n2173), .ZN(n4979) );
  OAI21_X1 U5138 ( .B1(n2174), .B2(n2175), .A(n12548), .ZN(n2173) );
  NAND4_X1 U5139 ( .A1(n2176), .A2(n2177), .A3(n2178), .A4(n2179), .ZN(n2175)
         );
  NAND4_X1 U5140 ( .A1(n2184), .A2(n2185), .A3(n2186), .A4(n2187), .ZN(n2174)
         );
  OAI21_X1 U5141 ( .B1(n4774), .B2(n12539), .A(n2154), .ZN(n4980) );
  OAI21_X1 U5142 ( .B1(n2155), .B2(n2156), .A(n12548), .ZN(n2154) );
  NAND4_X1 U5143 ( .A1(n2157), .A2(n2158), .A3(n2159), .A4(n2160), .ZN(n2156)
         );
  NAND4_X1 U5144 ( .A1(n2165), .A2(n2166), .A3(n2167), .A4(n2168), .ZN(n2155)
         );
  OAI21_X1 U5145 ( .B1(n4773), .B2(n12539), .A(n2135), .ZN(n4981) );
  OAI21_X1 U5146 ( .B1(n2136), .B2(n2137), .A(n12548), .ZN(n2135) );
  NAND4_X1 U5147 ( .A1(n2138), .A2(n2139), .A3(n2140), .A4(n2141), .ZN(n2137)
         );
  NAND4_X1 U5148 ( .A1(n2146), .A2(n2147), .A3(n2148), .A4(n2149), .ZN(n2136)
         );
  OAI21_X1 U5149 ( .B1(n4772), .B2(n12539), .A(n2116), .ZN(n4982) );
  OAI21_X1 U5150 ( .B1(n2117), .B2(n2118), .A(n12548), .ZN(n2116) );
  NAND4_X1 U5151 ( .A1(n2119), .A2(n2120), .A3(n2121), .A4(n2122), .ZN(n2118)
         );
  NAND4_X1 U5152 ( .A1(n2127), .A2(n2128), .A3(n2129), .A4(n2130), .ZN(n2117)
         );
  OAI21_X1 U5153 ( .B1(n4771), .B2(n12539), .A(n2097), .ZN(n4983) );
  OAI21_X1 U5154 ( .B1(n2098), .B2(n2099), .A(n12548), .ZN(n2097) );
  NAND4_X1 U5155 ( .A1(n2100), .A2(n2101), .A3(n2102), .A4(n2103), .ZN(n2099)
         );
  NAND4_X1 U5156 ( .A1(n2108), .A2(n2109), .A3(n2110), .A4(n2111), .ZN(n2098)
         );
  OAI21_X1 U5157 ( .B1(n4770), .B2(n12539), .A(n2078), .ZN(n4984) );
  OAI21_X1 U5158 ( .B1(n2079), .B2(n2080), .A(n12548), .ZN(n2078) );
  NAND4_X1 U5159 ( .A1(n2081), .A2(n2082), .A3(n2083), .A4(n2084), .ZN(n2080)
         );
  NAND4_X1 U5160 ( .A1(n2089), .A2(n2090), .A3(n2091), .A4(n2092), .ZN(n2079)
         );
  OAI21_X1 U5161 ( .B1(n4769), .B2(n12539), .A(n2059), .ZN(n4985) );
  OAI21_X1 U5162 ( .B1(n2060), .B2(n2061), .A(n12549), .ZN(n2059) );
  NAND4_X1 U5163 ( .A1(n2062), .A2(n2063), .A3(n2064), .A4(n2065), .ZN(n2061)
         );
  NAND4_X1 U5164 ( .A1(n2070), .A2(n2071), .A3(n2072), .A4(n2073), .ZN(n2060)
         );
  OAI21_X1 U5165 ( .B1(n4768), .B2(n12539), .A(n2040), .ZN(n4986) );
  OAI21_X1 U5166 ( .B1(n2041), .B2(n2042), .A(n12549), .ZN(n2040) );
  NAND4_X1 U5167 ( .A1(n2043), .A2(n2044), .A3(n2045), .A4(n2046), .ZN(n2042)
         );
  NAND4_X1 U5168 ( .A1(n2051), .A2(n2052), .A3(n2053), .A4(n2054), .ZN(n2041)
         );
  OAI21_X1 U5169 ( .B1(n4767), .B2(n12539), .A(n2021), .ZN(n4987) );
  OAI21_X1 U5170 ( .B1(n2022), .B2(n2023), .A(n12549), .ZN(n2021) );
  NAND4_X1 U5171 ( .A1(n2024), .A2(n2025), .A3(n2026), .A4(n2027), .ZN(n2023)
         );
  NAND4_X1 U5172 ( .A1(n2032), .A2(n2033), .A3(n2034), .A4(n2035), .ZN(n2022)
         );
  OAI21_X1 U5173 ( .B1(n4766), .B2(n12539), .A(n2002), .ZN(n4988) );
  OAI21_X1 U5174 ( .B1(n2003), .B2(n2004), .A(n12549), .ZN(n2002) );
  NAND4_X1 U5175 ( .A1(n2005), .A2(n2006), .A3(n2007), .A4(n2008), .ZN(n2004)
         );
  NAND4_X1 U5176 ( .A1(n2013), .A2(n2014), .A3(n2015), .A4(n2016), .ZN(n2003)
         );
  OAI21_X1 U5177 ( .B1(n4765), .B2(n12541), .A(n1951), .ZN(n4989) );
  OAI21_X1 U5178 ( .B1(n1952), .B2(n1953), .A(n12549), .ZN(n1951) );
  NAND4_X1 U5179 ( .A1(n1954), .A2(n1955), .A3(n1956), .A4(n1957), .ZN(n1953)
         );
  NAND4_X1 U5180 ( .A1(n1978), .A2(n1979), .A3(n1980), .A4(n1981), .ZN(n1952)
         );
  NOR3_X1 U5181 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n13387), .ZN(n4465) );
  NOR3_X1 U5182 ( .A1(n13387), .A2(ADD_RD2[3]), .A3(n13391), .ZN(n4466) );
  NOR2_X1 U5183 ( .A1(n13390), .A2(ADD_RD2[2]), .ZN(n4452) );
  NOR3_X1 U5184 ( .A1(n13387), .A2(ADD_RD2[0]), .A3(n13388), .ZN(n4469) );
  NOR3_X1 U5185 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n13391), .ZN(n4449) );
  NOR3_X1 U5186 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(n4451) );
  NOR3_X1 U5187 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n13388), .ZN(n4457) );
  NOR3_X1 U5188 ( .A1(n13391), .A2(ADD_RD2[4]), .A3(n13388), .ZN(n4458) );
  AOI221_X1 U5189 ( .B1(n12230), .B2(n4642), .C1(n12224), .C2(n4643), .A(n4464), .ZN(n4463) );
  OAI22_X1 U5190 ( .A1(n8577), .A2(n12218), .B1(n8578), .B2(n12212), .ZN(n4464) );
  AOI221_X1 U5191 ( .B1(n12230), .B2(n4646), .C1(n12224), .C2(n4647), .A(n4437), .ZN(n4436) );
  OAI22_X1 U5192 ( .A1(n8560), .A2(n12218), .B1(n8561), .B2(n12212), .ZN(n4437) );
  AOI221_X1 U5193 ( .B1(n12230), .B2(n4652), .C1(n12224), .C2(n4653), .A(n4418), .ZN(n4417) );
  OAI22_X1 U5194 ( .A1(n8543), .A2(n12218), .B1(n8544), .B2(n12212), .ZN(n4418) );
  AOI221_X1 U5195 ( .B1(n12230), .B2(n4654), .C1(n12224), .C2(n4655), .A(n4399), .ZN(n4398) );
  OAI22_X1 U5196 ( .A1(n8526), .A2(n12218), .B1(n8527), .B2(n12212), .ZN(n4399) );
  AOI221_X1 U5197 ( .B1(n12230), .B2(n8599), .C1(n12224), .C2(n8600), .A(n4380), .ZN(n4379) );
  OAI22_X1 U5198 ( .A1(n8509), .A2(n12218), .B1(n8510), .B2(n12212), .ZN(n4380) );
  AOI221_X1 U5199 ( .B1(n12230), .B2(n8603), .C1(n12224), .C2(n8604), .A(n4361), .ZN(n4360) );
  OAI22_X1 U5200 ( .A1(n8492), .A2(n12218), .B1(n8493), .B2(n12212), .ZN(n4361) );
  AOI221_X1 U5201 ( .B1(n12230), .B2(n8611), .C1(n12224), .C2(n8612), .A(n4342), .ZN(n4341) );
  OAI22_X1 U5202 ( .A1(n8475), .A2(n12218), .B1(n8476), .B2(n12212), .ZN(n4342) );
  AOI221_X1 U5203 ( .B1(n12230), .B2(n8617), .C1(n12224), .C2(n8618), .A(n4323), .ZN(n4322) );
  OAI22_X1 U5204 ( .A1(n8458), .A2(n12218), .B1(n8459), .B2(n12212), .ZN(n4323) );
  AOI221_X1 U5205 ( .B1(n12230), .B2(n8619), .C1(n12224), .C2(n8620), .A(n4304), .ZN(n4303) );
  OAI22_X1 U5206 ( .A1(n8441), .A2(n12218), .B1(n8442), .B2(n12212), .ZN(n4304) );
  AOI221_X1 U5207 ( .B1(n12230), .B2(n8621), .C1(n12224), .C2(n8622), .A(n4285), .ZN(n4284) );
  OAI22_X1 U5208 ( .A1(n8424), .A2(n12218), .B1(n8425), .B2(n12212), .ZN(n4285) );
  AOI221_X1 U5209 ( .B1(n12230), .B2(n8623), .C1(n12224), .C2(n8624), .A(n4266), .ZN(n4265) );
  OAI22_X1 U5210 ( .A1(n8407), .A2(n12218), .B1(n8408), .B2(n12212), .ZN(n4266) );
  AOI221_X1 U5211 ( .B1(n12230), .B2(n8625), .C1(n12224), .C2(n8626), .A(n4247), .ZN(n4246) );
  OAI22_X1 U5212 ( .A1(n8390), .A2(n12218), .B1(n8391), .B2(n12212), .ZN(n4247) );
  AOI221_X1 U5213 ( .B1(n12231), .B2(n8627), .C1(n12225), .C2(n8628), .A(n4228), .ZN(n4227) );
  OAI22_X1 U5214 ( .A1(n8373), .A2(n12219), .B1(n8374), .B2(n12213), .ZN(n4228) );
  AOI221_X1 U5215 ( .B1(n12327), .B2(n9999), .C1(n12321), .C2(n9935), .A(n4201), .ZN(n4200) );
  OAI22_X1 U5216 ( .A1(n14305), .A2(n12315), .B1(n13417), .B2(n12309), .ZN(
        n4201) );
  AOI221_X1 U5217 ( .B1(n12231), .B2(n8629), .C1(n12225), .C2(n8630), .A(n4209), .ZN(n4208) );
  OAI22_X1 U5218 ( .A1(n8356), .A2(n12219), .B1(n8357), .B2(n12213), .ZN(n4209) );
  AOI221_X1 U5219 ( .B1(n12327), .B2(n9998), .C1(n12321), .C2(n9934), .A(n4182), .ZN(n4181) );
  OAI22_X1 U5220 ( .A1(n14304), .A2(n12315), .B1(n13416), .B2(n12309), .ZN(
        n4182) );
  AOI221_X1 U5221 ( .B1(n12231), .B2(n8631), .C1(n12225), .C2(n8632), .A(n4190), .ZN(n4189) );
  OAI22_X1 U5222 ( .A1(n8339), .A2(n12219), .B1(n8340), .B2(n12213), .ZN(n4190) );
  AOI221_X1 U5223 ( .B1(n12327), .B2(n9997), .C1(n12321), .C2(n9933), .A(n4163), .ZN(n4162) );
  OAI22_X1 U5224 ( .A1(n14303), .A2(n12315), .B1(n13415), .B2(n12309), .ZN(
        n4163) );
  AOI221_X1 U5225 ( .B1(n12231), .B2(n8633), .C1(n12225), .C2(n8634), .A(n4171), .ZN(n4170) );
  OAI22_X1 U5226 ( .A1(n8322), .A2(n12219), .B1(n8323), .B2(n12213), .ZN(n4171) );
  AOI221_X1 U5227 ( .B1(n12327), .B2(n9996), .C1(n12321), .C2(n9932), .A(n4144), .ZN(n4143) );
  OAI22_X1 U5228 ( .A1(n14302), .A2(n12315), .B1(n13414), .B2(n12309), .ZN(
        n4144) );
  AOI221_X1 U5229 ( .B1(n12231), .B2(n8635), .C1(n12225), .C2(n8636), .A(n4152), .ZN(n4151) );
  OAI22_X1 U5230 ( .A1(n8305), .A2(n12219), .B1(n8306), .B2(n12213), .ZN(n4152) );
  AOI221_X1 U5231 ( .B1(n12327), .B2(n9995), .C1(n12321), .C2(n9931), .A(n4125), .ZN(n4124) );
  OAI22_X1 U5232 ( .A1(n14301), .A2(n12315), .B1(n13413), .B2(n12309), .ZN(
        n4125) );
  AOI221_X1 U5233 ( .B1(n12231), .B2(n8637), .C1(n12225), .C2(n8638), .A(n4133), .ZN(n4132) );
  OAI22_X1 U5234 ( .A1(n8288), .A2(n12219), .B1(n8289), .B2(n12213), .ZN(n4133) );
  AOI221_X1 U5235 ( .B1(n12327), .B2(n9994), .C1(n12321), .C2(n9930), .A(n4106), .ZN(n4105) );
  OAI22_X1 U5236 ( .A1(n14300), .A2(n12315), .B1(n13412), .B2(n12309), .ZN(
        n4106) );
  AOI221_X1 U5237 ( .B1(n12231), .B2(n8639), .C1(n12225), .C2(n8640), .A(n4114), .ZN(n4113) );
  OAI22_X1 U5238 ( .A1(n8271), .A2(n12219), .B1(n8272), .B2(n12213), .ZN(n4114) );
  AOI221_X1 U5239 ( .B1(n12327), .B2(n9993), .C1(n12321), .C2(n9929), .A(n4087), .ZN(n4086) );
  OAI22_X1 U5240 ( .A1(n14299), .A2(n12315), .B1(n13411), .B2(n12309), .ZN(
        n4087) );
  AOI221_X1 U5241 ( .B1(n12231), .B2(n8641), .C1(n12225), .C2(n8642), .A(n4095), .ZN(n4094) );
  OAI22_X1 U5242 ( .A1(n8254), .A2(n12219), .B1(n8255), .B2(n12213), .ZN(n4095) );
  AOI221_X1 U5243 ( .B1(n12327), .B2(n9992), .C1(n12321), .C2(n9928), .A(n4068), .ZN(n4067) );
  OAI22_X1 U5244 ( .A1(n14298), .A2(n12315), .B1(n13410), .B2(n12309), .ZN(
        n4068) );
  AOI221_X1 U5245 ( .B1(n12231), .B2(n8643), .C1(n12225), .C2(n8644), .A(n4076), .ZN(n4075) );
  OAI22_X1 U5246 ( .A1(n8237), .A2(n12219), .B1(n8238), .B2(n12213), .ZN(n4076) );
  AOI221_X1 U5247 ( .B1(n12327), .B2(n9991), .C1(n12321), .C2(n9927), .A(n4049), .ZN(n4048) );
  OAI22_X1 U5248 ( .A1(n14297), .A2(n12315), .B1(n13409), .B2(n12309), .ZN(
        n4049) );
  AOI221_X1 U5249 ( .B1(n12231), .B2(n8645), .C1(n12225), .C2(n8646), .A(n4057), .ZN(n4056) );
  OAI22_X1 U5250 ( .A1(n8220), .A2(n12219), .B1(n8221), .B2(n12213), .ZN(n4057) );
  AOI221_X1 U5251 ( .B1(n12327), .B2(n9990), .C1(n12321), .C2(n9926), .A(n4030), .ZN(n4029) );
  OAI22_X1 U5252 ( .A1(n14296), .A2(n12315), .B1(n13408), .B2(n12309), .ZN(
        n4030) );
  AOI221_X1 U5253 ( .B1(n12231), .B2(n8647), .C1(n12225), .C2(n8648), .A(n4038), .ZN(n4037) );
  OAI22_X1 U5254 ( .A1(n8203), .A2(n12219), .B1(n8204), .B2(n12213), .ZN(n4038) );
  AOI221_X1 U5255 ( .B1(n12327), .B2(n9989), .C1(n12321), .C2(n9925), .A(n4011), .ZN(n4010) );
  OAI22_X1 U5256 ( .A1(n14295), .A2(n12315), .B1(n13407), .B2(n12309), .ZN(
        n4011) );
  AOI221_X1 U5257 ( .B1(n12231), .B2(n8649), .C1(n12225), .C2(n8650), .A(n4019), .ZN(n4018) );
  OAI22_X1 U5258 ( .A1(n8186), .A2(n12219), .B1(n8187), .B2(n12213), .ZN(n4019) );
  AOI221_X1 U5259 ( .B1(n12328), .B2(n9988), .C1(n12322), .C2(n9924), .A(n3992), .ZN(n3991) );
  OAI22_X1 U5260 ( .A1(n14294), .A2(n12316), .B1(n13406), .B2(n12310), .ZN(
        n3992) );
  AOI221_X1 U5261 ( .B1(n12232), .B2(n8651), .C1(n12226), .C2(n8652), .A(n4000), .ZN(n3999) );
  OAI22_X1 U5262 ( .A1(n8169), .A2(n12220), .B1(n8170), .B2(n12214), .ZN(n4000) );
  AOI221_X1 U5263 ( .B1(n12328), .B2(n9987), .C1(n12322), .C2(n9923), .A(n3973), .ZN(n3972) );
  OAI22_X1 U5264 ( .A1(n14293), .A2(n12316), .B1(n13405), .B2(n12310), .ZN(
        n3973) );
  AOI221_X1 U5265 ( .B1(n12232), .B2(n8653), .C1(n12226), .C2(n8654), .A(n3981), .ZN(n3980) );
  OAI22_X1 U5266 ( .A1(n8152), .A2(n12220), .B1(n8153), .B2(n12214), .ZN(n3981) );
  AOI221_X1 U5267 ( .B1(n12328), .B2(n9986), .C1(n12322), .C2(n9922), .A(n3954), .ZN(n3953) );
  OAI22_X1 U5268 ( .A1(n14292), .A2(n12316), .B1(n13404), .B2(n12310), .ZN(
        n3954) );
  AOI221_X1 U5269 ( .B1(n12232), .B2(n8655), .C1(n12226), .C2(n8656), .A(n3962), .ZN(n3961) );
  OAI22_X1 U5270 ( .A1(n8135), .A2(n12220), .B1(n8136), .B2(n12214), .ZN(n3962) );
  AOI221_X1 U5271 ( .B1(n12328), .B2(n9985), .C1(n12322), .C2(n9921), .A(n3935), .ZN(n3934) );
  OAI22_X1 U5272 ( .A1(n14291), .A2(n12316), .B1(n13403), .B2(n12310), .ZN(
        n3935) );
  AOI221_X1 U5273 ( .B1(n12232), .B2(n8657), .C1(n12226), .C2(n8658), .A(n3943), .ZN(n3942) );
  OAI22_X1 U5274 ( .A1(n8118), .A2(n12220), .B1(n8119), .B2(n12214), .ZN(n3943) );
  AOI221_X1 U5275 ( .B1(n12328), .B2(n9984), .C1(n12322), .C2(n9920), .A(n3916), .ZN(n3915) );
  OAI22_X1 U5276 ( .A1(n14290), .A2(n12316), .B1(n13402), .B2(n12310), .ZN(
        n3916) );
  AOI221_X1 U5277 ( .B1(n12232), .B2(n8659), .C1(n12226), .C2(n8660), .A(n3924), .ZN(n3923) );
  OAI22_X1 U5278 ( .A1(n8101), .A2(n12220), .B1(n8102), .B2(n12214), .ZN(n3924) );
  AOI221_X1 U5279 ( .B1(n12328), .B2(n9983), .C1(n12322), .C2(n9919), .A(n3897), .ZN(n3896) );
  OAI22_X1 U5280 ( .A1(n14289), .A2(n12316), .B1(n14322), .B2(n12310), .ZN(
        n3897) );
  AOI221_X1 U5281 ( .B1(n12232), .B2(n8661), .C1(n12226), .C2(n8662), .A(n3905), .ZN(n3904) );
  OAI22_X1 U5282 ( .A1(n8084), .A2(n12220), .B1(n8085), .B2(n12214), .ZN(n3905) );
  AOI221_X1 U5283 ( .B1(n12328), .B2(n9982), .C1(n12322), .C2(n9918), .A(n3878), .ZN(n3877) );
  OAI22_X1 U5284 ( .A1(n14456), .A2(n12316), .B1(n14321), .B2(n12310), .ZN(
        n3878) );
  AOI221_X1 U5285 ( .B1(n12232), .B2(n8663), .C1(n12226), .C2(n8664), .A(n3886), .ZN(n3885) );
  OAI22_X1 U5286 ( .A1(n8067), .A2(n12220), .B1(n8068), .B2(n12214), .ZN(n3886) );
  AOI221_X1 U5287 ( .B1(n12328), .B2(n9981), .C1(n12322), .C2(n9917), .A(n3859), .ZN(n3858) );
  OAI22_X1 U5288 ( .A1(n14455), .A2(n12316), .B1(n14320), .B2(n12310), .ZN(
        n3859) );
  AOI221_X1 U5289 ( .B1(n12232), .B2(n8665), .C1(n12226), .C2(n8666), .A(n3867), .ZN(n3866) );
  OAI22_X1 U5290 ( .A1(n8050), .A2(n12220), .B1(n8051), .B2(n12214), .ZN(n3867) );
  AOI221_X1 U5291 ( .B1(n12328), .B2(n9980), .C1(n12322), .C2(n9916), .A(n3840), .ZN(n3839) );
  OAI22_X1 U5292 ( .A1(n14454), .A2(n12316), .B1(n14319), .B2(n12310), .ZN(
        n3840) );
  AOI221_X1 U5293 ( .B1(n12232), .B2(n8667), .C1(n12226), .C2(n8668), .A(n3848), .ZN(n3847) );
  OAI22_X1 U5294 ( .A1(n8033), .A2(n12220), .B1(n8034), .B2(n12214), .ZN(n3848) );
  AOI221_X1 U5295 ( .B1(n12328), .B2(n9979), .C1(n12322), .C2(n9915), .A(n3821), .ZN(n3820) );
  OAI22_X1 U5296 ( .A1(n14453), .A2(n12316), .B1(n14318), .B2(n12310), .ZN(
        n3821) );
  AOI221_X1 U5297 ( .B1(n12232), .B2(n8669), .C1(n12226), .C2(n8670), .A(n3829), .ZN(n3828) );
  OAI22_X1 U5298 ( .A1(n8016), .A2(n12220), .B1(n8017), .B2(n12214), .ZN(n3829) );
  AOI221_X1 U5299 ( .B1(n12328), .B2(n9978), .C1(n12322), .C2(n9914), .A(n3802), .ZN(n3801) );
  OAI22_X1 U5300 ( .A1(n14452), .A2(n12316), .B1(n14317), .B2(n12310), .ZN(
        n3802) );
  AOI221_X1 U5301 ( .B1(n12232), .B2(n8671), .C1(n12226), .C2(n8672), .A(n3810), .ZN(n3809) );
  OAI22_X1 U5302 ( .A1(n7999), .A2(n12220), .B1(n8000), .B2(n12214), .ZN(n3810) );
  AOI221_X1 U5303 ( .B1(n12328), .B2(n9977), .C1(n12322), .C2(n9913), .A(n3783), .ZN(n3782) );
  OAI22_X1 U5304 ( .A1(n14451), .A2(n12316), .B1(n14316), .B2(n12310), .ZN(
        n3783) );
  AOI221_X1 U5305 ( .B1(n12232), .B2(n8673), .C1(n12226), .C2(n8674), .A(n3791), .ZN(n3790) );
  OAI22_X1 U5306 ( .A1(n7982), .A2(n12220), .B1(n7983), .B2(n12214), .ZN(n3791) );
  AOI221_X1 U5307 ( .B1(n12329), .B2(n9976), .C1(n12323), .C2(n9912), .A(n3764), .ZN(n3763) );
  OAI22_X1 U5308 ( .A1(n14450), .A2(n12317), .B1(n14315), .B2(n12311), .ZN(
        n3764) );
  AOI221_X1 U5309 ( .B1(n12233), .B2(n8675), .C1(n12227), .C2(n8676), .A(n3772), .ZN(n3771) );
  OAI22_X1 U5310 ( .A1(n7965), .A2(n12221), .B1(n7966), .B2(n12215), .ZN(n3772) );
  AOI221_X1 U5311 ( .B1(n12329), .B2(n9975), .C1(n12323), .C2(n9911), .A(n3745), .ZN(n3744) );
  OAI22_X1 U5312 ( .A1(n14449), .A2(n12317), .B1(n14314), .B2(n12311), .ZN(
        n3745) );
  AOI221_X1 U5313 ( .B1(n12233), .B2(n8677), .C1(n12227), .C2(n8678), .A(n3753), .ZN(n3752) );
  OAI22_X1 U5314 ( .A1(n7948), .A2(n12221), .B1(n7949), .B2(n12215), .ZN(n3753) );
  AOI221_X1 U5315 ( .B1(n12329), .B2(n9974), .C1(n12323), .C2(n9910), .A(n3726), .ZN(n3725) );
  OAI22_X1 U5316 ( .A1(n14448), .A2(n12317), .B1(n14313), .B2(n12311), .ZN(
        n3726) );
  AOI221_X1 U5317 ( .B1(n12233), .B2(n8679), .C1(n12227), .C2(n8680), .A(n3734), .ZN(n3733) );
  OAI22_X1 U5318 ( .A1(n7931), .A2(n12221), .B1(n7932), .B2(n12215), .ZN(n3734) );
  AOI221_X1 U5319 ( .B1(n12329), .B2(n9973), .C1(n12323), .C2(n9909), .A(n3707), .ZN(n3706) );
  OAI22_X1 U5320 ( .A1(n14447), .A2(n12317), .B1(n14312), .B2(n12311), .ZN(
        n3707) );
  AOI221_X1 U5321 ( .B1(n12233), .B2(n8681), .C1(n12227), .C2(n8682), .A(n3715), .ZN(n3714) );
  OAI22_X1 U5322 ( .A1(n7914), .A2(n12221), .B1(n7915), .B2(n12215), .ZN(n3715) );
  AOI221_X1 U5323 ( .B1(n12329), .B2(n9972), .C1(n12323), .C2(n9908), .A(n3688), .ZN(n3687) );
  OAI22_X1 U5324 ( .A1(n14446), .A2(n12317), .B1(n14432), .B2(n12311), .ZN(
        n3688) );
  AOI221_X1 U5325 ( .B1(n12233), .B2(n8683), .C1(n12227), .C2(n8684), .A(n3696), .ZN(n3695) );
  OAI22_X1 U5326 ( .A1(n7897), .A2(n12221), .B1(n7898), .B2(n12215), .ZN(n3696) );
  AOI221_X1 U5327 ( .B1(n12329), .B2(n9971), .C1(n12323), .C2(n9907), .A(n3669), .ZN(n3668) );
  OAI22_X1 U5328 ( .A1(n14445), .A2(n12317), .B1(n14431), .B2(n12311), .ZN(
        n3669) );
  AOI221_X1 U5329 ( .B1(n12233), .B2(n8685), .C1(n12227), .C2(n8686), .A(n3677), .ZN(n3676) );
  OAI22_X1 U5330 ( .A1(n7880), .A2(n12221), .B1(n7881), .B2(n12215), .ZN(n3677) );
  AOI221_X1 U5331 ( .B1(n12329), .B2(n9970), .C1(n12323), .C2(n9906), .A(n3650), .ZN(n3649) );
  OAI22_X1 U5332 ( .A1(n14444), .A2(n12317), .B1(n14430), .B2(n12311), .ZN(
        n3650) );
  AOI221_X1 U5333 ( .B1(n12233), .B2(n8687), .C1(n12227), .C2(n8688), .A(n3658), .ZN(n3657) );
  OAI22_X1 U5334 ( .A1(n7863), .A2(n12221), .B1(n7864), .B2(n12215), .ZN(n3658) );
  AOI221_X1 U5335 ( .B1(n12329), .B2(n9969), .C1(n12323), .C2(n9905), .A(n3631), .ZN(n3630) );
  OAI22_X1 U5336 ( .A1(n14443), .A2(n12317), .B1(n14429), .B2(n12311), .ZN(
        n3631) );
  AOI221_X1 U5337 ( .B1(n12233), .B2(n8689), .C1(n12227), .C2(n8690), .A(n3639), .ZN(n3638) );
  OAI22_X1 U5338 ( .A1(n7846), .A2(n12221), .B1(n7847), .B2(n12215), .ZN(n3639) );
  AOI221_X1 U5339 ( .B1(n12329), .B2(n9968), .C1(n12323), .C2(n9904), .A(n3612), .ZN(n3611) );
  OAI22_X1 U5340 ( .A1(n14442), .A2(n12317), .B1(n14428), .B2(n12311), .ZN(
        n3612) );
  AOI221_X1 U5341 ( .B1(n12233), .B2(n8691), .C1(n12227), .C2(n8692), .A(n3620), .ZN(n3619) );
  OAI22_X1 U5342 ( .A1(n7829), .A2(n12221), .B1(n7830), .B2(n12215), .ZN(n3620) );
  AOI221_X1 U5343 ( .B1(n12329), .B2(n9967), .C1(n12323), .C2(n9903), .A(n3593), .ZN(n3592) );
  OAI22_X1 U5344 ( .A1(n14441), .A2(n12317), .B1(n14427), .B2(n12311), .ZN(
        n3593) );
  AOI221_X1 U5345 ( .B1(n12233), .B2(n8693), .C1(n12227), .C2(n8694), .A(n3601), .ZN(n3600) );
  OAI22_X1 U5346 ( .A1(n7812), .A2(n12221), .B1(n7813), .B2(n12215), .ZN(n3601) );
  AOI221_X1 U5347 ( .B1(n12329), .B2(n9966), .C1(n12323), .C2(n9902), .A(n3574), .ZN(n3573) );
  OAI22_X1 U5348 ( .A1(n13401), .A2(n12317), .B1(n14426), .B2(n12311), .ZN(
        n3574) );
  AOI221_X1 U5349 ( .B1(n12233), .B2(n8695), .C1(n12227), .C2(n8696), .A(n3582), .ZN(n3581) );
  OAI22_X1 U5350 ( .A1(n7795), .A2(n12221), .B1(n7796), .B2(n12215), .ZN(n3582) );
  AOI221_X1 U5351 ( .B1(n12329), .B2(n9965), .C1(n12323), .C2(n9901), .A(n3555), .ZN(n3554) );
  OAI22_X1 U5352 ( .A1(n13400), .A2(n12317), .B1(n14425), .B2(n12311), .ZN(
        n3555) );
  AOI221_X1 U5353 ( .B1(n12233), .B2(n4656), .C1(n12227), .C2(n4657), .A(n3563), .ZN(n3562) );
  OAI22_X1 U5354 ( .A1(n7778), .A2(n12221), .B1(n7779), .B2(n12215), .ZN(n3563) );
  AOI221_X1 U5355 ( .B1(n12330), .B2(n9964), .C1(n12324), .C2(n9900), .A(n3536), .ZN(n3535) );
  OAI22_X1 U5356 ( .A1(n13399), .A2(n12318), .B1(n14424), .B2(n12312), .ZN(
        n3536) );
  AOI221_X1 U5357 ( .B1(n12234), .B2(n4658), .C1(n12228), .C2(n4659), .A(n3544), .ZN(n3543) );
  OAI22_X1 U5358 ( .A1(n7761), .A2(n12222), .B1(n7762), .B2(n12216), .ZN(n3544) );
  AOI221_X1 U5359 ( .B1(n12330), .B2(n9963), .C1(n12324), .C2(n9899), .A(n3517), .ZN(n3516) );
  OAI22_X1 U5360 ( .A1(n13398), .A2(n12318), .B1(n14423), .B2(n12312), .ZN(
        n3517) );
  AOI221_X1 U5361 ( .B1(n12234), .B2(n4660), .C1(n12228), .C2(n4661), .A(n3525), .ZN(n3524) );
  OAI22_X1 U5362 ( .A1(n7744), .A2(n12222), .B1(n7745), .B2(n12216), .ZN(n3525) );
  AOI221_X1 U5363 ( .B1(n12330), .B2(n9962), .C1(n12324), .C2(n9898), .A(n3498), .ZN(n3497) );
  OAI22_X1 U5364 ( .A1(n13397), .A2(n12318), .B1(n14422), .B2(n12312), .ZN(
        n3498) );
  AOI221_X1 U5365 ( .B1(n12234), .B2(n4662), .C1(n12228), .C2(n4663), .A(n3506), .ZN(n3505) );
  OAI22_X1 U5366 ( .A1(n7642), .A2(n12222), .B1(n7643), .B2(n12216), .ZN(n3506) );
  AOI221_X1 U5367 ( .B1(n12330), .B2(n9961), .C1(n12324), .C2(n9897), .A(n3479), .ZN(n3478) );
  OAI22_X1 U5368 ( .A1(n13396), .A2(n12318), .B1(n14421), .B2(n12312), .ZN(
        n3479) );
  AOI221_X1 U5369 ( .B1(n12234), .B2(n4664), .C1(n12228), .C2(n4665), .A(n3487), .ZN(n3486) );
  OAI22_X1 U5370 ( .A1(n7625), .A2(n12222), .B1(n7626), .B2(n12216), .ZN(n3487) );
  AOI221_X1 U5371 ( .B1(n12330), .B2(n9960), .C1(n12324), .C2(n9896), .A(n3460), .ZN(n3459) );
  OAI22_X1 U5372 ( .A1(n13395), .A2(n12318), .B1(n14420), .B2(n12312), .ZN(
        n3460) );
  AOI221_X1 U5373 ( .B1(n12234), .B2(n4666), .C1(n12228), .C2(n4667), .A(n3468), .ZN(n3467) );
  OAI22_X1 U5374 ( .A1(n7521), .A2(n12222), .B1(n7522), .B2(n12216), .ZN(n3468) );
  AOI221_X1 U5375 ( .B1(n12330), .B2(n9959), .C1(n12324), .C2(n9895), .A(n3441), .ZN(n3440) );
  OAI22_X1 U5376 ( .A1(n13394), .A2(n12318), .B1(n14419), .B2(n12312), .ZN(
        n3441) );
  AOI221_X1 U5377 ( .B1(n12234), .B2(n4668), .C1(n12228), .C2(n4669), .A(n3449), .ZN(n3448) );
  OAI22_X1 U5378 ( .A1(n7504), .A2(n12222), .B1(n7505), .B2(n12216), .ZN(n3449) );
  AOI221_X1 U5379 ( .B1(n12330), .B2(n9958), .C1(n12324), .C2(n9894), .A(n3422), .ZN(n3421) );
  OAI22_X1 U5380 ( .A1(n13393), .A2(n12318), .B1(n14418), .B2(n12312), .ZN(
        n3422) );
  AOI221_X1 U5381 ( .B1(n12234), .B2(n4670), .C1(n12228), .C2(n4671), .A(n3430), .ZN(n3429) );
  OAI22_X1 U5382 ( .A1(n7402), .A2(n12222), .B1(n7403), .B2(n12216), .ZN(n3430) );
  AOI221_X1 U5383 ( .B1(n12330), .B2(n9957), .C1(n12324), .C2(n9893), .A(n3403), .ZN(n3402) );
  OAI22_X1 U5384 ( .A1(n14440), .A2(n12318), .B1(n14417), .B2(n12312), .ZN(
        n3403) );
  AOI221_X1 U5385 ( .B1(n12234), .B2(n4672), .C1(n12228), .C2(n4673), .A(n3411), .ZN(n3410) );
  OAI22_X1 U5386 ( .A1(n7385), .A2(n12222), .B1(n7386), .B2(n12216), .ZN(n3411) );
  AOI221_X1 U5387 ( .B1(n12330), .B2(n9956), .C1(n12324), .C2(n9892), .A(n3384), .ZN(n3383) );
  OAI22_X1 U5388 ( .A1(n14439), .A2(n12318), .B1(n14416), .B2(n12312), .ZN(
        n3384) );
  AOI221_X1 U5389 ( .B1(n12234), .B2(n4674), .C1(n12228), .C2(n4675), .A(n3392), .ZN(n3391) );
  OAI22_X1 U5390 ( .A1(n7368), .A2(n12222), .B1(n7369), .B2(n12216), .ZN(n3392) );
  AOI221_X1 U5391 ( .B1(n12330), .B2(n9955), .C1(n12324), .C2(n9891), .A(n3365), .ZN(n3364) );
  OAI22_X1 U5392 ( .A1(n14438), .A2(n12318), .B1(n14415), .B2(n12312), .ZN(
        n3365) );
  AOI221_X1 U5393 ( .B1(n12234), .B2(n4676), .C1(n12228), .C2(n4677), .A(n3373), .ZN(n3372) );
  OAI22_X1 U5394 ( .A1(n7269), .A2(n12222), .B1(n7270), .B2(n12216), .ZN(n3373) );
  AOI221_X1 U5395 ( .B1(n12330), .B2(n9954), .C1(n12324), .C2(n9890), .A(n3346), .ZN(n3345) );
  OAI22_X1 U5396 ( .A1(n14437), .A2(n12318), .B1(n14414), .B2(n12312), .ZN(
        n3346) );
  AOI221_X1 U5397 ( .B1(n12234), .B2(n4678), .C1(n12228), .C2(n4679), .A(n3354), .ZN(n3353) );
  OAI22_X1 U5398 ( .A1(n7252), .A2(n12222), .B1(n7253), .B2(n12216), .ZN(n3354) );
  AOI221_X1 U5399 ( .B1(n12330), .B2(n9953), .C1(n12324), .C2(n9889), .A(n3327), .ZN(n3326) );
  OAI22_X1 U5400 ( .A1(n14436), .A2(n12318), .B1(n14413), .B2(n12312), .ZN(
        n3327) );
  AOI221_X1 U5401 ( .B1(n12234), .B2(n4682), .C1(n12228), .C2(n4683), .A(n3335), .ZN(n3334) );
  OAI22_X1 U5402 ( .A1(n7235), .A2(n12222), .B1(n7236), .B2(n12216), .ZN(n3335) );
  AOI221_X1 U5403 ( .B1(n12235), .B2(n4472), .C1(n12229), .C2(n4473), .A(n3316), .ZN(n3315) );
  OAI22_X1 U5404 ( .A1(n7138), .A2(n12223), .B1(n7139), .B2(n12217), .ZN(n3316) );
  AOI221_X1 U5405 ( .B1(n12331), .B2(n9952), .C1(n12325), .C2(n9888), .A(n3308), .ZN(n3307) );
  OAI22_X1 U5406 ( .A1(n14435), .A2(n12319), .B1(n14412), .B2(n12313), .ZN(
        n3308) );
  AOI221_X1 U5407 ( .B1(n12235), .B2(n4474), .C1(n12229), .C2(n4475), .A(n3297), .ZN(n3296) );
  OAI22_X1 U5408 ( .A1(n7121), .A2(n12223), .B1(n7122), .B2(n12217), .ZN(n3297) );
  AOI221_X1 U5409 ( .B1(n12331), .B2(n9951), .C1(n12325), .C2(n9887), .A(n3289), .ZN(n3288) );
  OAI22_X1 U5410 ( .A1(n14434), .A2(n12319), .B1(n14411), .B2(n12313), .ZN(
        n3289) );
  AOI221_X1 U5411 ( .B1(n12235), .B2(n4476), .C1(n12229), .C2(n4477), .A(n3278), .ZN(n3277) );
  OAI22_X1 U5412 ( .A1(n4860), .A2(n12223), .B1(n4861), .B2(n12217), .ZN(n3278) );
  AOI221_X1 U5413 ( .B1(n12331), .B2(n9950), .C1(n12325), .C2(n9886), .A(n3270), .ZN(n3269) );
  OAI22_X1 U5414 ( .A1(n14433), .A2(n12319), .B1(n14410), .B2(n12313), .ZN(
        n3270) );
  AOI221_X1 U5415 ( .B1(n12235), .B2(n4478), .C1(n12229), .C2(n4479), .A(n3245), .ZN(n3242) );
  OAI22_X1 U5416 ( .A1(n4843), .A2(n12223), .B1(n4844), .B2(n12217), .ZN(n3245) );
  AOI221_X1 U5417 ( .B1(n12331), .B2(n9949), .C1(n12325), .C2(n9885), .A(n3221), .ZN(n3218) );
  OAI22_X1 U5418 ( .A1(n13392), .A2(n12319), .B1(n14409), .B2(n12313), .ZN(
        n3221) );
  AOI221_X1 U5419 ( .B1(n12326), .B2(n11766), .C1(n12320), .C2(n9948), .A(
        n4448), .ZN(n4447) );
  OAI22_X1 U5420 ( .A1(n14216), .A2(n12314), .B1(n13430), .B2(n12308), .ZN(
        n4448) );
  AOI221_X1 U5421 ( .B1(n12326), .B2(n11767), .C1(n12320), .C2(n9947), .A(
        n4429), .ZN(n4428) );
  OAI22_X1 U5422 ( .A1(n14328), .A2(n12314), .B1(n13429), .B2(n12308), .ZN(
        n4429) );
  AOI221_X1 U5423 ( .B1(n12326), .B2(n11768), .C1(n12320), .C2(n9946), .A(
        n4410), .ZN(n4409) );
  OAI22_X1 U5424 ( .A1(n14327), .A2(n12314), .B1(n13428), .B2(n12308), .ZN(
        n4410) );
  AOI221_X1 U5425 ( .B1(n12326), .B2(n11769), .C1(n12320), .C2(n9945), .A(
        n4391), .ZN(n4390) );
  OAI22_X1 U5426 ( .A1(n14326), .A2(n12314), .B1(n13427), .B2(n12308), .ZN(
        n4391) );
  AOI221_X1 U5427 ( .B1(n12326), .B2(n11770), .C1(n12320), .C2(n9944), .A(
        n4372), .ZN(n4371) );
  OAI22_X1 U5428 ( .A1(n14325), .A2(n12314), .B1(n13426), .B2(n12308), .ZN(
        n4372) );
  AOI221_X1 U5429 ( .B1(n12326), .B2(n11771), .C1(n12320), .C2(n9943), .A(
        n4353), .ZN(n4352) );
  OAI22_X1 U5430 ( .A1(n14324), .A2(n12314), .B1(n13425), .B2(n12308), .ZN(
        n4353) );
  AOI221_X1 U5431 ( .B1(n12326), .B2(n11772), .C1(n12320), .C2(n9942), .A(
        n4334), .ZN(n4333) );
  OAI22_X1 U5432 ( .A1(n14311), .A2(n12314), .B1(n13424), .B2(n12308), .ZN(
        n4334) );
  AOI221_X1 U5433 ( .B1(n12326), .B2(n11773), .C1(n12320), .C2(n9941), .A(
        n4315), .ZN(n4314) );
  OAI22_X1 U5434 ( .A1(n14310), .A2(n12314), .B1(n13423), .B2(n12308), .ZN(
        n4315) );
  AOI221_X1 U5435 ( .B1(n12326), .B2(n11774), .C1(n12320), .C2(n9940), .A(
        n4296), .ZN(n4295) );
  OAI22_X1 U5436 ( .A1(n14323), .A2(n12314), .B1(n13422), .B2(n12308), .ZN(
        n4296) );
  AOI221_X1 U5437 ( .B1(n12326), .B2(n11775), .C1(n12320), .C2(n9939), .A(
        n4277), .ZN(n4276) );
  OAI22_X1 U5438 ( .A1(n14309), .A2(n12314), .B1(n13421), .B2(n12308), .ZN(
        n4277) );
  AOI221_X1 U5439 ( .B1(n12326), .B2(n11776), .C1(n12320), .C2(n9938), .A(
        n4258), .ZN(n4257) );
  OAI22_X1 U5440 ( .A1(n14308), .A2(n12314), .B1(n13420), .B2(n12308), .ZN(
        n4258) );
  AOI221_X1 U5441 ( .B1(n12326), .B2(n11777), .C1(n12320), .C2(n9937), .A(
        n4239), .ZN(n4238) );
  OAI22_X1 U5442 ( .A1(n14307), .A2(n12314), .B1(n13419), .B2(n12308), .ZN(
        n4239) );
  AOI221_X1 U5443 ( .B1(n12327), .B2(n11778), .C1(n12321), .C2(n9936), .A(
        n4220), .ZN(n4219) );
  OAI22_X1 U5444 ( .A1(n14306), .A2(n12315), .B1(n13418), .B2(n12309), .ZN(
        n4220) );
  AOI221_X1 U5445 ( .B1(n12206), .B2(n4480), .C1(n12200), .C2(n4481), .A(n4467), .ZN(n4462) );
  OAI22_X1 U5446 ( .A1(n8579), .A2(n12194), .B1(n8580), .B2(n12188), .ZN(n4467) );
  AOI221_X1 U5447 ( .B1(n12206), .B2(n4648), .C1(n12200), .C2(n4649), .A(n4438), .ZN(n4435) );
  OAI22_X1 U5448 ( .A1(n8562), .A2(n12194), .B1(n8563), .B2(n12188), .ZN(n4438) );
  AOI221_X1 U5449 ( .B1(n12206), .B2(n4482), .C1(n12200), .C2(n4483), .A(n4419), .ZN(n4416) );
  OAI22_X1 U5450 ( .A1(n8545), .A2(n12194), .B1(n8546), .B2(n12188), .ZN(n4419) );
  AOI221_X1 U5451 ( .B1(n12206), .B2(n4484), .C1(n12200), .C2(n4485), .A(n4400), .ZN(n4397) );
  OAI22_X1 U5452 ( .A1(n8528), .A2(n12194), .B1(n8529), .B2(n12188), .ZN(n4400) );
  AOI221_X1 U5453 ( .B1(n12206), .B2(n7080), .C1(n12200), .C2(n7081), .A(n4381), .ZN(n4378) );
  OAI22_X1 U5454 ( .A1(n8511), .A2(n12194), .B1(n8512), .B2(n12188), .ZN(n4381) );
  AOI221_X1 U5455 ( .B1(n12206), .B2(n8605), .C1(n12200), .C2(n8606), .A(n4362), .ZN(n4359) );
  OAI22_X1 U5456 ( .A1(n8494), .A2(n12194), .B1(n8495), .B2(n12188), .ZN(n4362) );
  AOI221_X1 U5457 ( .B1(n12206), .B2(n8613), .C1(n12200), .C2(n8614), .A(n4343), .ZN(n4340) );
  OAI22_X1 U5458 ( .A1(n8477), .A2(n12194), .B1(n8478), .B2(n12188), .ZN(n4343) );
  AOI221_X1 U5459 ( .B1(n12206), .B2(n7084), .C1(n12200), .C2(n7085), .A(n4324), .ZN(n4321) );
  OAI22_X1 U5460 ( .A1(n8460), .A2(n12194), .B1(n8461), .B2(n12188), .ZN(n4324) );
  AOI221_X1 U5461 ( .B1(n12206), .B2(n7088), .C1(n12200), .C2(n7089), .A(n4305), .ZN(n4302) );
  OAI22_X1 U5462 ( .A1(n8443), .A2(n12194), .B1(n8444), .B2(n12188), .ZN(n4305) );
  AOI221_X1 U5463 ( .B1(n12206), .B2(n7092), .C1(n12200), .C2(n7093), .A(n4286), .ZN(n4283) );
  OAI22_X1 U5464 ( .A1(n8426), .A2(n12194), .B1(n8427), .B2(n12188), .ZN(n4286) );
  AOI221_X1 U5465 ( .B1(n12206), .B2(n7096), .C1(n12200), .C2(n7097), .A(n4267), .ZN(n4264) );
  OAI22_X1 U5466 ( .A1(n8409), .A2(n12194), .B1(n8410), .B2(n12188), .ZN(n4267) );
  AOI221_X1 U5467 ( .B1(n12206), .B2(n7100), .C1(n12200), .C2(n7101), .A(n4248), .ZN(n4245) );
  OAI22_X1 U5468 ( .A1(n8392), .A2(n12194), .B1(n8393), .B2(n12188), .ZN(n4248) );
  AOI221_X1 U5469 ( .B1(n12207), .B2(n7104), .C1(n12201), .C2(n7105), .A(n4229), .ZN(n4226) );
  OAI22_X1 U5470 ( .A1(n8375), .A2(n12195), .B1(n8376), .B2(n12189), .ZN(n4229) );
  AOI221_X1 U5471 ( .B1(n12207), .B2(n7130), .C1(n12201), .C2(n7131), .A(n4210), .ZN(n4207) );
  OAI22_X1 U5472 ( .A1(n8358), .A2(n12195), .B1(n8359), .B2(n12189), .ZN(n4210) );
  AOI221_X1 U5473 ( .B1(n12207), .B2(n7154), .C1(n12201), .C2(n7155), .A(n4191), .ZN(n4188) );
  OAI22_X1 U5474 ( .A1(n8341), .A2(n12195), .B1(n8342), .B2(n12189), .ZN(n4191) );
  AOI221_X1 U5475 ( .B1(n12207), .B2(n7158), .C1(n12201), .C2(n7159), .A(n4172), .ZN(n4169) );
  OAI22_X1 U5476 ( .A1(n8324), .A2(n12195), .B1(n8325), .B2(n12189), .ZN(n4172) );
  AOI221_X1 U5477 ( .B1(n12207), .B2(n7162), .C1(n12201), .C2(n7163), .A(n4153), .ZN(n4150) );
  OAI22_X1 U5478 ( .A1(n8307), .A2(n12195), .B1(n8308), .B2(n12189), .ZN(n4153) );
  AOI221_X1 U5479 ( .B1(n12207), .B2(n7166), .C1(n12201), .C2(n7167), .A(n4134), .ZN(n4131) );
  OAI22_X1 U5480 ( .A1(n8290), .A2(n12195), .B1(n8291), .B2(n12189), .ZN(n4134) );
  AOI221_X1 U5481 ( .B1(n12207), .B2(n7170), .C1(n12201), .C2(n7171), .A(n4115), .ZN(n4112) );
  OAI22_X1 U5482 ( .A1(n8273), .A2(n12195), .B1(n8274), .B2(n12189), .ZN(n4115) );
  AOI221_X1 U5483 ( .B1(n12207), .B2(n7174), .C1(n12201), .C2(n7175), .A(n4096), .ZN(n4093) );
  OAI22_X1 U5484 ( .A1(n8256), .A2(n12195), .B1(n8257), .B2(n12189), .ZN(n4096) );
  AOI221_X1 U5485 ( .B1(n12207), .B2(n7178), .C1(n12201), .C2(n7179), .A(n4077), .ZN(n4074) );
  OAI22_X1 U5486 ( .A1(n8239), .A2(n12195), .B1(n8240), .B2(n12189), .ZN(n4077) );
  AOI221_X1 U5487 ( .B1(n12207), .B2(n7182), .C1(n12201), .C2(n7183), .A(n4058), .ZN(n4055) );
  OAI22_X1 U5488 ( .A1(n8222), .A2(n12195), .B1(n8223), .B2(n12189), .ZN(n4058) );
  AOI221_X1 U5489 ( .B1(n12207), .B2(n7186), .C1(n12201), .C2(n7187), .A(n4039), .ZN(n4036) );
  OAI22_X1 U5490 ( .A1(n8205), .A2(n12195), .B1(n8206), .B2(n12189), .ZN(n4039) );
  AOI221_X1 U5491 ( .B1(n12207), .B2(n7190), .C1(n12201), .C2(n7191), .A(n4020), .ZN(n4017) );
  OAI22_X1 U5492 ( .A1(n8188), .A2(n12195), .B1(n8189), .B2(n12189), .ZN(n4020) );
  AOI221_X1 U5493 ( .B1(n12208), .B2(n7194), .C1(n12202), .C2(n7195), .A(n4001), .ZN(n3998) );
  OAI22_X1 U5494 ( .A1(n8171), .A2(n12196), .B1(n8172), .B2(n12190), .ZN(n4001) );
  AOI221_X1 U5495 ( .B1(n12208), .B2(n7198), .C1(n12202), .C2(n7199), .A(n3982), .ZN(n3979) );
  OAI22_X1 U5496 ( .A1(n8154), .A2(n12196), .B1(n8155), .B2(n12190), .ZN(n3982) );
  AOI221_X1 U5497 ( .B1(n12208), .B2(n7202), .C1(n12202), .C2(n8708), .A(n3963), .ZN(n3960) );
  OAI22_X1 U5498 ( .A1(n8137), .A2(n12196), .B1(n8138), .B2(n12190), .ZN(n3963) );
  AOI221_X1 U5499 ( .B1(n12208), .B2(n7205), .C1(n12202), .C2(n8707), .A(n3944), .ZN(n3941) );
  OAI22_X1 U5500 ( .A1(n8120), .A2(n12196), .B1(n8121), .B2(n12190), .ZN(n3944) );
  AOI221_X1 U5501 ( .B1(n12208), .B2(n7208), .C1(n12202), .C2(n8706), .A(n3925), .ZN(n3922) );
  OAI22_X1 U5502 ( .A1(n8103), .A2(n12196), .B1(n8104), .B2(n12190), .ZN(n3925) );
  AOI221_X1 U5503 ( .B1(n12208), .B2(n7211), .C1(n12202), .C2(n8705), .A(n3906), .ZN(n3903) );
  OAI22_X1 U5504 ( .A1(n8086), .A2(n12196), .B1(n8087), .B2(n12190), .ZN(n3906) );
  AOI221_X1 U5505 ( .B1(n12208), .B2(n7214), .C1(n12202), .C2(n8704), .A(n3887), .ZN(n3884) );
  OAI22_X1 U5506 ( .A1(n8069), .A2(n12196), .B1(n8070), .B2(n12190), .ZN(n3887) );
  AOI221_X1 U5507 ( .B1(n12208), .B2(n7217), .C1(n12202), .C2(n8703), .A(n3868), .ZN(n3865) );
  OAI22_X1 U5508 ( .A1(n8052), .A2(n12196), .B1(n8053), .B2(n12190), .ZN(n3868) );
  AOI221_X1 U5509 ( .B1(n12208), .B2(n7220), .C1(n12202), .C2(n8702), .A(n3849), .ZN(n3846) );
  OAI22_X1 U5510 ( .A1(n8035), .A2(n12196), .B1(n8036), .B2(n12190), .ZN(n3849) );
  AOI221_X1 U5511 ( .B1(n12208), .B2(n7223), .C1(n12202), .C2(n8701), .A(n3830), .ZN(n3827) );
  OAI22_X1 U5512 ( .A1(n8018), .A2(n12196), .B1(n8019), .B2(n12190), .ZN(n3830) );
  AOI221_X1 U5513 ( .B1(n12208), .B2(n7226), .C1(n12202), .C2(n8700), .A(n3811), .ZN(n3808) );
  OAI22_X1 U5514 ( .A1(n8001), .A2(n12196), .B1(n8002), .B2(n12190), .ZN(n3811) );
  AOI221_X1 U5515 ( .B1(n12208), .B2(n7229), .C1(n12202), .C2(n8699), .A(n3792), .ZN(n3789) );
  OAI22_X1 U5516 ( .A1(n7984), .A2(n12196), .B1(n7985), .B2(n12190), .ZN(n3792) );
  AOI221_X1 U5517 ( .B1(n12209), .B2(n7232), .C1(n12203), .C2(n8698), .A(n3773), .ZN(n3770) );
  OAI22_X1 U5518 ( .A1(n7967), .A2(n12197), .B1(n7968), .B2(n12191), .ZN(n3773) );
  AOI221_X1 U5519 ( .B1(n12209), .B2(n7245), .C1(n12203), .C2(n8697), .A(n3754), .ZN(n3751) );
  OAI22_X1 U5520 ( .A1(n7950), .A2(n12197), .B1(n7951), .B2(n12191), .ZN(n3754) );
  AOI221_X1 U5521 ( .B1(n12209), .B2(n7278), .C1(n12203), .C2(n7279), .A(n3735), .ZN(n3732) );
  OAI22_X1 U5522 ( .A1(n7933), .A2(n12197), .B1(n7934), .B2(n12191), .ZN(n3735) );
  AOI221_X1 U5523 ( .B1(n12209), .B2(n7282), .C1(n12203), .C2(n7283), .A(n3716), .ZN(n3713) );
  OAI22_X1 U5524 ( .A1(n7916), .A2(n12197), .B1(n7917), .B2(n12191), .ZN(n3716) );
  AOI221_X1 U5525 ( .B1(n12209), .B2(n7286), .C1(n12203), .C2(n7287), .A(n3697), .ZN(n3694) );
  OAI22_X1 U5526 ( .A1(n7899), .A2(n12197), .B1(n7900), .B2(n12191), .ZN(n3697) );
  AOI221_X1 U5527 ( .B1(n12209), .B2(n7290), .C1(n12203), .C2(n7291), .A(n3678), .ZN(n3675) );
  OAI22_X1 U5528 ( .A1(n7882), .A2(n12197), .B1(n7883), .B2(n12191), .ZN(n3678) );
  AOI221_X1 U5529 ( .B1(n12209), .B2(n7294), .C1(n12203), .C2(n7295), .A(n3659), .ZN(n3656) );
  OAI22_X1 U5530 ( .A1(n7865), .A2(n12197), .B1(n7866), .B2(n12191), .ZN(n3659) );
  AOI221_X1 U5531 ( .B1(n12209), .B2(n7298), .C1(n12203), .C2(n7299), .A(n3640), .ZN(n3637) );
  OAI22_X1 U5532 ( .A1(n7848), .A2(n12197), .B1(n7849), .B2(n12191), .ZN(n3640) );
  AOI221_X1 U5533 ( .B1(n12209), .B2(n7302), .C1(n12203), .C2(n7303), .A(n3621), .ZN(n3618) );
  OAI22_X1 U5534 ( .A1(n7831), .A2(n12197), .B1(n7832), .B2(n12191), .ZN(n3621) );
  AOI221_X1 U5535 ( .B1(n12209), .B2(n7306), .C1(n12203), .C2(n7307), .A(n3602), .ZN(n3599) );
  OAI22_X1 U5536 ( .A1(n7814), .A2(n12197), .B1(n7815), .B2(n12191), .ZN(n3602) );
  AOI221_X1 U5537 ( .B1(n12209), .B2(n7310), .C1(n12203), .C2(n7311), .A(n3583), .ZN(n3580) );
  OAI22_X1 U5538 ( .A1(n7797), .A2(n12197), .B1(n7798), .B2(n12191), .ZN(n3583) );
  AOI221_X1 U5539 ( .B1(n12209), .B2(n7314), .C1(n12203), .C2(n7315), .A(n3564), .ZN(n3561) );
  OAI22_X1 U5540 ( .A1(n7780), .A2(n12197), .B1(n7781), .B2(n12191), .ZN(n3564) );
  AOI221_X1 U5541 ( .B1(n12210), .B2(n7318), .C1(n12204), .C2(n7319), .A(n3545), .ZN(n3542) );
  OAI22_X1 U5542 ( .A1(n7763), .A2(n12198), .B1(n7764), .B2(n12192), .ZN(n3545) );
  AOI221_X1 U5543 ( .B1(n12210), .B2(n7322), .C1(n12204), .C2(n7323), .A(n3526), .ZN(n3523) );
  OAI22_X1 U5544 ( .A1(n7746), .A2(n12198), .B1(n7747), .B2(n12192), .ZN(n3526) );
  AOI221_X1 U5545 ( .B1(n12210), .B2(n4486), .C1(n12204), .C2(n4487), .A(n3507), .ZN(n3504) );
  OAI22_X1 U5546 ( .A1(n7644), .A2(n12198), .B1(n7645), .B2(n12192), .ZN(n3507) );
  AOI221_X1 U5547 ( .B1(n12210), .B2(n4488), .C1(n12204), .C2(n4489), .A(n3488), .ZN(n3485) );
  OAI22_X1 U5548 ( .A1(n7627), .A2(n12198), .B1(n7628), .B2(n12192), .ZN(n3488) );
  AOI221_X1 U5549 ( .B1(n12210), .B2(n4490), .C1(n12204), .C2(n4491), .A(n3469), .ZN(n3466) );
  OAI22_X1 U5550 ( .A1(n7523), .A2(n12198), .B1(n7524), .B2(n12192), .ZN(n3469) );
  AOI221_X1 U5551 ( .B1(n12210), .B2(n4492), .C1(n12204), .C2(n4493), .A(n3450), .ZN(n3447) );
  OAI22_X1 U5552 ( .A1(n7506), .A2(n12198), .B1(n7507), .B2(n12192), .ZN(n3450) );
  AOI221_X1 U5553 ( .B1(n12210), .B2(n4494), .C1(n12204), .C2(n4495), .A(n3431), .ZN(n3428) );
  OAI22_X1 U5554 ( .A1(n7404), .A2(n12198), .B1(n7490), .B2(n12192), .ZN(n3431) );
  AOI221_X1 U5555 ( .B1(n12210), .B2(n4496), .C1(n12204), .C2(n4497), .A(n3412), .ZN(n3409) );
  OAI22_X1 U5556 ( .A1(n7387), .A2(n12198), .B1(n7388), .B2(n12192), .ZN(n3412) );
  AOI221_X1 U5557 ( .B1(n12210), .B2(n4498), .C1(n12204), .C2(n4499), .A(n3393), .ZN(n3390) );
  OAI22_X1 U5558 ( .A1(n7370), .A2(n12198), .B1(n7371), .B2(n12192), .ZN(n3393) );
  AOI221_X1 U5559 ( .B1(n12210), .B2(n4500), .C1(n12204), .C2(n4501), .A(n3374), .ZN(n3371) );
  OAI22_X1 U5560 ( .A1(n7271), .A2(n12198), .B1(n7272), .B2(n12192), .ZN(n3374) );
  AOI221_X1 U5561 ( .B1(n12210), .B2(n4502), .C1(n12204), .C2(n4503), .A(n3355), .ZN(n3352) );
  OAI22_X1 U5562 ( .A1(n7254), .A2(n12198), .B1(n7255), .B2(n12192), .ZN(n3355) );
  AOI221_X1 U5563 ( .B1(n12210), .B2(n4684), .C1(n12204), .C2(n4685), .A(n3336), .ZN(n3333) );
  OAI22_X1 U5564 ( .A1(n7237), .A2(n12198), .B1(n7238), .B2(n12192), .ZN(n3336) );
  AOI221_X1 U5565 ( .B1(n12211), .B2(n4504), .C1(n12205), .C2(n4505), .A(n3317), .ZN(n3314) );
  OAI22_X1 U5566 ( .A1(n7140), .A2(n12199), .B1(n7141), .B2(n12193), .ZN(n3317) );
  AOI221_X1 U5567 ( .B1(n12211), .B2(n4506), .C1(n12205), .C2(n4507), .A(n3298), .ZN(n3295) );
  OAI22_X1 U5568 ( .A1(n7123), .A2(n12199), .B1(n7124), .B2(n12193), .ZN(n3298) );
  AOI221_X1 U5569 ( .B1(n12211), .B2(n4508), .C1(n12205), .C2(n4509), .A(n3279), .ZN(n3276) );
  OAI22_X1 U5570 ( .A1(n7106), .A2(n12199), .B1(n7107), .B2(n12193), .ZN(n3279) );
  AOI221_X1 U5571 ( .B1(n12211), .B2(n4510), .C1(n12205), .C2(n4511), .A(n3250), .ZN(n3241) );
  OAI22_X1 U5572 ( .A1(n4845), .A2(n12199), .B1(n4846), .B2(n12193), .ZN(n3250) );
  INV_X1 U5573 ( .A(ADD_RD2[3]), .ZN(n13388) );
  INV_X1 U5574 ( .A(ADD_RD2[0]), .ZN(n13391) );
  INV_X1 U5575 ( .A(ADD_RD2[4]), .ZN(n13387) );
  AND2_X1 U5576 ( .A1(WR), .A2(ENABLE), .ZN(n1922) );
  NAND2_X1 U5577 ( .A1(DATAIN[63]), .A2(n12132), .ZN(n1841) );
  OAI21_X1 U5578 ( .B1(n8568), .B2(n12339), .A(n4441), .ZN(n4862) );
  OAI21_X1 U5579 ( .B1(n4442), .B2(n4443), .A(n12344), .ZN(n4441) );
  NAND4_X1 U5580 ( .A1(n4460), .A2(n4461), .A3(n4462), .A4(n4463), .ZN(n4442)
         );
  NAND4_X1 U5581 ( .A1(n4444), .A2(n4445), .A3(n4446), .A4(n4447), .ZN(n4443)
         );
  OAI21_X1 U5582 ( .B1(n8551), .B2(n12338), .A(n4422), .ZN(n4863) );
  OAI21_X1 U5583 ( .B1(n4423), .B2(n4424), .A(n12344), .ZN(n4422) );
  NAND4_X1 U5584 ( .A1(n4433), .A2(n4434), .A3(n4435), .A4(n4436), .ZN(n4423)
         );
  NAND4_X1 U5585 ( .A1(n4425), .A2(n4426), .A3(n4427), .A4(n4428), .ZN(n4424)
         );
  OAI21_X1 U5586 ( .B1(n8534), .B2(n12339), .A(n4403), .ZN(n4864) );
  OAI21_X1 U5587 ( .B1(n4404), .B2(n4405), .A(n12344), .ZN(n4403) );
  NAND4_X1 U5588 ( .A1(n4414), .A2(n4415), .A3(n4416), .A4(n4417), .ZN(n4404)
         );
  NAND4_X1 U5589 ( .A1(n4406), .A2(n4407), .A3(n4408), .A4(n4409), .ZN(n4405)
         );
  OAI21_X1 U5590 ( .B1(n8517), .B2(n12338), .A(n4384), .ZN(n4865) );
  OAI21_X1 U5591 ( .B1(n4385), .B2(n4386), .A(n12343), .ZN(n4384) );
  NAND4_X1 U5592 ( .A1(n4395), .A2(n4396), .A3(n4397), .A4(n4398), .ZN(n4385)
         );
  NAND4_X1 U5593 ( .A1(n4387), .A2(n4388), .A3(n4389), .A4(n4390), .ZN(n4386)
         );
  OAI21_X1 U5594 ( .B1(n8500), .B2(n12338), .A(n4365), .ZN(n4866) );
  OAI21_X1 U5595 ( .B1(n4366), .B2(n4367), .A(n12343), .ZN(n4365) );
  NAND4_X1 U5596 ( .A1(n4376), .A2(n4377), .A3(n4378), .A4(n4379), .ZN(n4366)
         );
  NAND4_X1 U5597 ( .A1(n4368), .A2(n4369), .A3(n4370), .A4(n4371), .ZN(n4367)
         );
  OAI21_X1 U5598 ( .B1(n8483), .B2(n12339), .A(n4346), .ZN(n4867) );
  OAI21_X1 U5599 ( .B1(n4347), .B2(n4348), .A(n12343), .ZN(n4346) );
  NAND4_X1 U5600 ( .A1(n4357), .A2(n4358), .A3(n4359), .A4(n4360), .ZN(n4347)
         );
  NAND4_X1 U5601 ( .A1(n4349), .A2(n4350), .A3(n4351), .A4(n4352), .ZN(n4348)
         );
  OAI21_X1 U5602 ( .B1(n8466), .B2(n12339), .A(n4327), .ZN(n4868) );
  OAI21_X1 U5603 ( .B1(n4328), .B2(n4329), .A(n12343), .ZN(n4327) );
  NAND4_X1 U5604 ( .A1(n4338), .A2(n4339), .A3(n4340), .A4(n4341), .ZN(n4328)
         );
  NAND4_X1 U5605 ( .A1(n4330), .A2(n4331), .A3(n4332), .A4(n4333), .ZN(n4329)
         );
  OAI21_X1 U5606 ( .B1(n8449), .B2(n12338), .A(n4308), .ZN(n4869) );
  OAI21_X1 U5607 ( .B1(n4309), .B2(n4310), .A(n12343), .ZN(n4308) );
  NAND4_X1 U5608 ( .A1(n4319), .A2(n4320), .A3(n4321), .A4(n4322), .ZN(n4309)
         );
  NAND4_X1 U5609 ( .A1(n4311), .A2(n4312), .A3(n4313), .A4(n4314), .ZN(n4310)
         );
  OAI21_X1 U5610 ( .B1(n8432), .B2(n12338), .A(n4289), .ZN(n4870) );
  OAI21_X1 U5611 ( .B1(n4290), .B2(n4291), .A(n12342), .ZN(n4289) );
  NAND4_X1 U5612 ( .A1(n4300), .A2(n4301), .A3(n4302), .A4(n4303), .ZN(n4290)
         );
  NAND4_X1 U5613 ( .A1(n4292), .A2(n4293), .A3(n4294), .A4(n4295), .ZN(n4291)
         );
  OAI21_X1 U5614 ( .B1(n8415), .B2(n12338), .A(n4270), .ZN(n4871) );
  OAI21_X1 U5615 ( .B1(n4271), .B2(n4272), .A(n12342), .ZN(n4270) );
  NAND4_X1 U5616 ( .A1(n4281), .A2(n4282), .A3(n4283), .A4(n4284), .ZN(n4271)
         );
  NAND4_X1 U5617 ( .A1(n4273), .A2(n4274), .A3(n4275), .A4(n4276), .ZN(n4272)
         );
  OAI21_X1 U5618 ( .B1(n8398), .B2(n12337), .A(n4251), .ZN(n4872) );
  OAI21_X1 U5619 ( .B1(n4252), .B2(n4253), .A(n12341), .ZN(n4251) );
  NAND4_X1 U5620 ( .A1(n4262), .A2(n4263), .A3(n4264), .A4(n4265), .ZN(n4252)
         );
  NAND4_X1 U5621 ( .A1(n4254), .A2(n4255), .A3(n4256), .A4(n4257), .ZN(n4253)
         );
  OAI21_X1 U5622 ( .B1(n8381), .B2(n12338), .A(n4232), .ZN(n4873) );
  OAI21_X1 U5623 ( .B1(n4233), .B2(n4234), .A(n12341), .ZN(n4232) );
  NAND4_X1 U5624 ( .A1(n4243), .A2(n4244), .A3(n4245), .A4(n4246), .ZN(n4233)
         );
  NAND4_X1 U5625 ( .A1(n4235), .A2(n4236), .A3(n4237), .A4(n4238), .ZN(n4234)
         );
  OAI21_X1 U5626 ( .B1(n8364), .B2(n12338), .A(n4213), .ZN(n4874) );
  OAI21_X1 U5627 ( .B1(n4214), .B2(n4215), .A(n12341), .ZN(n4213) );
  NAND4_X1 U5628 ( .A1(n4224), .A2(n4225), .A3(n4226), .A4(n4227), .ZN(n4214)
         );
  NAND4_X1 U5629 ( .A1(n4216), .A2(n4217), .A3(n4218), .A4(n4219), .ZN(n4215)
         );
  OAI21_X1 U5630 ( .B1(n8347), .B2(n12338), .A(n4194), .ZN(n4875) );
  OAI21_X1 U5631 ( .B1(n4195), .B2(n4196), .A(n12340), .ZN(n4194) );
  NAND4_X1 U5632 ( .A1(n4205), .A2(n4206), .A3(n4207), .A4(n4208), .ZN(n4195)
         );
  NAND4_X1 U5633 ( .A1(n4197), .A2(n4198), .A3(n4199), .A4(n4200), .ZN(n4196)
         );
  OAI21_X1 U5634 ( .B1(n8330), .B2(n12338), .A(n4175), .ZN(n4876) );
  OAI21_X1 U5635 ( .B1(n4176), .B2(n4177), .A(n12342), .ZN(n4175) );
  NAND4_X1 U5636 ( .A1(n4186), .A2(n4187), .A3(n4188), .A4(n4189), .ZN(n4176)
         );
  NAND4_X1 U5637 ( .A1(n4178), .A2(n4179), .A3(n4180), .A4(n4181), .ZN(n4177)
         );
  OAI21_X1 U5638 ( .B1(n8313), .B2(n12338), .A(n4156), .ZN(n4877) );
  OAI21_X1 U5639 ( .B1(n4157), .B2(n4158), .A(n12341), .ZN(n4156) );
  NAND4_X1 U5640 ( .A1(n4167), .A2(n4168), .A3(n4169), .A4(n4170), .ZN(n4157)
         );
  NAND4_X1 U5641 ( .A1(n4159), .A2(n4160), .A3(n4161), .A4(n4162), .ZN(n4158)
         );
  OAI21_X1 U5642 ( .B1(n8296), .B2(n12337), .A(n4137), .ZN(n4878) );
  OAI21_X1 U5643 ( .B1(n4138), .B2(n4139), .A(n12339), .ZN(n4137) );
  NAND4_X1 U5644 ( .A1(n4148), .A2(n4149), .A3(n4150), .A4(n4151), .ZN(n4138)
         );
  NAND4_X1 U5645 ( .A1(n4140), .A2(n4141), .A3(n4142), .A4(n4143), .ZN(n4139)
         );
  OAI21_X1 U5646 ( .B1(n8279), .B2(n12337), .A(n4118), .ZN(n4879) );
  OAI21_X1 U5647 ( .B1(n4119), .B2(n4120), .A(n12341), .ZN(n4118) );
  NAND4_X1 U5648 ( .A1(n4129), .A2(n4130), .A3(n4131), .A4(n4132), .ZN(n4119)
         );
  NAND4_X1 U5649 ( .A1(n4121), .A2(n4122), .A3(n4123), .A4(n4124), .ZN(n4120)
         );
  OAI21_X1 U5650 ( .B1(n8262), .B2(n12338), .A(n4099), .ZN(n4880) );
  OAI21_X1 U5651 ( .B1(n4100), .B2(n4101), .A(n12340), .ZN(n4099) );
  NAND4_X1 U5652 ( .A1(n4110), .A2(n4111), .A3(n4112), .A4(n4113), .ZN(n4100)
         );
  NAND4_X1 U5653 ( .A1(n4102), .A2(n4103), .A3(n4104), .A4(n4105), .ZN(n4101)
         );
  OAI21_X1 U5654 ( .B1(n8245), .B2(n12337), .A(n4080), .ZN(n4881) );
  OAI21_X1 U5655 ( .B1(n4081), .B2(n4082), .A(n12341), .ZN(n4080) );
  NAND4_X1 U5656 ( .A1(n4091), .A2(n4092), .A3(n4093), .A4(n4094), .ZN(n4081)
         );
  NAND4_X1 U5657 ( .A1(n4083), .A2(n4084), .A3(n4085), .A4(n4086), .ZN(n4082)
         );
  OAI21_X1 U5658 ( .B1(n8228), .B2(n12337), .A(n4061), .ZN(n4882) );
  OAI21_X1 U5659 ( .B1(n4062), .B2(n4063), .A(n12339), .ZN(n4061) );
  NAND4_X1 U5660 ( .A1(n4072), .A2(n4073), .A3(n4074), .A4(n4075), .ZN(n4062)
         );
  NAND4_X1 U5661 ( .A1(n4064), .A2(n4065), .A3(n4066), .A4(n4067), .ZN(n4063)
         );
  OAI21_X1 U5662 ( .B1(n8211), .B2(n12337), .A(n4042), .ZN(n4883) );
  OAI21_X1 U5663 ( .B1(n4043), .B2(n4044), .A(n12340), .ZN(n4042) );
  NAND4_X1 U5664 ( .A1(n4053), .A2(n4054), .A3(n4055), .A4(n4056), .ZN(n4043)
         );
  NAND4_X1 U5665 ( .A1(n4045), .A2(n4046), .A3(n4047), .A4(n4048), .ZN(n4044)
         );
  OAI21_X1 U5666 ( .B1(n8194), .B2(n12337), .A(n4023), .ZN(n4884) );
  OAI21_X1 U5667 ( .B1(n4024), .B2(n4025), .A(n12339), .ZN(n4023) );
  NAND4_X1 U5668 ( .A1(n4034), .A2(n4035), .A3(n4036), .A4(n4037), .ZN(n4024)
         );
  NAND4_X1 U5669 ( .A1(n4026), .A2(n4027), .A3(n4028), .A4(n4029), .ZN(n4025)
         );
  OAI21_X1 U5670 ( .B1(n8177), .B2(n12337), .A(n4004), .ZN(n4885) );
  OAI21_X1 U5671 ( .B1(n4005), .B2(n4006), .A(n12340), .ZN(n4004) );
  NAND4_X1 U5672 ( .A1(n4015), .A2(n4016), .A3(n4017), .A4(n4018), .ZN(n4005)
         );
  NAND4_X1 U5673 ( .A1(n4007), .A2(n4008), .A3(n4009), .A4(n4010), .ZN(n4006)
         );
  OAI21_X1 U5674 ( .B1(n8160), .B2(n12337), .A(n3985), .ZN(n4886) );
  OAI21_X1 U5675 ( .B1(n3986), .B2(n3987), .A(n12339), .ZN(n3985) );
  NAND4_X1 U5676 ( .A1(n3996), .A2(n3997), .A3(n3998), .A4(n3999), .ZN(n3986)
         );
  NAND4_X1 U5677 ( .A1(n3988), .A2(n3989), .A3(n3990), .A4(n3991), .ZN(n3987)
         );
  OAI21_X1 U5678 ( .B1(n8143), .B2(n12337), .A(n3966), .ZN(n4887) );
  OAI21_X1 U5679 ( .B1(n3967), .B2(n3968), .A(n12340), .ZN(n3966) );
  NAND4_X1 U5680 ( .A1(n3977), .A2(n3978), .A3(n3979), .A4(n3980), .ZN(n3967)
         );
  NAND4_X1 U5681 ( .A1(n3969), .A2(n3970), .A3(n3971), .A4(n3972), .ZN(n3968)
         );
  OAI21_X1 U5682 ( .B1(n8126), .B2(n12337), .A(n3947), .ZN(n4888) );
  OAI21_X1 U5683 ( .B1(n3948), .B2(n3949), .A(n12340), .ZN(n3947) );
  NAND4_X1 U5684 ( .A1(n3958), .A2(n3959), .A3(n3960), .A4(n3961), .ZN(n3948)
         );
  NAND4_X1 U5685 ( .A1(n3950), .A2(n3951), .A3(n3952), .A4(n3953), .ZN(n3949)
         );
  OAI21_X1 U5686 ( .B1(n8109), .B2(n12336), .A(n3928), .ZN(n4889) );
  OAI21_X1 U5687 ( .B1(n3929), .B2(n3930), .A(n12339), .ZN(n3928) );
  NAND4_X1 U5688 ( .A1(n3939), .A2(n3940), .A3(n3941), .A4(n3942), .ZN(n3929)
         );
  NAND4_X1 U5689 ( .A1(n3931), .A2(n3932), .A3(n3933), .A4(n3934), .ZN(n3930)
         );
  OAI21_X1 U5690 ( .B1(n8092), .B2(n12336), .A(n3909), .ZN(n4890) );
  OAI21_X1 U5691 ( .B1(n3910), .B2(n3911), .A(n12339), .ZN(n3909) );
  NAND4_X1 U5692 ( .A1(n3920), .A2(n3921), .A3(n3922), .A4(n3923), .ZN(n3910)
         );
  NAND4_X1 U5693 ( .A1(n3912), .A2(n3913), .A3(n3914), .A4(n3915), .ZN(n3911)
         );
  OAI21_X1 U5694 ( .B1(n8075), .B2(n12336), .A(n3890), .ZN(n4891) );
  OAI21_X1 U5695 ( .B1(n3891), .B2(n3892), .A(n12340), .ZN(n3890) );
  NAND4_X1 U5696 ( .A1(n3901), .A2(n3902), .A3(n3903), .A4(n3904), .ZN(n3891)
         );
  NAND4_X1 U5697 ( .A1(n3893), .A2(n3894), .A3(n3895), .A4(n3896), .ZN(n3892)
         );
  OAI21_X1 U5698 ( .B1(n8058), .B2(n12336), .A(n3871), .ZN(n4892) );
  OAI21_X1 U5699 ( .B1(n3872), .B2(n3873), .A(n12339), .ZN(n3871) );
  NAND4_X1 U5700 ( .A1(n3882), .A2(n3883), .A3(n3884), .A4(n3885), .ZN(n3872)
         );
  NAND4_X1 U5701 ( .A1(n3874), .A2(n3875), .A3(n3876), .A4(n3877), .ZN(n3873)
         );
  OAI21_X1 U5702 ( .B1(n8041), .B2(n12337), .A(n3852), .ZN(n4893) );
  OAI21_X1 U5703 ( .B1(n3853), .B2(n3854), .A(n12339), .ZN(n3852) );
  NAND4_X1 U5704 ( .A1(n3863), .A2(n3864), .A3(n3865), .A4(n3866), .ZN(n3853)
         );
  NAND4_X1 U5705 ( .A1(n3855), .A2(n3856), .A3(n3857), .A4(n3858), .ZN(n3854)
         );
  OAI21_X1 U5706 ( .B1(n8024), .B2(n12336), .A(n3833), .ZN(n4894) );
  OAI21_X1 U5707 ( .B1(n3834), .B2(n3835), .A(n12340), .ZN(n3833) );
  NAND4_X1 U5708 ( .A1(n3844), .A2(n3845), .A3(n3846), .A4(n3847), .ZN(n3834)
         );
  NAND4_X1 U5709 ( .A1(n3836), .A2(n3837), .A3(n3838), .A4(n3839), .ZN(n3835)
         );
  OAI21_X1 U5710 ( .B1(n8007), .B2(n12336), .A(n3814), .ZN(n4895) );
  OAI21_X1 U5711 ( .B1(n3815), .B2(n3816), .A(n12340), .ZN(n3814) );
  NAND4_X1 U5712 ( .A1(n3825), .A2(n3826), .A3(n3827), .A4(n3828), .ZN(n3815)
         );
  NAND4_X1 U5713 ( .A1(n3817), .A2(n3818), .A3(n3819), .A4(n3820), .ZN(n3816)
         );
  OAI21_X1 U5714 ( .B1(n7990), .B2(n12336), .A(n3795), .ZN(n4896) );
  OAI21_X1 U5715 ( .B1(n3796), .B2(n3797), .A(n12340), .ZN(n3795) );
  NAND4_X1 U5716 ( .A1(n3806), .A2(n3807), .A3(n3808), .A4(n3809), .ZN(n3796)
         );
  NAND4_X1 U5717 ( .A1(n3798), .A2(n3799), .A3(n3800), .A4(n3801), .ZN(n3797)
         );
  OAI21_X1 U5718 ( .B1(n7973), .B2(n12336), .A(n3776), .ZN(n4897) );
  OAI21_X1 U5719 ( .B1(n3777), .B2(n3778), .A(n12341), .ZN(n3776) );
  NAND4_X1 U5720 ( .A1(n3787), .A2(n3788), .A3(n3789), .A4(n3790), .ZN(n3777)
         );
  NAND4_X1 U5721 ( .A1(n3779), .A2(n3780), .A3(n3781), .A4(n3782), .ZN(n3778)
         );
  OAI21_X1 U5722 ( .B1(n7956), .B2(n12336), .A(n3757), .ZN(n4898) );
  OAI21_X1 U5723 ( .B1(n3758), .B2(n3759), .A(n12340), .ZN(n3757) );
  NAND4_X1 U5724 ( .A1(n3768), .A2(n3769), .A3(n3770), .A4(n3771), .ZN(n3758)
         );
  NAND4_X1 U5725 ( .A1(n3760), .A2(n3761), .A3(n3762), .A4(n3763), .ZN(n3759)
         );
  OAI21_X1 U5726 ( .B1(n7939), .B2(n12336), .A(n3738), .ZN(n4899) );
  OAI21_X1 U5727 ( .B1(n3739), .B2(n3740), .A(n12340), .ZN(n3738) );
  NAND4_X1 U5728 ( .A1(n3749), .A2(n3750), .A3(n3751), .A4(n3752), .ZN(n3739)
         );
  NAND4_X1 U5729 ( .A1(n3741), .A2(n3742), .A3(n3743), .A4(n3744), .ZN(n3740)
         );
  OAI21_X1 U5730 ( .B1(n7922), .B2(n12336), .A(n3719), .ZN(n4900) );
  OAI21_X1 U5731 ( .B1(n3720), .B2(n3721), .A(n12342), .ZN(n3719) );
  NAND4_X1 U5732 ( .A1(n3730), .A2(n3731), .A3(n3732), .A4(n3733), .ZN(n3720)
         );
  NAND4_X1 U5733 ( .A1(n3722), .A2(n3723), .A3(n3724), .A4(n3725), .ZN(n3721)
         );
  OAI21_X1 U5734 ( .B1(n7905), .B2(n12335), .A(n3700), .ZN(n4901) );
  OAI21_X1 U5735 ( .B1(n3701), .B2(n3702), .A(n12342), .ZN(n3700) );
  NAND4_X1 U5736 ( .A1(n3711), .A2(n3712), .A3(n3713), .A4(n3714), .ZN(n3701)
         );
  NAND4_X1 U5737 ( .A1(n3703), .A2(n3704), .A3(n3705), .A4(n3706), .ZN(n3702)
         );
  OAI21_X1 U5738 ( .B1(n7888), .B2(n12335), .A(n3681), .ZN(n4902) );
  OAI21_X1 U5739 ( .B1(n3682), .B2(n3683), .A(n12341), .ZN(n3681) );
  NAND4_X1 U5740 ( .A1(n3692), .A2(n3693), .A3(n3694), .A4(n3695), .ZN(n3682)
         );
  NAND4_X1 U5741 ( .A1(n3684), .A2(n3685), .A3(n3686), .A4(n3687), .ZN(n3683)
         );
  OAI21_X1 U5742 ( .B1(n7871), .B2(n12335), .A(n3662), .ZN(n4903) );
  OAI21_X1 U5743 ( .B1(n3663), .B2(n3664), .A(n12341), .ZN(n3662) );
  NAND4_X1 U5744 ( .A1(n3673), .A2(n3674), .A3(n3675), .A4(n3676), .ZN(n3663)
         );
  NAND4_X1 U5745 ( .A1(n3665), .A2(n3666), .A3(n3667), .A4(n3668), .ZN(n3664)
         );
  OAI21_X1 U5746 ( .B1(n7854), .B2(n12335), .A(n3643), .ZN(n4904) );
  OAI21_X1 U5747 ( .B1(n3644), .B2(n3645), .A(n12341), .ZN(n3643) );
  NAND4_X1 U5748 ( .A1(n3654), .A2(n3655), .A3(n3656), .A4(n3657), .ZN(n3644)
         );
  NAND4_X1 U5749 ( .A1(n3646), .A2(n3647), .A3(n3648), .A4(n3649), .ZN(n3645)
         );
  OAI21_X1 U5750 ( .B1(n7837), .B2(n12335), .A(n3624), .ZN(n4905) );
  OAI21_X1 U5751 ( .B1(n3625), .B2(n3626), .A(n12341), .ZN(n3624) );
  NAND4_X1 U5752 ( .A1(n3635), .A2(n3636), .A3(n3637), .A4(n3638), .ZN(n3625)
         );
  NAND4_X1 U5753 ( .A1(n3627), .A2(n3628), .A3(n3629), .A4(n3630), .ZN(n3626)
         );
  OAI21_X1 U5754 ( .B1(n7820), .B2(n12335), .A(n3605), .ZN(n4906) );
  OAI21_X1 U5755 ( .B1(n3606), .B2(n3607), .A(n12342), .ZN(n3605) );
  NAND4_X1 U5756 ( .A1(n3616), .A2(n3617), .A3(n3618), .A4(n3619), .ZN(n3606)
         );
  NAND4_X1 U5757 ( .A1(n3608), .A2(n3609), .A3(n3610), .A4(n3611), .ZN(n3607)
         );
  OAI21_X1 U5758 ( .B1(n7803), .B2(n12335), .A(n3586), .ZN(n4907) );
  OAI21_X1 U5759 ( .B1(n3587), .B2(n3588), .A(n12341), .ZN(n3586) );
  NAND4_X1 U5760 ( .A1(n3597), .A2(n3598), .A3(n3599), .A4(n3600), .ZN(n3587)
         );
  NAND4_X1 U5761 ( .A1(n3589), .A2(n3590), .A3(n3591), .A4(n3592), .ZN(n3588)
         );
  OAI21_X1 U5762 ( .B1(n7786), .B2(n12335), .A(n3567), .ZN(n4908) );
  OAI21_X1 U5763 ( .B1(n3568), .B2(n3569), .A(n12342), .ZN(n3567) );
  NAND4_X1 U5764 ( .A1(n3578), .A2(n3579), .A3(n3580), .A4(n3581), .ZN(n3568)
         );
  NAND4_X1 U5765 ( .A1(n3570), .A2(n3571), .A3(n3572), .A4(n3573), .ZN(n3569)
         );
  OAI21_X1 U5766 ( .B1(n7769), .B2(n12335), .A(n3548), .ZN(n4909) );
  OAI21_X1 U5767 ( .B1(n3549), .B2(n3550), .A(n12342), .ZN(n3548) );
  NAND4_X1 U5768 ( .A1(n3559), .A2(n3560), .A3(n3561), .A4(n3562), .ZN(n3549)
         );
  NAND4_X1 U5769 ( .A1(n3551), .A2(n3552), .A3(n3553), .A4(n3554), .ZN(n3550)
         );
  OAI21_X1 U5770 ( .B1(n7752), .B2(n12335), .A(n3529), .ZN(n4910) );
  OAI21_X1 U5771 ( .B1(n3530), .B2(n3531), .A(n12342), .ZN(n3529) );
  NAND4_X1 U5772 ( .A1(n3540), .A2(n3541), .A3(n3542), .A4(n3543), .ZN(n3530)
         );
  NAND4_X1 U5773 ( .A1(n3532), .A2(n3533), .A3(n3534), .A4(n3535), .ZN(n3531)
         );
  OAI21_X1 U5774 ( .B1(n7650), .B2(n12335), .A(n3510), .ZN(n4911) );
  OAI21_X1 U5775 ( .B1(n3511), .B2(n3512), .A(n12342), .ZN(n3510) );
  NAND4_X1 U5776 ( .A1(n3521), .A2(n3522), .A3(n3523), .A4(n3524), .ZN(n3511)
         );
  NAND4_X1 U5777 ( .A1(n3513), .A2(n3514), .A3(n3515), .A4(n3516), .ZN(n3512)
         );
  OAI21_X1 U5778 ( .B1(n7633), .B2(n12335), .A(n3491), .ZN(n4912) );
  OAI21_X1 U5779 ( .B1(n3492), .B2(n3493), .A(n12343), .ZN(n3491) );
  NAND4_X1 U5780 ( .A1(n3502), .A2(n3503), .A3(n3504), .A4(n3505), .ZN(n3492)
         );
  NAND4_X1 U5781 ( .A1(n3494), .A2(n3495), .A3(n3496), .A4(n3497), .ZN(n3493)
         );
  OAI21_X1 U5782 ( .B1(n7529), .B2(n12334), .A(n3472), .ZN(n4913) );
  OAI21_X1 U5783 ( .B1(n3473), .B2(n3474), .A(n12342), .ZN(n3472) );
  NAND4_X1 U5784 ( .A1(n3483), .A2(n3484), .A3(n3485), .A4(n3486), .ZN(n3473)
         );
  NAND4_X1 U5785 ( .A1(n3475), .A2(n3476), .A3(n3477), .A4(n3478), .ZN(n3474)
         );
  OAI21_X1 U5786 ( .B1(n7512), .B2(n12334), .A(n3453), .ZN(n4914) );
  OAI21_X1 U5787 ( .B1(n3454), .B2(n3455), .A(n12342), .ZN(n3453) );
  NAND4_X1 U5788 ( .A1(n3464), .A2(n3465), .A3(n3466), .A4(n3467), .ZN(n3454)
         );
  NAND4_X1 U5789 ( .A1(n3456), .A2(n3457), .A3(n3458), .A4(n3459), .ZN(n3455)
         );
  OAI21_X1 U5790 ( .B1(n7495), .B2(n12334), .A(n3434), .ZN(n4915) );
  OAI21_X1 U5791 ( .B1(n3435), .B2(n3436), .A(n12343), .ZN(n3434) );
  NAND4_X1 U5792 ( .A1(n3445), .A2(n3446), .A3(n3447), .A4(n3448), .ZN(n3435)
         );
  NAND4_X1 U5793 ( .A1(n3437), .A2(n3438), .A3(n3439), .A4(n3440), .ZN(n3436)
         );
  OAI21_X1 U5794 ( .B1(n7393), .B2(n12334), .A(n3415), .ZN(n4916) );
  OAI21_X1 U5795 ( .B1(n3416), .B2(n3417), .A(n12343), .ZN(n3415) );
  NAND4_X1 U5796 ( .A1(n3426), .A2(n3427), .A3(n3428), .A4(n3429), .ZN(n3416)
         );
  NAND4_X1 U5797 ( .A1(n3418), .A2(n3419), .A3(n3420), .A4(n3421), .ZN(n3417)
         );
  OAI21_X1 U5798 ( .B1(n7376), .B2(n12334), .A(n3396), .ZN(n4917) );
  OAI21_X1 U5799 ( .B1(n3397), .B2(n3398), .A(n12343), .ZN(n3396) );
  NAND4_X1 U5800 ( .A1(n3407), .A2(n3408), .A3(n3409), .A4(n3410), .ZN(n3397)
         );
  NAND4_X1 U5801 ( .A1(n3399), .A2(n3400), .A3(n3401), .A4(n3402), .ZN(n3398)
         );
  OAI21_X1 U5802 ( .B1(n7277), .B2(n12334), .A(n3377), .ZN(n4918) );
  OAI21_X1 U5803 ( .B1(n3378), .B2(n3379), .A(n12343), .ZN(n3377) );
  NAND4_X1 U5804 ( .A1(n3388), .A2(n3389), .A3(n3390), .A4(n3391), .ZN(n3378)
         );
  NAND4_X1 U5805 ( .A1(n3380), .A2(n3381), .A3(n3382), .A4(n3383), .ZN(n3379)
         );
  OAI21_X1 U5806 ( .B1(n7260), .B2(n12334), .A(n3358), .ZN(n4919) );
  OAI21_X1 U5807 ( .B1(n3359), .B2(n3360), .A(n12343), .ZN(n3358) );
  NAND4_X1 U5808 ( .A1(n3369), .A2(n3370), .A3(n3371), .A4(n3372), .ZN(n3359)
         );
  NAND4_X1 U5809 ( .A1(n3361), .A2(n3362), .A3(n3363), .A4(n3364), .ZN(n3360)
         );
  OAI21_X1 U5810 ( .B1(n7243), .B2(n12334), .A(n3339), .ZN(n4920) );
  OAI21_X1 U5811 ( .B1(n3340), .B2(n3341), .A(n12343), .ZN(n3339) );
  NAND4_X1 U5812 ( .A1(n3350), .A2(n3351), .A3(n3352), .A4(n3353), .ZN(n3340)
         );
  NAND4_X1 U5813 ( .A1(n3342), .A2(n3343), .A3(n3344), .A4(n3345), .ZN(n3341)
         );
  OAI21_X1 U5814 ( .B1(n7146), .B2(n12334), .A(n3320), .ZN(n4921) );
  OAI21_X1 U5815 ( .B1(n3321), .B2(n3322), .A(n12344), .ZN(n3320) );
  NAND4_X1 U5816 ( .A1(n3331), .A2(n3332), .A3(n3333), .A4(n3334), .ZN(n3321)
         );
  NAND4_X1 U5817 ( .A1(n3323), .A2(n3324), .A3(n3325), .A4(n3326), .ZN(n3322)
         );
  OAI21_X1 U5818 ( .B1(n7129), .B2(n12334), .A(n3301), .ZN(n4922) );
  OAI21_X1 U5819 ( .B1(n3302), .B2(n3303), .A(n12344), .ZN(n3301) );
  NAND4_X1 U5820 ( .A1(n3304), .A2(n3305), .A3(n3306), .A4(n3307), .ZN(n3303)
         );
  NAND4_X1 U5821 ( .A1(n3312), .A2(n3313), .A3(n3314), .A4(n3315), .ZN(n3302)
         );
  OAI21_X1 U5822 ( .B1(n7112), .B2(n12334), .A(n3282), .ZN(n4923) );
  OAI21_X1 U5823 ( .B1(n3283), .B2(n3284), .A(n12344), .ZN(n3282) );
  NAND4_X1 U5824 ( .A1(n3285), .A2(n3286), .A3(n3287), .A4(n3288), .ZN(n3284)
         );
  NAND4_X1 U5825 ( .A1(n3293), .A2(n3294), .A3(n3295), .A4(n3296), .ZN(n3283)
         );
  OAI21_X1 U5826 ( .B1(n4851), .B2(n12334), .A(n3263), .ZN(n4924) );
  OAI21_X1 U5827 ( .B1(n3264), .B2(n3265), .A(n12344), .ZN(n3263) );
  NAND4_X1 U5828 ( .A1(n3266), .A2(n3267), .A3(n3268), .A4(n3269), .ZN(n3265)
         );
  NAND4_X1 U5829 ( .A1(n3274), .A2(n3275), .A3(n3276), .A4(n3277), .ZN(n3264)
         );
  OAI21_X1 U5830 ( .B1(n4834), .B2(n12336), .A(n3212), .ZN(n4925) );
  OAI21_X1 U5831 ( .B1(n3213), .B2(n3214), .A(n12344), .ZN(n3212) );
  NAND4_X1 U5832 ( .A1(n3215), .A2(n3216), .A3(n3217), .A4(n3218), .ZN(n3214)
         );
  NAND4_X1 U5833 ( .A1(n3239), .A2(n3240), .A3(n3241), .A4(n3242), .ZN(n3213)
         );
  INV_X1 U5834 ( .A(ADD_RD2[1]), .ZN(n13390) );
  INV_X1 U5835 ( .A(ADD_RD2[2]), .ZN(n13389) );
  NAND2_X1 U5836 ( .A1(DATAIN[29]), .A2(n12134), .ZN(n1876) );
  NAND2_X1 U5837 ( .A1(DATAIN[30]), .A2(n12134), .ZN(n1875) );
  NAND2_X1 U5838 ( .A1(DATAIN[31]), .A2(n12134), .ZN(n1874) );
  NAND2_X1 U5839 ( .A1(DATAIN[32]), .A2(n12134), .ZN(n1873) );
  NAND2_X1 U5840 ( .A1(DATAIN[33]), .A2(n12134), .ZN(n1872) );
  NAND2_X1 U5841 ( .A1(DATAIN[34]), .A2(n12134), .ZN(n1871) );
  NAND2_X1 U5842 ( .A1(DATAIN[35]), .A2(n12134), .ZN(n1870) );
  NAND2_X1 U5843 ( .A1(DATAIN[36]), .A2(n12134), .ZN(n1869) );
  NAND2_X1 U5844 ( .A1(DATAIN[37]), .A2(n12134), .ZN(n1868) );
  NAND2_X1 U5845 ( .A1(DATAIN[38]), .A2(n12134), .ZN(n1867) );
  NAND2_X1 U5846 ( .A1(DATAIN[39]), .A2(n12134), .ZN(n1866) );
  NAND2_X1 U5847 ( .A1(DATAIN[40]), .A2(n12133), .ZN(n1865) );
  NAND2_X1 U5848 ( .A1(DATAIN[41]), .A2(n12133), .ZN(n1864) );
  NAND2_X1 U5849 ( .A1(DATAIN[42]), .A2(n12133), .ZN(n1863) );
  NAND2_X1 U5850 ( .A1(DATAIN[43]), .A2(n12133), .ZN(n1862) );
  NAND2_X1 U5851 ( .A1(DATAIN[44]), .A2(n12133), .ZN(n1861) );
  NAND2_X1 U5852 ( .A1(DATAIN[45]), .A2(n12133), .ZN(n1860) );
  NAND2_X1 U5853 ( .A1(DATAIN[55]), .A2(n12132), .ZN(n1850) );
  NAND2_X1 U5854 ( .A1(DATAIN[56]), .A2(n12132), .ZN(n1849) );
  NAND2_X1 U5855 ( .A1(DATAIN[57]), .A2(n12132), .ZN(n1848) );
  NAND2_X1 U5856 ( .A1(DATAIN[58]), .A2(n12132), .ZN(n1847) );
  NAND2_X1 U5857 ( .A1(DATAIN[59]), .A2(n12132), .ZN(n1846) );
  NAND2_X1 U5858 ( .A1(DATAIN[0]), .A2(n12137), .ZN(n1905) );
  NAND2_X1 U5859 ( .A1(DATAIN[1]), .A2(n12137), .ZN(n1904) );
  NAND2_X1 U5860 ( .A1(DATAIN[2]), .A2(n12137), .ZN(n1903) );
  NAND2_X1 U5861 ( .A1(DATAIN[3]), .A2(n12136), .ZN(n1902) );
  NAND2_X1 U5862 ( .A1(DATAIN[4]), .A2(n12137), .ZN(n1901) );
  NAND2_X1 U5863 ( .A1(DATAIN[5]), .A2(n12136), .ZN(n1900) );
  NAND2_X1 U5864 ( .A1(DATAIN[6]), .A2(n12136), .ZN(n1899) );
  NAND2_X1 U5865 ( .A1(DATAIN[7]), .A2(n12136), .ZN(n1898) );
  NAND2_X1 U5866 ( .A1(DATAIN[8]), .A2(n12136), .ZN(n1897) );
  NAND2_X1 U5867 ( .A1(DATAIN[9]), .A2(n12136), .ZN(n1896) );
  NAND2_X1 U5868 ( .A1(DATAIN[10]), .A2(n12136), .ZN(n1895) );
  NAND2_X1 U5869 ( .A1(DATAIN[11]), .A2(n12136), .ZN(n1894) );
  NAND2_X1 U5870 ( .A1(DATAIN[12]), .A2(n12136), .ZN(n1893) );
  NAND2_X1 U5871 ( .A1(DATAIN[13]), .A2(n12136), .ZN(n1892) );
  NAND2_X1 U5872 ( .A1(DATAIN[14]), .A2(n12136), .ZN(n1891) );
  NAND2_X1 U5873 ( .A1(DATAIN[15]), .A2(n12135), .ZN(n1890) );
  NAND2_X1 U5874 ( .A1(DATAIN[16]), .A2(n12136), .ZN(n1889) );
  NAND2_X1 U5875 ( .A1(DATAIN[17]), .A2(n12135), .ZN(n1888) );
  NAND2_X1 U5876 ( .A1(DATAIN[18]), .A2(n12135), .ZN(n1887) );
  NAND2_X1 U5877 ( .A1(DATAIN[19]), .A2(n12135), .ZN(n1886) );
  NAND2_X1 U5878 ( .A1(DATAIN[20]), .A2(n12135), .ZN(n1885) );
  NAND2_X1 U5879 ( .A1(DATAIN[21]), .A2(n12134), .ZN(n1884) );
  NAND2_X1 U5880 ( .A1(DATAIN[22]), .A2(n12135), .ZN(n1883) );
  NAND2_X1 U5881 ( .A1(DATAIN[23]), .A2(n12135), .ZN(n1882) );
  NAND2_X1 U5882 ( .A1(DATAIN[24]), .A2(n12135), .ZN(n1881) );
  NAND2_X1 U5883 ( .A1(DATAIN[25]), .A2(n12135), .ZN(n1880) );
  NAND2_X1 U5884 ( .A1(DATAIN[26]), .A2(n12135), .ZN(n1879) );
  NAND2_X1 U5885 ( .A1(DATAIN[27]), .A2(n12135), .ZN(n1878) );
  NAND2_X1 U5886 ( .A1(DATAIN[28]), .A2(n12135), .ZN(n1877) );
  NAND2_X1 U5887 ( .A1(DATAIN[46]), .A2(n12133), .ZN(n1859) );
  NAND2_X1 U5888 ( .A1(DATAIN[47]), .A2(n12133), .ZN(n1858) );
  NAND2_X1 U5889 ( .A1(DATAIN[48]), .A2(n12133), .ZN(n1857) );
  NAND2_X1 U5890 ( .A1(DATAIN[49]), .A2(n12133), .ZN(n1856) );
  NAND2_X1 U5891 ( .A1(DATAIN[50]), .A2(n12133), .ZN(n1855) );
  NAND2_X1 U5892 ( .A1(DATAIN[51]), .A2(n12133), .ZN(n1854) );
  NAND2_X1 U5893 ( .A1(DATAIN[52]), .A2(n12132), .ZN(n1853) );
  NAND2_X1 U5894 ( .A1(DATAIN[53]), .A2(n12132), .ZN(n1852) );
  NAND2_X1 U5895 ( .A1(DATAIN[54]), .A2(n12132), .ZN(n1851) );
  NAND2_X1 U5896 ( .A1(DATAIN[60]), .A2(n12132), .ZN(n1845) );
  NAND2_X1 U5897 ( .A1(DATAIN[61]), .A2(n12132), .ZN(n1844) );
  NAND2_X1 U5898 ( .A1(DATAIN[62]), .A2(n12132), .ZN(n1843) );
  AND3_X1 U5899 ( .A1(ENABLE), .A2(n12139), .A3(RD1), .ZN(n1950) );
  INV_X1 U5900 ( .A(RESET), .ZN(n14466) );
  OAI22_X1 U5901 ( .A1(n13027), .A2(n13170), .B1(n8574), .B2(n1923), .ZN(n6462) );
  OAI22_X1 U5902 ( .A1(n13027), .A2(n13173), .B1(n8557), .B2(n1923), .ZN(n6463) );
  OAI22_X1 U5903 ( .A1(n13027), .A2(n13176), .B1(n8540), .B2(n1923), .ZN(n6464) );
  OAI22_X1 U5904 ( .A1(n13027), .A2(n13179), .B1(n8523), .B2(n1923), .ZN(n6465) );
  OAI22_X1 U5905 ( .A1(n13026), .A2(n13182), .B1(n8506), .B2(n1923), .ZN(n6466) );
  OAI22_X1 U5906 ( .A1(n13026), .A2(n13185), .B1(n8489), .B2(n1923), .ZN(n6467) );
  OAI22_X1 U5907 ( .A1(n13026), .A2(n13188), .B1(n8472), .B2(n13010), .ZN(
        n6468) );
  OAI22_X1 U5908 ( .A1(n13026), .A2(n13191), .B1(n8455), .B2(n13014), .ZN(
        n6469) );
  OAI22_X1 U5909 ( .A1(n13026), .A2(n13194), .B1(n8438), .B2(n13013), .ZN(
        n6470) );
  OAI22_X1 U5910 ( .A1(n13025), .A2(n13197), .B1(n8421), .B2(n13011), .ZN(
        n6471) );
  OAI22_X1 U5911 ( .A1(n13025), .A2(n13200), .B1(n8404), .B2(n13014), .ZN(
        n6472) );
  OAI22_X1 U5912 ( .A1(n13025), .A2(n13203), .B1(n8387), .B2(n13013), .ZN(
        n6473) );
  OAI22_X1 U5913 ( .A1(n12945), .A2(n13207), .B1(n8372), .B2(n12931), .ZN(
        n6218) );
  OAI22_X1 U5914 ( .A1(n12943), .A2(n13240), .B1(n8185), .B2(n12931), .ZN(
        n6229) );
  OAI22_X1 U5915 ( .A1(n12943), .A2(n13237), .B1(n8202), .B2(n12931), .ZN(
        n6228) );
  OAI22_X1 U5916 ( .A1(n12943), .A2(n13234), .B1(n8219), .B2(n12931), .ZN(
        n6227) );
  OAI22_X1 U5917 ( .A1(n12943), .A2(n13231), .B1(n8236), .B2(n12931), .ZN(
        n6226) );
  OAI22_X1 U5918 ( .A1(n12943), .A2(n13228), .B1(n8253), .B2(n12931), .ZN(
        n6225) );
  OAI22_X1 U5919 ( .A1(n13047), .A2(n13170), .B1(n8572), .B2(n1920), .ZN(n6526) );
  OAI22_X1 U5920 ( .A1(n13047), .A2(n13173), .B1(n8555), .B2(n1920), .ZN(n6527) );
  OAI22_X1 U5921 ( .A1(n13047), .A2(n13176), .B1(n8538), .B2(n1920), .ZN(n6528) );
  OAI22_X1 U5922 ( .A1(n13047), .A2(n13179), .B1(n8521), .B2(n1920), .ZN(n6529) );
  OAI22_X1 U5923 ( .A1(n13046), .A2(n13182), .B1(n8504), .B2(n1920), .ZN(n6530) );
  OAI22_X1 U5924 ( .A1(n13046), .A2(n13185), .B1(n8487), .B2(n1920), .ZN(n6531) );
  OAI22_X1 U5925 ( .A1(n13046), .A2(n13188), .B1(n8470), .B2(n13030), .ZN(
        n6532) );
  OAI22_X1 U5926 ( .A1(n13046), .A2(n13191), .B1(n8453), .B2(n13034), .ZN(
        n6533) );
  OAI22_X1 U5927 ( .A1(n13046), .A2(n13194), .B1(n8436), .B2(n13033), .ZN(
        n6534) );
  OAI22_X1 U5928 ( .A1(n13045), .A2(n13197), .B1(n8419), .B2(n13031), .ZN(
        n6535) );
  OAI22_X1 U5929 ( .A1(n13045), .A2(n13200), .B1(n8402), .B2(n13034), .ZN(
        n6536) );
  OAI22_X1 U5930 ( .A1(n13045), .A2(n13203), .B1(n8385), .B2(n13033), .ZN(
        n6537) );
  OAI22_X1 U5931 ( .A1(n13067), .A2(n13170), .B1(n8571), .B2(n1918), .ZN(n6590) );
  OAI22_X1 U5932 ( .A1(n13067), .A2(n13176), .B1(n8537), .B2(n1918), .ZN(n6592) );
  OAI22_X1 U5933 ( .A1(n13067), .A2(n13179), .B1(n8520), .B2(n1918), .ZN(n6593) );
  OAI22_X1 U5934 ( .A1(n13066), .A2(n13182), .B1(n8503), .B2(n1918), .ZN(n6594) );
  OAI22_X1 U5935 ( .A1(n13066), .A2(n13185), .B1(n8486), .B2(n1918), .ZN(n6595) );
  OAI22_X1 U5936 ( .A1(n13066), .A2(n13188), .B1(n8469), .B2(n1918), .ZN(n6596) );
  OAI22_X1 U5937 ( .A1(n13066), .A2(n13191), .B1(n8452), .B2(n13050), .ZN(
        n6597) );
  OAI22_X1 U5938 ( .A1(n13066), .A2(n13194), .B1(n8435), .B2(n13054), .ZN(
        n6598) );
  OAI22_X1 U5939 ( .A1(n13065), .A2(n13197), .B1(n8418), .B2(n13053), .ZN(
        n6599) );
  OAI22_X1 U5940 ( .A1(n13065), .A2(n13200), .B1(n8401), .B2(n13051), .ZN(
        n6600) );
  OAI22_X1 U5941 ( .A1(n13065), .A2(n13203), .B1(n8384), .B2(n13054), .ZN(
        n6601) );
  OAI22_X1 U5942 ( .A1(n13067), .A2(n13173), .B1(n8554), .B2(n13053), .ZN(
        n6591) );
  OAI21_X1 U5943 ( .B1(n1909), .B2(n1924), .A(n12139), .ZN(n1925) );
  OAI21_X1 U5944 ( .B1(n1907), .B2(n1924), .A(n12139), .ZN(n1923) );
  OAI21_X1 U5945 ( .B1(n1915), .B2(n1924), .A(n12138), .ZN(n1928) );
  OAI22_X1 U5946 ( .A1(n12945), .A2(n13204), .B1(n8389), .B2(n1928), .ZN(n6217) );
  OAI22_X1 U5947 ( .A1(n12945), .A2(n13201), .B1(n8406), .B2(n1928), .ZN(n6216) );
  OAI22_X1 U5948 ( .A1(n12945), .A2(n13198), .B1(n8423), .B2(n1928), .ZN(n6215) );
  OAI22_X1 U5949 ( .A1(n12946), .A2(n13195), .B1(n8440), .B2(n1928), .ZN(n6214) );
  OAI22_X1 U5950 ( .A1(n12946), .A2(n13192), .B1(n8457), .B2(n1928), .ZN(n6213) );
  OAI22_X1 U5951 ( .A1(n12946), .A2(n13189), .B1(n8474), .B2(n1928), .ZN(n6212) );
  AND2_X1 U5952 ( .A1(n3194), .A2(n3204), .ZN(n1987) );
  AND2_X1 U5953 ( .A1(n3191), .A2(n3204), .ZN(n1982) );
  NAND2_X1 U5954 ( .A1(n3193), .A2(n3204), .ZN(n1991) );
  NAND2_X1 U5955 ( .A1(n3189), .A2(n3204), .ZN(n1986) );
  NAND3_X2 U5956 ( .A1(ADD_WR[3]), .A2(n1922), .A3(ADD_WR[4]), .ZN(n1942) );
  OAI22_X1 U5957 ( .A1(n12867), .A2(n13171), .B1(n8578), .B2(n1932), .ZN(n5950) );
  OAI22_X1 U5958 ( .A1(n12867), .A2(n13174), .B1(n8561), .B2(n1932), .ZN(n5951) );
  OAI22_X1 U5959 ( .A1(n12867), .A2(n13177), .B1(n8544), .B2(n1932), .ZN(n5952) );
  OAI22_X1 U5960 ( .A1(n12867), .A2(n13180), .B1(n8527), .B2(n1932), .ZN(n5953) );
  OAI22_X1 U5961 ( .A1(n12866), .A2(n13183), .B1(n8510), .B2(n1932), .ZN(n5954) );
  OAI22_X1 U5962 ( .A1(n12866), .A2(n13186), .B1(n8493), .B2(n1932), .ZN(n5955) );
  OAI22_X1 U5963 ( .A1(n12866), .A2(n13189), .B1(n8476), .B2(n12850), .ZN(
        n5956) );
  OAI22_X1 U5964 ( .A1(n12866), .A2(n13192), .B1(n8459), .B2(n12854), .ZN(
        n5957) );
  OAI22_X1 U5965 ( .A1(n12866), .A2(n13195), .B1(n8442), .B2(n12853), .ZN(
        n5958) );
  OAI22_X1 U5966 ( .A1(n12865), .A2(n13198), .B1(n8425), .B2(n12851), .ZN(
        n5959) );
  OAI22_X1 U5967 ( .A1(n12865), .A2(n13201), .B1(n8408), .B2(n12854), .ZN(
        n5960) );
  OAI22_X1 U5968 ( .A1(n12865), .A2(n13204), .B1(n8391), .B2(n12853), .ZN(
        n5961) );
  OAI21_X1 U5969 ( .B1(n1911), .B2(n1933), .A(n12138), .ZN(n1935) );
  OAI21_X1 U5970 ( .B1(n1913), .B2(n1933), .A(n12138), .ZN(n1936) );
  OAI21_X1 U5971 ( .B1(n1919), .B2(n1933), .A(n12138), .ZN(n1939) );
  OAI21_X1 U5972 ( .B1(n1921), .B2(n1933), .A(n12138), .ZN(n1940) );
  OAI21_X1 U5973 ( .B1(n1909), .B2(n1933), .A(n12138), .ZN(n1934) );
  OAI21_X1 U5974 ( .B1(n1915), .B2(n1933), .A(n12138), .ZN(n1937) );
  OAI21_X1 U5975 ( .B1(n1917), .B2(n1933), .A(n12138), .ZN(n1938) );
  OAI21_X1 U5976 ( .B1(n1907), .B2(n1933), .A(n12138), .ZN(n1932) );
  OAI22_X1 U5977 ( .A1(n13127), .A2(n13170), .B1(n8570), .B2(n1912), .ZN(n6782) );
  OAI22_X1 U5978 ( .A1(n13127), .A2(n13173), .B1(n8553), .B2(n1912), .ZN(n6783) );
  OAI22_X1 U5979 ( .A1(n13127), .A2(n13176), .B1(n8536), .B2(n1912), .ZN(n6784) );
  OAI22_X1 U5980 ( .A1(n13127), .A2(n13179), .B1(n8519), .B2(n1912), .ZN(n6785) );
  OAI22_X1 U5981 ( .A1(n13126), .A2(n13182), .B1(n8502), .B2(n1912), .ZN(n6786) );
  OAI22_X1 U5982 ( .A1(n13126), .A2(n13185), .B1(n8485), .B2(n1912), .ZN(n6787) );
  OAI22_X1 U5983 ( .A1(n13126), .A2(n13188), .B1(n8468), .B2(n1912), .ZN(n6788) );
  OAI22_X1 U5984 ( .A1(n13126), .A2(n13191), .B1(n8451), .B2(n1912), .ZN(n6789) );
  OAI22_X1 U5985 ( .A1(n13126), .A2(n13194), .B1(n8434), .B2(n13110), .ZN(
        n6790) );
  OAI22_X1 U5986 ( .A1(n13125), .A2(n13197), .B1(n8417), .B2(n13111), .ZN(
        n6791) );
  OAI22_X1 U5987 ( .A1(n13125), .A2(n13200), .B1(n8400), .B2(n13114), .ZN(
        n6792) );
  OAI22_X1 U5988 ( .A1(n13125), .A2(n13203), .B1(n8383), .B2(n13113), .ZN(
        n6793) );
  OAI21_X1 U5989 ( .B1(n1906), .B2(n1907), .A(n12137), .ZN(n1842) );
  OAI21_X1 U5990 ( .B1(n1906), .B2(n1909), .A(n12139), .ZN(n1908) );
  OAI21_X1 U5991 ( .B1(n1906), .B2(n1911), .A(n12139), .ZN(n1910) );
  OAI21_X1 U5992 ( .B1(n1906), .B2(n1915), .A(n12139), .ZN(n1914) );
  OAI21_X1 U5993 ( .B1(n1906), .B2(n1917), .A(n12139), .ZN(n1916) );
  OAI21_X1 U5994 ( .B1(n1906), .B2(n1919), .A(n12139), .ZN(n1918) );
  OAI21_X1 U5995 ( .B1(n1906), .B2(n1921), .A(n12139), .ZN(n1920) );
  OAI21_X1 U5996 ( .B1(n1906), .B2(n1913), .A(n12139), .ZN(n1912) );
  INV_X1 U5997 ( .A(ADD_WR[4]), .ZN(n13382) );
  NAND3_X2 U5998 ( .A1(n1922), .A2(n13382), .A3(ADD_WR[3]), .ZN(n1924) );
  CLKBUF_X1 U5999 ( .A(n14466), .Z(n12129) );
  CLKBUF_X1 U6000 ( .A(n14466), .Z(n12130) );
  CLKBUF_X1 U6001 ( .A(n14466), .Z(n12131) );
  CLKBUF_X1 U6002 ( .A(n3262), .Z(n12145) );
  CLKBUF_X1 U6003 ( .A(n3261), .Z(n12151) );
  CLKBUF_X1 U6004 ( .A(n3259), .Z(n12157) );
  CLKBUF_X1 U6005 ( .A(n3258), .Z(n12163) );
  CLKBUF_X1 U6006 ( .A(n3257), .Z(n12169) );
  CLKBUF_X1 U6007 ( .A(n3256), .Z(n12175) );
  CLKBUF_X1 U6008 ( .A(n3254), .Z(n12181) );
  CLKBUF_X1 U6009 ( .A(n3253), .Z(n12187) );
  CLKBUF_X1 U6010 ( .A(n3252), .Z(n12193) );
  CLKBUF_X1 U6011 ( .A(n3251), .Z(n12199) );
  CLKBUF_X1 U6012 ( .A(n3249), .Z(n12205) );
  CLKBUF_X1 U6013 ( .A(n3248), .Z(n12211) );
  CLKBUF_X1 U6014 ( .A(n3247), .Z(n12217) );
  CLKBUF_X1 U6015 ( .A(n3246), .Z(n12223) );
  CLKBUF_X1 U6016 ( .A(n3244), .Z(n12229) );
  CLKBUF_X1 U6017 ( .A(n3243), .Z(n12235) );
  CLKBUF_X1 U6018 ( .A(n3238), .Z(n12241) );
  CLKBUF_X1 U6019 ( .A(n3237), .Z(n12247) );
  CLKBUF_X1 U6020 ( .A(n3235), .Z(n12253) );
  CLKBUF_X1 U6021 ( .A(n3234), .Z(n12259) );
  CLKBUF_X1 U6022 ( .A(n3233), .Z(n12265) );
  CLKBUF_X1 U6023 ( .A(n3232), .Z(n12271) );
  CLKBUF_X1 U6024 ( .A(n3230), .Z(n12277) );
  CLKBUF_X1 U6025 ( .A(n3229), .Z(n12283) );
  CLKBUF_X1 U6026 ( .A(n3228), .Z(n12289) );
  CLKBUF_X1 U6027 ( .A(n3227), .Z(n12295) );
  CLKBUF_X1 U6028 ( .A(n3225), .Z(n12301) );
  CLKBUF_X1 U6029 ( .A(n3224), .Z(n12307) );
  CLKBUF_X1 U6030 ( .A(n3223), .Z(n12313) );
  CLKBUF_X1 U6031 ( .A(n3222), .Z(n12319) );
  CLKBUF_X1 U6032 ( .A(n3220), .Z(n12325) );
  CLKBUF_X1 U6033 ( .A(n3219), .Z(n12331) );
  CLKBUF_X1 U6034 ( .A(n12333), .Z(n12344) );
  CLKBUF_X1 U6035 ( .A(n2001), .Z(n12350) );
  CLKBUF_X1 U6036 ( .A(n2000), .Z(n12356) );
  CLKBUF_X1 U6037 ( .A(n1998), .Z(n12362) );
  CLKBUF_X1 U6038 ( .A(n1997), .Z(n12368) );
  CLKBUF_X1 U6039 ( .A(n1996), .Z(n12374) );
  CLKBUF_X1 U6040 ( .A(n1995), .Z(n12380) );
  CLKBUF_X1 U6041 ( .A(n1993), .Z(n12386) );
  CLKBUF_X1 U6042 ( .A(n1992), .Z(n12392) );
  CLKBUF_X1 U6043 ( .A(n1991), .Z(n12398) );
  CLKBUF_X1 U6044 ( .A(n1990), .Z(n12404) );
  CLKBUF_X1 U6045 ( .A(n1988), .Z(n12410) );
  CLKBUF_X1 U6046 ( .A(n1987), .Z(n12416) );
  CLKBUF_X1 U6047 ( .A(n1986), .Z(n12422) );
  CLKBUF_X1 U6048 ( .A(n1985), .Z(n12428) );
  CLKBUF_X1 U6049 ( .A(n1983), .Z(n12434) );
  CLKBUF_X1 U6050 ( .A(n1982), .Z(n12440) );
  CLKBUF_X1 U6051 ( .A(n1977), .Z(n12446) );
  CLKBUF_X1 U6052 ( .A(n1976), .Z(n12452) );
  CLKBUF_X1 U6053 ( .A(n1974), .Z(n12458) );
  CLKBUF_X1 U6054 ( .A(n1973), .Z(n12464) );
  CLKBUF_X1 U6055 ( .A(n1972), .Z(n12470) );
  CLKBUF_X1 U6056 ( .A(n1971), .Z(n12476) );
  CLKBUF_X1 U6057 ( .A(n1969), .Z(n12482) );
  CLKBUF_X1 U6058 ( .A(n1968), .Z(n12488) );
  CLKBUF_X1 U6059 ( .A(n1967), .Z(n12494) );
  CLKBUF_X1 U6060 ( .A(n1966), .Z(n12500) );
  CLKBUF_X1 U6061 ( .A(n1964), .Z(n12506) );
  CLKBUF_X1 U6062 ( .A(n1963), .Z(n12512) );
  CLKBUF_X1 U6063 ( .A(n1962), .Z(n12518) );
  CLKBUF_X1 U6064 ( .A(n1961), .Z(n12524) );
  CLKBUF_X1 U6065 ( .A(n1959), .Z(n12530) );
  CLKBUF_X1 U6066 ( .A(n1958), .Z(n12536) );
  CLKBUF_X1 U6067 ( .A(n12538), .Z(n12549) );
  INV_X1 U6068 ( .A(n12573), .ZN(n12556) );
endmodule


module MUX21_generic_N5 ( A, B, sel, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input sel;
  wire   n7, n8, n9, n10, n11, n22;

  INV_X1 U1 ( .A(n11), .ZN(Y[0]) );
  AOI22_X1 U2 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n22), .ZN(n11) );
  INV_X1 U3 ( .A(n9), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n22), .ZN(n9) );
  INV_X1 U5 ( .A(n10), .ZN(Y[1]) );
  AOI22_X1 U6 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n22), .ZN(n10) );
  INV_X1 U7 ( .A(n8), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n22), .ZN(n8) );
  INV_X1 U9 ( .A(sel), .ZN(n22) );
  INV_X1 U10 ( .A(n7), .ZN(Y[4]) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[4]), .B1(B[4]), .B2(n22), .ZN(n7) );
endmodule


module address_conversion_M8_N4_N_bit64_F3_DW01_addsub_0 ( A, B, CI, ADD_SUB, 
        SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  FA_X1 U1_4 ( .A(A[4]), .B(B_AS[4]), .CI(carry[4]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA_X1 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA_X1 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA_X1 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0])
         );
  XOR2_X1 U1 ( .A(B[4]), .B(carry[0]), .Z(B_AS[4]) );
  XOR2_X1 U2 ( .A(B[3]), .B(carry[0]), .Z(B_AS[3]) );
  XOR2_X1 U3 ( .A(B[2]), .B(carry[0]), .Z(B_AS[2]) );
  XOR2_X1 U4 ( .A(B[1]), .B(carry[0]), .Z(B_AS[1]) );
  XOR2_X1 U5 ( .A(B[0]), .B(carry[0]), .Z(B_AS[0]) );
endmodule


module address_conversion_M8_N4_N_bit64_F3_DW01_addsub_1 ( A, B, CI, ADD_SUB, 
        SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  FA_X1 U1_4 ( .A(A[4]), .B(B_AS[4]), .CI(carry[4]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA_X1 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA_X1 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA_X1 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0])
         );
  XOR2_X1 U1 ( .A(B[4]), .B(carry[0]), .Z(B_AS[4]) );
  XOR2_X1 U2 ( .A(B[3]), .B(carry[0]), .Z(B_AS[3]) );
  XOR2_X1 U3 ( .A(B[2]), .B(carry[0]), .Z(B_AS[2]) );
  XOR2_X1 U4 ( .A(B[1]), .B(carry[0]), .Z(B_AS[1]) );
  XOR2_X1 U5 ( .A(B[0]), .B(carry[0]), .Z(B_AS[0]) );
endmodule


module address_conversion_M8_N4_N_bit64_F3_DW01_addsub_2 ( A, B, CI, ADD_SUB, 
        SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  FA_X1 U1_4 ( .A(A[4]), .B(B_AS[4]), .CI(carry[4]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA_X1 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA_X1 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA_X1 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0])
         );
  XOR2_X1 U1 ( .A(B[4]), .B(carry[0]), .Z(B_AS[4]) );
  XOR2_X1 U2 ( .A(B[3]), .B(carry[0]), .Z(B_AS[3]) );
  XOR2_X1 U3 ( .A(B[2]), .B(carry[0]), .Z(B_AS[2]) );
  XOR2_X1 U4 ( .A(B[1]), .B(carry[0]), .Z(B_AS[1]) );
  XOR2_X1 U5 ( .A(B[0]), .B(carry[0]), .Z(B_AS[0]) );
endmodule


module address_conversion_M8_N4_N_bit64_F3_DW01_add_0 ( A, B, CI, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI;
  output CO;
  wire   n4, n5, n6, n10, n11, n12;
  wire   [4:1] carry;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  AOI21_X1 U1 ( .B1(A[1]), .B2(B[1]), .A(n11), .ZN(n4) );
  INV_X1 U2 ( .A(n6), .ZN(n11) );
  OAI211_X1 U3 ( .C1(A[1]), .C2(B[1]), .A(A[0]), .B(B[0]), .ZN(n6) );
  OAI21_X1 U4 ( .B1(n4), .B2(n12), .A(n5), .ZN(carry[3]) );
  OAI21_X1 U5 ( .B1(A[2]), .B2(n10), .A(B[2]), .ZN(n5) );
  INV_X1 U6 ( .A(n4), .ZN(n10) );
  INV_X1 U7 ( .A(A[2]), .ZN(n12) );
endmodule


module address_conversion_M8_N4_N_bit64_F3_DW01_add_1 ( A, B, CI, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI;
  output CO;
  wire   n4, n5, n6, n10, n11, n12;
  wire   [4:1] carry;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  INV_X1 U1 ( .A(n6), .ZN(n11) );
  INV_X1 U2 ( .A(A[2]), .ZN(n12) );
  OAI21_X1 U3 ( .B1(A[2]), .B2(n10), .A(B[2]), .ZN(n5) );
  AOI21_X1 U4 ( .B1(A[1]), .B2(B[1]), .A(n11), .ZN(n4) );
  OAI211_X1 U5 ( .C1(A[1]), .C2(B[1]), .A(A[0]), .B(B[0]), .ZN(n6) );
  OAI21_X1 U6 ( .B1(n4), .B2(n12), .A(n5), .ZN(carry[3]) );
  INV_X1 U7 ( .A(n4), .ZN(n10) );
endmodule


module address_conversion_M8_N4_N_bit64_F3_DW01_add_2 ( A, B, CI, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI;
  output CO;
  wire   n4, n5, n6, n10, n11, n12;
  wire   [4:1] carry;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  INV_X1 U1 ( .A(A[2]), .ZN(n12) );
  OAI21_X1 U2 ( .B1(A[2]), .B2(n10), .A(B[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(A[1]), .B2(B[1]), .A(n11), .ZN(n4) );
  INV_X1 U4 ( .A(n6), .ZN(n11) );
  OAI211_X1 U5 ( .C1(A[1]), .C2(B[1]), .A(A[0]), .B(B[0]), .ZN(n6) );
  OAI21_X1 U6 ( .B1(n4), .B2(n12), .A(n5), .ZN(carry[3]) );
  INV_X1 U7 ( .A(n4), .ZN(n10) );
endmodule


module address_conversion_M8_N4_N_bit64_F3 ( spill_fill_count, wait_count, 
        start_write, clck, address_input_1, address_input_3, address_output_1, 
        address_output_2, address_output_3, swp, cwp );
  input [4:0] address_input_1;
  input [4:0] address_input_3;
  output [4:0] address_output_1;
  output [4:0] address_output_2;
  output [4:0] address_output_3;
  input [4:0] swp;
  input [4:0] cwp;
  input spill_fill_count, clck;
  output wait_count, start_write;
  wire   N15, N16, N45, N46, N77, N78, N91, N92, N93, N94, N95, N97, N98, N99,
         \U3/U1/Z_0 , \U3/U1/Z_1 , \U3/U1/Z_2 , \U3/U1/Z_3 , \U3/U1/Z_4 ,
         \U3/U2/Z_0 , \U3/U3/Z_0 , \U3/U3/Z_1 , \U3/U3/Z_2 , \U3/U3/Z_3 ,
         \U3/U3/Z_4 , \U3/U4/Z_0 , \U3/U5/Z_0 , \U3/U5/Z_1 , \U3/U5/Z_2 ,
         \U3/U5/Z_3 , \U3/U5/Z_4 , n76, \add_101/carry[4] , \add_101/carry[3] ,
         \add_101/carry[2] , n2, n20, n21, n22, n23, n24, n25, n27, n28, n30,
         n31, n33, n34, n35, n36, n42, n43, n44, n45, n46, n47, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66;
  wire   [4:0] ADDRESS_WRITE_cpu;
  wire   [4:0] i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8;

  DFFR_X1 wait_s_reg ( .D(1'b1), .CK(spill_fill_count), .RN(n36), .Q(
        wait_count) );
  DLL_X1 \ADDRESS_COUNT_reg[4]  ( .D(N95), .GN(n55), .Q(address_output_2[4])
         );
  DLL_X1 \ADDRESS_COUNT_reg[3]  ( .D(N94), .GN(n55), .Q(address_output_2[3])
         );
  DLL_X1 \ADDRESS_COUNT_reg[2]  ( .D(N93), .GN(n55), .Q(address_output_2[2])
         );
  DLL_X1 \ADDRESS_COUNT_reg[1]  ( .D(N92), .GN(n55), .Q(address_output_2[1])
         );
  DLL_X1 \ADDRESS_COUNT_reg[0]  ( .D(N91), .GN(n55), .Q(address_output_2[0])
         );
  DLL_X1 start_reg ( .D(n56), .GN(n76), .Q(start_write) );
  HA_X1 \add_101/U1_1_1  ( .A(i[1]), .B(i[0]), .CO(\add_101/carry[2] ), .S(N97) );
  HA_X1 \add_101/U1_1_2  ( .A(i[2]), .B(\add_101/carry[2] ), .CO(
        \add_101/carry[3] ), .S(N98) );
  HA_X1 \add_101/U1_1_3  ( .A(i[3]), .B(\add_101/carry[3] ), .CO(
        \add_101/carry[4] ), .S(N99) );
  MUX21_generic_N5 ADDRESS_multiplexer_write ( .A(address_output_2), .B(
        ADDRESS_WRITE_cpu), .sel(wait_count), .Y(address_output_3) );
  address_conversion_M8_N4_N_bit64_F3_DW01_addsub_0 r150 ( .A(address_input_1), 
        .B({\U3/U1/Z_4 , \U3/U1/Z_3 , \U3/U1/Z_2 , \U3/U1/Z_1 , \U3/U1/Z_0 }), 
        .CI(1'b0), .ADD_SUB(\U3/U2/Z_0 ), .SUM(address_output_1) );
  address_conversion_M8_N4_N_bit64_F3_DW01_addsub_1 r160 ( .A(address_input_3), 
        .B({\U3/U3/Z_4 , \U3/U3/Z_3 , \U3/U3/Z_2 , \U3/U3/Z_1 , \U3/U3/Z_0 }), 
        .CI(1'b0), .ADD_SUB(\U3/U4/Z_0 ), .SUM(ADDRESS_WRITE_cpu) );
  address_conversion_M8_N4_N_bit64_F3_DW01_addsub_2 r174 ( .A(i), .B({
        \U3/U5/Z_4 , \U3/U5/Z_3 , \U3/U5/Z_2 , \U3/U5/Z_1 , \U3/U5/Z_0 }), 
        .CI(1'b0), .ADD_SUB(n57), .SUM({N95, N94, N93, N92, N91}) );
  address_conversion_M8_N4_N_bit64_F3_DW01_add_0 add_96 ( .A(swp), .B(i), .CI(
        1'b0), .SUM({N78, N77, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2}) );
  address_conversion_M8_N4_N_bit64_F3_DW01_add_1 add_52 ( .A(address_input_1), 
        .B(cwp), .CI(1'b0), .SUM({N16, N15, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5}) );
  address_conversion_M8_N4_N_bit64_F3_DW01_add_2 add_61 ( .A(address_input_3), 
        .B(cwp), .CI(1'b0), .SUM({N46, N45, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8}) );
  DFFRS_X1 \i_reg[4]  ( .D(1'b0), .CK(spill_fill_count), .RN(n25), .SN(n27), 
        .Q(i[4]), .QN(n22) );
  DFFRS_X1 \i_reg[2]  ( .D(1'b0), .CK(spill_fill_count), .RN(n31), .SN(n33), 
        .Q(i[2]) );
  DFFRS_X1 \i_reg[0]  ( .D(1'b0), .CK(spill_fill_count), .RN(n23), .SN(n24), 
        .Q(i[0]), .QN(n21) );
  DFFRS_X1 \i_reg[3]  ( .D(1'b0), .CK(spill_fill_count), .RN(n28), .SN(n30), 
        .Q(i[3]), .QN(n20) );
  DFFRS_X1 \i_reg[1]  ( .D(1'b0), .CK(spill_fill_count), .RN(n34), .SN(n35), 
        .Q(i[1]) );
  OR2_X1 U3 ( .A1(n55), .A2(n21), .ZN(n23) );
  NAND2_X1 U4 ( .A1(n21), .A2(n2), .ZN(n24) );
  OR2_X1 U18 ( .A1(n56), .A2(n76), .ZN(n36) );
  OR2_X1 U12 ( .A1(n55), .A2(N98), .ZN(n31) );
  OR2_X1 U8 ( .A1(n55), .A2(N99), .ZN(n28) );
  OR2_X1 U15 ( .A1(n55), .A2(N97), .ZN(n34) );
  OR2_X1 U5 ( .A1(\add_101/carry[4] ), .A2(n55), .ZN(n25) );
  NAND2_X1 U6 ( .A1(\add_101/carry[4] ), .A2(n2), .ZN(n27) );
  NAND2_X1 U13 ( .A1(N98), .A2(n2), .ZN(n33) );
  NAND2_X1 U10 ( .A1(N99), .A2(n2), .ZN(n30) );
  NAND2_X1 U16 ( .A1(N97), .A2(n2), .ZN(n35) );
  INV_X1 U19 ( .A(n47), .ZN(n59) );
  INV_X1 U21 ( .A(n2), .ZN(n55) );
  INV_X1 U22 ( .A(n44), .ZN(n65) );
  AOI21_X1 U23 ( .B1(N15), .B2(N16), .A(n66), .ZN(n47) );
  INV_X1 U24 ( .A(n46), .ZN(n66) );
  AND3_X1 U25 ( .A1(N16), .A2(n46), .A3(N15), .ZN(\U3/U2/Z_0 ) );
  NOR2_X1 U26 ( .A1(n42), .A2(n76), .ZN(n2) );
  INV_X1 U27 ( .A(n43), .ZN(n57) );
  INV_X1 U28 ( .A(n42), .ZN(n56) );
  OAI21_X1 U29 ( .B1(n64), .B2(n59), .A(n46), .ZN(\U3/U1/Z_4 ) );
  NOR2_X1 U30 ( .A1(n61), .A2(n59), .ZN(\U3/U1/Z_2 ) );
  NOR2_X1 U31 ( .A1(n62), .A2(n59), .ZN(\U3/U1/Z_1 ) );
  NOR2_X1 U32 ( .A1(n63), .A2(n59), .ZN(\U3/U1/Z_0 ) );
  INV_X1 U33 ( .A(cwp[2]), .ZN(n61) );
  INV_X1 U34 ( .A(cwp[4]), .ZN(n64) );
  INV_X1 U35 ( .A(cwp[0]), .ZN(n63) );
  INV_X1 U36 ( .A(cwp[3]), .ZN(n60) );
  AOI21_X1 U37 ( .B1(address_input_1[3]), .B2(address_input_1[2]), .A(
        address_input_1[4]), .ZN(n46) );
  AOI21_X1 U38 ( .B1(address_input_3[3]), .B2(address_input_3[2]), .A(
        address_input_3[4]), .ZN(n44) );
  NAND2_X1 U39 ( .A1(N78), .A2(N77), .ZN(n43) );
  AND2_X1 U40 ( .A1(swp[0]), .A2(n43), .ZN(\U3/U5/Z_0 ) );
  AND2_X1 U41 ( .A1(swp[1]), .A2(n43), .ZN(\U3/U5/Z_1 ) );
  AND2_X1 U42 ( .A1(swp[2]), .A2(n43), .ZN(\U3/U5/Z_2 ) );
  OR2_X1 U43 ( .A1(n57), .A2(swp[3]), .ZN(\U3/U5/Z_3 ) );
  NAND2_X1 U44 ( .A1(n22), .A2(n20), .ZN(n42) );
  NAND2_X1 U45 ( .A1(wait_count), .A2(clck), .ZN(n76) );
  AND2_X1 U46 ( .A1(swp[4]), .A2(n43), .ZN(\U3/U5/Z_4 ) );
  INV_X1 U47 ( .A(cwp[1]), .ZN(n62) );
  AND3_X1 U48 ( .A1(N46), .A2(n44), .A3(N45), .ZN(\U3/U4/Z_0 ) );
  NAND2_X1 U49 ( .A1(n47), .A2(n60), .ZN(\U3/U1/Z_3 ) );
  AOI21_X1 U50 ( .B1(N45), .B2(N46), .A(n65), .ZN(n45) );
  OAI21_X1 U51 ( .B1(n58), .B2(n64), .A(n44), .ZN(\U3/U3/Z_4 ) );
  NAND2_X1 U52 ( .A1(n45), .A2(n60), .ZN(\U3/U3/Z_3 ) );
  NOR2_X1 U53 ( .A1(n58), .A2(n61), .ZN(\U3/U3/Z_2 ) );
  NOR2_X1 U54 ( .A1(n58), .A2(n62), .ZN(\U3/U3/Z_1 ) );
  INV_X1 U55 ( .A(n45), .ZN(n58) );
  NOR2_X1 U56 ( .A1(n58), .A2(n63), .ZN(\U3/U3/Z_0 ) );
endmodule


module MUX21_generic_N64 ( A, B, sel, Y );
  input [63:0] A;
  input [63:0] B;
  output [63:0] Y;
  input sel;
  wire   n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246;

  INV_X1 U1 ( .A(n243), .ZN(n221) );
  INV_X1 U2 ( .A(n243), .ZN(n222) );
  INV_X1 U3 ( .A(n243), .ZN(n223) );
  INV_X1 U4 ( .A(n243), .ZN(n224) );
  INV_X1 U5 ( .A(n243), .ZN(n225) );
  BUF_X1 U6 ( .A(n244), .Z(n243) );
  BUF_X1 U7 ( .A(n245), .Z(n234) );
  BUF_X1 U8 ( .A(n245), .Z(n233) );
  BUF_X1 U9 ( .A(n245), .Z(n232) );
  BUF_X1 U10 ( .A(n246), .Z(n242) );
  BUF_X1 U11 ( .A(n245), .Z(n241) );
  BUF_X1 U12 ( .A(n245), .Z(n240) );
  BUF_X1 U13 ( .A(n244), .Z(n239) );
  BUF_X1 U14 ( .A(n245), .Z(n238) );
  BUF_X1 U15 ( .A(n244), .Z(n237) );
  BUF_X1 U16 ( .A(n244), .Z(n236) );
  BUF_X1 U17 ( .A(n244), .Z(n235) );
  BUF_X1 U18 ( .A(n246), .Z(n231) );
  BUF_X1 U19 ( .A(n246), .Z(n230) );
  BUF_X1 U20 ( .A(n246), .Z(n229) );
  BUF_X1 U21 ( .A(n246), .Z(n228) );
  BUF_X1 U22 ( .A(n246), .Z(n227) );
  INV_X1 U23 ( .A(n220), .ZN(n245) );
  INV_X1 U24 ( .A(n220), .ZN(n244) );
  INV_X1 U25 ( .A(n220), .ZN(n246) );
  BUF_X1 U26 ( .A(sel), .Z(n220) );
  INV_X1 U27 ( .A(n66), .ZN(Y[63]) );
  AOI22_X1 U28 ( .A1(n226), .A2(A[63]), .B1(B[63]), .B2(n227), .ZN(n66) );
  INV_X1 U29 ( .A(n100), .ZN(Y[29]) );
  AOI22_X1 U30 ( .A1(A[29]), .A2(n223), .B1(B[29]), .B2(n235), .ZN(n100) );
  INV_X1 U31 ( .A(n99), .ZN(Y[30]) );
  AOI22_X1 U32 ( .A1(A[30]), .A2(n223), .B1(B[30]), .B2(n235), .ZN(n99) );
  INV_X1 U33 ( .A(n98), .ZN(Y[31]) );
  AOI22_X1 U34 ( .A1(A[31]), .A2(n223), .B1(B[31]), .B2(n235), .ZN(n98) );
  INV_X1 U35 ( .A(n97), .ZN(Y[32]) );
  AOI22_X1 U36 ( .A1(A[32]), .A2(n223), .B1(B[32]), .B2(n234), .ZN(n97) );
  INV_X1 U37 ( .A(n96), .ZN(Y[33]) );
  AOI22_X1 U38 ( .A1(A[33]), .A2(n223), .B1(B[33]), .B2(n234), .ZN(n96) );
  INV_X1 U39 ( .A(n95), .ZN(Y[34]) );
  AOI22_X1 U40 ( .A1(A[34]), .A2(n223), .B1(B[34]), .B2(n234), .ZN(n95) );
  INV_X1 U41 ( .A(n94), .ZN(Y[35]) );
  AOI22_X1 U42 ( .A1(A[35]), .A2(n223), .B1(B[35]), .B2(n234), .ZN(n94) );
  INV_X1 U43 ( .A(n93), .ZN(Y[36]) );
  AOI22_X1 U44 ( .A1(A[36]), .A2(n224), .B1(B[36]), .B2(n233), .ZN(n93) );
  INV_X1 U45 ( .A(n92), .ZN(Y[37]) );
  AOI22_X1 U46 ( .A1(A[37]), .A2(n224), .B1(B[37]), .B2(n233), .ZN(n92) );
  INV_X1 U47 ( .A(n91), .ZN(Y[38]) );
  AOI22_X1 U48 ( .A1(A[38]), .A2(n224), .B1(B[38]), .B2(n233), .ZN(n91) );
  INV_X1 U49 ( .A(n90), .ZN(Y[39]) );
  AOI22_X1 U50 ( .A1(A[39]), .A2(n224), .B1(B[39]), .B2(n233), .ZN(n90) );
  INV_X1 U51 ( .A(n89), .ZN(Y[40]) );
  AOI22_X1 U52 ( .A1(A[40]), .A2(n224), .B1(B[40]), .B2(n232), .ZN(n89) );
  INV_X1 U53 ( .A(n88), .ZN(Y[41]) );
  AOI22_X1 U54 ( .A1(A[41]), .A2(n224), .B1(B[41]), .B2(n232), .ZN(n88) );
  INV_X1 U55 ( .A(n87), .ZN(Y[42]) );
  AOI22_X1 U56 ( .A1(A[42]), .A2(n224), .B1(B[42]), .B2(n232), .ZN(n87) );
  INV_X1 U57 ( .A(n86), .ZN(Y[43]) );
  AOI22_X1 U58 ( .A1(A[43]), .A2(n224), .B1(B[43]), .B2(n232), .ZN(n86) );
  INV_X1 U59 ( .A(n85), .ZN(Y[44]) );
  AOI22_X1 U60 ( .A1(A[44]), .A2(n224), .B1(B[44]), .B2(n231), .ZN(n85) );
  INV_X1 U61 ( .A(n84), .ZN(Y[45]) );
  AOI22_X1 U62 ( .A1(A[45]), .A2(n224), .B1(B[45]), .B2(n231), .ZN(n84) );
  INV_X1 U63 ( .A(n74), .ZN(Y[55]) );
  AOI22_X1 U64 ( .A1(A[55]), .A2(n225), .B1(B[55]), .B2(n229), .ZN(n74) );
  INV_X1 U65 ( .A(n73), .ZN(Y[56]) );
  AOI22_X1 U66 ( .A1(A[56]), .A2(n225), .B1(B[56]), .B2(n228), .ZN(n73) );
  INV_X1 U67 ( .A(n72), .ZN(Y[57]) );
  AOI22_X1 U68 ( .A1(A[57]), .A2(n225), .B1(B[57]), .B2(n228), .ZN(n72) );
  INV_X1 U69 ( .A(n71), .ZN(Y[58]) );
  AOI22_X1 U70 ( .A1(A[58]), .A2(n225), .B1(B[58]), .B2(n228), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(Y[59]) );
  AOI22_X1 U72 ( .A1(A[59]), .A2(n225), .B1(B[59]), .B2(n228), .ZN(n70) );
  INV_X1 U73 ( .A(n129), .ZN(Y[0]) );
  AOI22_X1 U74 ( .A1(A[0]), .A2(n221), .B1(B[0]), .B2(n242), .ZN(n129) );
  INV_X1 U75 ( .A(n128), .ZN(Y[1]) );
  AOI22_X1 U76 ( .A1(A[1]), .A2(n221), .B1(B[1]), .B2(n242), .ZN(n128) );
  INV_X1 U77 ( .A(n127), .ZN(Y[2]) );
  AOI22_X1 U78 ( .A1(A[2]), .A2(n221), .B1(B[2]), .B2(n242), .ZN(n127) );
  INV_X1 U79 ( .A(n126), .ZN(Y[3]) );
  AOI22_X1 U80 ( .A1(A[3]), .A2(n221), .B1(B[3]), .B2(n242), .ZN(n126) );
  INV_X1 U81 ( .A(n125), .ZN(Y[4]) );
  AOI22_X1 U82 ( .A1(A[4]), .A2(n221), .B1(B[4]), .B2(n241), .ZN(n125) );
  INV_X1 U83 ( .A(n124), .ZN(Y[5]) );
  AOI22_X1 U84 ( .A1(A[5]), .A2(n221), .B1(B[5]), .B2(n241), .ZN(n124) );
  INV_X1 U85 ( .A(n123), .ZN(Y[6]) );
  AOI22_X1 U86 ( .A1(A[6]), .A2(n221), .B1(B[6]), .B2(n241), .ZN(n123) );
  INV_X1 U87 ( .A(n122), .ZN(Y[7]) );
  AOI22_X1 U88 ( .A1(A[7]), .A2(n221), .B1(B[7]), .B2(n241), .ZN(n122) );
  INV_X1 U89 ( .A(n121), .ZN(Y[8]) );
  AOI22_X1 U90 ( .A1(A[8]), .A2(n221), .B1(B[8]), .B2(n240), .ZN(n121) );
  INV_X1 U91 ( .A(n120), .ZN(Y[9]) );
  AOI22_X1 U92 ( .A1(A[9]), .A2(n221), .B1(B[9]), .B2(n240), .ZN(n120) );
  INV_X1 U93 ( .A(n119), .ZN(Y[10]) );
  AOI22_X1 U94 ( .A1(A[10]), .A2(n221), .B1(B[10]), .B2(n240), .ZN(n119) );
  INV_X1 U95 ( .A(n118), .ZN(Y[11]) );
  AOI22_X1 U96 ( .A1(A[11]), .A2(n221), .B1(B[11]), .B2(n240), .ZN(n118) );
  INV_X1 U97 ( .A(n117), .ZN(Y[12]) );
  AOI22_X1 U98 ( .A1(A[12]), .A2(n222), .B1(B[12]), .B2(n239), .ZN(n117) );
  INV_X1 U99 ( .A(n116), .ZN(Y[13]) );
  AOI22_X1 U100 ( .A1(A[13]), .A2(n222), .B1(B[13]), .B2(n239), .ZN(n116) );
  INV_X1 U101 ( .A(n115), .ZN(Y[14]) );
  AOI22_X1 U102 ( .A1(A[14]), .A2(n222), .B1(B[14]), .B2(n239), .ZN(n115) );
  INV_X1 U103 ( .A(n114), .ZN(Y[15]) );
  AOI22_X1 U104 ( .A1(A[15]), .A2(n222), .B1(B[15]), .B2(n239), .ZN(n114) );
  INV_X1 U105 ( .A(n113), .ZN(Y[16]) );
  AOI22_X1 U106 ( .A1(A[16]), .A2(n222), .B1(B[16]), .B2(n238), .ZN(n113) );
  INV_X1 U107 ( .A(n112), .ZN(Y[17]) );
  AOI22_X1 U108 ( .A1(A[17]), .A2(n222), .B1(B[17]), .B2(n238), .ZN(n112) );
  INV_X1 U109 ( .A(n111), .ZN(Y[18]) );
  AOI22_X1 U110 ( .A1(A[18]), .A2(n222), .B1(B[18]), .B2(n238), .ZN(n111) );
  INV_X1 U111 ( .A(n110), .ZN(Y[19]) );
  AOI22_X1 U112 ( .A1(A[19]), .A2(n222), .B1(B[19]), .B2(n238), .ZN(n110) );
  INV_X1 U113 ( .A(n109), .ZN(Y[20]) );
  AOI22_X1 U114 ( .A1(A[20]), .A2(n222), .B1(B[20]), .B2(n237), .ZN(n109) );
  INV_X1 U115 ( .A(n108), .ZN(Y[21]) );
  AOI22_X1 U116 ( .A1(A[21]), .A2(n222), .B1(B[21]), .B2(n237), .ZN(n108) );
  INV_X1 U117 ( .A(n107), .ZN(Y[22]) );
  AOI22_X1 U118 ( .A1(A[22]), .A2(n222), .B1(B[22]), .B2(n237), .ZN(n107) );
  INV_X1 U119 ( .A(n106), .ZN(Y[23]) );
  AOI22_X1 U120 ( .A1(A[23]), .A2(n222), .B1(B[23]), .B2(n237), .ZN(n106) );
  INV_X1 U121 ( .A(n105), .ZN(Y[24]) );
  AOI22_X1 U122 ( .A1(A[24]), .A2(n223), .B1(B[24]), .B2(n236), .ZN(n105) );
  INV_X1 U123 ( .A(n104), .ZN(Y[25]) );
  AOI22_X1 U124 ( .A1(A[25]), .A2(n223), .B1(B[25]), .B2(n236), .ZN(n104) );
  INV_X1 U125 ( .A(n103), .ZN(Y[26]) );
  AOI22_X1 U126 ( .A1(A[26]), .A2(n223), .B1(B[26]), .B2(n236), .ZN(n103) );
  INV_X1 U127 ( .A(n102), .ZN(Y[27]) );
  AOI22_X1 U128 ( .A1(A[27]), .A2(n223), .B1(B[27]), .B2(n236), .ZN(n102) );
  INV_X1 U129 ( .A(n101), .ZN(Y[28]) );
  AOI22_X1 U130 ( .A1(A[28]), .A2(n223), .B1(B[28]), .B2(n235), .ZN(n101) );
  INV_X1 U131 ( .A(n83), .ZN(Y[46]) );
  AOI22_X1 U132 ( .A1(A[46]), .A2(n224), .B1(B[46]), .B2(n231), .ZN(n83) );
  INV_X1 U133 ( .A(n82), .ZN(Y[47]) );
  AOI22_X1 U134 ( .A1(A[47]), .A2(n224), .B1(B[47]), .B2(n231), .ZN(n82) );
  INV_X1 U135 ( .A(n81), .ZN(Y[48]) );
  AOI22_X1 U136 ( .A1(A[48]), .A2(n225), .B1(B[48]), .B2(n230), .ZN(n81) );
  INV_X1 U137 ( .A(n80), .ZN(Y[49]) );
  AOI22_X1 U138 ( .A1(A[49]), .A2(n225), .B1(B[49]), .B2(n230), .ZN(n80) );
  INV_X1 U139 ( .A(n79), .ZN(Y[50]) );
  AOI22_X1 U140 ( .A1(A[50]), .A2(n225), .B1(B[50]), .B2(n230), .ZN(n79) );
  INV_X1 U141 ( .A(n78), .ZN(Y[51]) );
  AOI22_X1 U142 ( .A1(A[51]), .A2(n225), .B1(B[51]), .B2(n230), .ZN(n78) );
  INV_X1 U143 ( .A(n77), .ZN(Y[52]) );
  AOI22_X1 U144 ( .A1(A[52]), .A2(n225), .B1(B[52]), .B2(n229), .ZN(n77) );
  INV_X1 U145 ( .A(n76), .ZN(Y[53]) );
  AOI22_X1 U146 ( .A1(A[53]), .A2(n225), .B1(B[53]), .B2(n229), .ZN(n76) );
  INV_X1 U147 ( .A(n75), .ZN(Y[54]) );
  AOI22_X1 U148 ( .A1(A[54]), .A2(n225), .B1(B[54]), .B2(n229), .ZN(n75) );
  INV_X1 U149 ( .A(n69), .ZN(Y[60]) );
  AOI22_X1 U150 ( .A1(A[60]), .A2(n226), .B1(B[60]), .B2(n227), .ZN(n69) );
  INV_X1 U151 ( .A(n68), .ZN(Y[61]) );
  AOI22_X1 U152 ( .A1(A[61]), .A2(n226), .B1(B[61]), .B2(n227), .ZN(n68) );
  INV_X1 U153 ( .A(n67), .ZN(Y[62]) );
  AOI22_X1 U154 ( .A1(A[62]), .A2(n226), .B1(B[62]), .B2(n227), .ZN(n67) );
  INV_X1 U155 ( .A(n243), .ZN(n226) );
endmodule


module windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_2 ( A, INC_DEC, SUM
 );
  input [31:0] A;
  output [31:0] SUM;
  input INC_DEC;
  wire   n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n360,
         n361;

  XOR2_X1 U128 ( .A(n241), .B(INC_DEC), .Z(n247) );
  XOR2_X1 U129 ( .A(n249), .B(n227), .Z(SUM[8]) );
  XOR2_X1 U130 ( .A(n239), .B(INC_DEC), .Z(n249) );
  XOR2_X1 U131 ( .A(n250), .B(n251), .Z(SUM[7]) );
  XOR2_X1 U132 ( .A(INC_DEC), .B(A[7]), .Z(n251) );
  XOR2_X1 U133 ( .A(n255), .B(n252), .Z(SUM[6]) );
  XOR2_X1 U134 ( .A(n256), .B(n258), .Z(SUM[5]) );
  XOR2_X1 U135 ( .A(n261), .B(n262), .Z(SUM[4]) );
  XOR2_X1 U136 ( .A(INC_DEC), .B(A[4]), .Z(n262) );
  XOR2_X1 U137 ( .A(n263), .B(n264), .Z(SUM[3]) );
  XOR2_X1 U138 ( .A(INC_DEC), .B(A[3]), .Z(n264) );
  XOR2_X1 U139 ( .A(n268), .B(n269), .Z(SUM[31]) );
  XOR2_X1 U140 ( .A(INC_DEC), .B(A[31]), .Z(n269) );
  XOR2_X1 U141 ( .A(INC_DEC), .B(A[30]), .Z(n272) );
  XOR2_X1 U142 ( .A(n274), .B(n265), .Z(SUM[2]) );
  XOR2_X1 U143 ( .A(n222), .B(n276), .Z(SUM[29]) );
  XOR2_X1 U144 ( .A(INC_DEC), .B(A[29]), .Z(n276) );
  XOR2_X1 U145 ( .A(n278), .B(n280), .Z(SUM[28]) );
  XOR2_X1 U146 ( .A(INC_DEC), .B(A[28]), .Z(n280) );
  XOR2_X1 U147 ( .A(n287), .B(n288), .Z(SUM[27]) );
  XOR2_X1 U148 ( .A(n217), .B(A[27]), .Z(n288) );
  XOR2_X1 U149 ( .A(n286), .B(n295), .Z(SUM[24]) );
  XOR2_X1 U150 ( .A(INC_DEC), .B(A[24]), .Z(n295) );
  XOR2_X1 U151 ( .A(n302), .B(n303), .Z(SUM[23]) );
  XOR2_X1 U152 ( .A(A[23]), .B(n219), .Z(n302) );
  XOR2_X1 U153 ( .A(n304), .B(n306), .Z(SUM[22]) );
  XOR2_X1 U154 ( .A(n309), .B(n307), .Z(SUM[21]) );
  XOR2_X1 U155 ( .A(A[20]), .B(n219), .Z(n310) );
  XOR2_X1 U156 ( .A(A[0]), .B(n316), .Z(SUM[1]) );
  XOR2_X1 U157 ( .A(INC_DEC), .B(A[1]), .Z(n316) );
  XOR2_X1 U158 ( .A(INC_DEC), .B(A[19]), .Z(n318) );
  XOR2_X1 U159 ( .A(n319), .B(n321), .Z(SUM[18]) );
  XOR2_X1 U160 ( .A(n217), .B(A[18]), .Z(n321) );
  XOR2_X1 U161 ( .A(n217), .B(A[17]), .Z(n324) );
  XOR2_X1 U162 ( .A(n313), .B(n325), .Z(SUM[16]) );
  XOR2_X1 U163 ( .A(n217), .B(A[16]), .Z(n325) );
  XOR2_X1 U164 ( .A(n336), .B(n337), .Z(SUM[15]) );
  XOR2_X1 U165 ( .A(n217), .B(A[15]), .Z(n337) );
  XOR2_X1 U166 ( .A(n217), .B(A[14]), .Z(n340) );
  XOR2_X1 U167 ( .A(n217), .B(A[13]), .Z(n343) );
  XOR2_X1 U168 ( .A(n344), .B(n346), .Z(SUM[12]) );
  XOR2_X1 U169 ( .A(n217), .B(A[12]), .Z(n346) );
  XOR2_X1 U170 ( .A(n349), .B(n350), .Z(SUM[11]) );
  XOR2_X1 U171 ( .A(n246), .B(INC_DEC), .Z(n349) );
  XOR2_X1 U172 ( .A(n353), .B(n352), .Z(SUM[10]) );
  NAND3_X1 U173 ( .A1(n333), .A2(n267), .A3(n358), .ZN(n261) );
  XOR2_X1 U174 ( .A(n245), .B(INC_DEC), .Z(n353) );
  INV_X1 U1 ( .A(INC_DEC), .ZN(n219) );
  OAI21_X1 U2 ( .B1(n227), .B2(n347), .A(n329), .ZN(n344) );
  NOR2_X1 U3 ( .A1(n330), .A2(n217), .ZN(n347) );
  INV_X1 U4 ( .A(n356), .ZN(n227) );
  NOR4_X1 U5 ( .A1(n246), .A2(n245), .A3(n241), .A4(n239), .ZN(n330) );
  NOR4_X1 U6 ( .A1(n332), .A2(n242), .A3(n244), .A4(n360), .ZN(n331) );
  NAND4_X1 U7 ( .A1(n245), .A2(n246), .A3(n239), .A4(n241), .ZN(n348) );
  OAI21_X1 U8 ( .B1(n332), .B2(n230), .A(n326), .ZN(n356) );
  AOI21_X1 U9 ( .B1(n235), .B2(n256), .A(n231), .ZN(n252) );
  INV_X1 U10 ( .A(n257), .ZN(n235) );
  AOI21_X1 U11 ( .B1(n304), .B2(n232), .A(n233), .ZN(n303) );
  INV_X1 U12 ( .A(n305), .ZN(n232) );
  OAI21_X1 U13 ( .B1(n289), .B2(n290), .A(n282), .ZN(n287) );
  NAND4_X1 U14 ( .A1(SUM[0]), .A2(n242), .A3(n244), .A4(n360), .ZN(n335) );
  INV_X1 U15 ( .A(n261), .ZN(n230) );
  INV_X1 U16 ( .A(n297), .ZN(n233) );
  INV_X1 U17 ( .A(n259), .ZN(n231) );
  INV_X1 U18 ( .A(n339), .ZN(n225) );
  INV_X1 U19 ( .A(n282), .ZN(n234) );
  OAI22_X1 U20 ( .A1(n227), .A2(n239), .B1(n355), .B2(n219), .ZN(n248) );
  NOR2_X1 U21 ( .A1(A[8]), .A2(n356), .ZN(n355) );
  AOI22_X1 U22 ( .A1(n344), .A2(A[12]), .B1(n345), .B2(n218), .ZN(n341) );
  OR2_X1 U23 ( .A1(A[12]), .A2(n344), .ZN(n345) );
  AOI22_X1 U24 ( .A1(n313), .A2(A[16]), .B1(n315), .B2(n218), .ZN(n322) );
  INV_X1 U25 ( .A(n299), .ZN(n220) );
  AOI22_X1 U26 ( .A1(n248), .A2(A[9]), .B1(n354), .B2(n218), .ZN(n352) );
  OR2_X1 U27 ( .A1(A[9]), .A2(n248), .ZN(n354) );
  OAI21_X1 U28 ( .B1(n322), .B2(n240), .A(n323), .ZN(n319) );
  INV_X1 U29 ( .A(A[17]), .ZN(n240) );
  OAI21_X1 U30 ( .B1(A[17]), .B2(n229), .A(n218), .ZN(n323) );
  INV_X1 U31 ( .A(n322), .ZN(n229) );
  AOI22_X1 U32 ( .A1(n222), .A2(A[29]), .B1(n273), .B2(n218), .ZN(n271) );
  OR2_X1 U33 ( .A1(n222), .A2(A[29]), .ZN(n273) );
  NAND4_X1 U34 ( .A1(n326), .A2(n327), .A3(n328), .A4(n329), .ZN(n313) );
  NAND4_X1 U35 ( .A1(n237), .A2(A[15]), .A3(n330), .A4(n331), .ZN(n328) );
  OAI21_X1 U36 ( .B1(n334), .B2(n335), .A(n218), .ZN(n327) );
  INV_X1 U37 ( .A(n333), .ZN(n237) );
  OAI21_X1 U38 ( .B1(A[3]), .B2(n275), .A(n217), .ZN(n358) );
  OAI21_X1 U39 ( .B1(n311), .B2(n219), .A(n312), .ZN(n301) );
  NAND4_X1 U40 ( .A1(A[16]), .A2(n313), .A3(A[17]), .A4(n314), .ZN(n312) );
  NOR4_X1 U41 ( .A1(A[19]), .A2(A[18]), .A3(A[17]), .A4(n315), .ZN(n311) );
  AND2_X1 U42 ( .A1(A[18]), .A2(A[19]), .ZN(n314) );
  NOR2_X1 U43 ( .A1(n257), .A2(n231), .ZN(n258) );
  NOR2_X1 U44 ( .A1(n217), .A2(A[5]), .ZN(n257) );
  OAI21_X1 U45 ( .B1(n221), .B2(n243), .A(n284), .ZN(n293) );
  INV_X1 U46 ( .A(A[24]), .ZN(n243) );
  AOI21_X1 U47 ( .B1(n238), .B2(n230), .A(n260), .ZN(n256) );
  INV_X1 U48 ( .A(A[4]), .ZN(n238) );
  AOI21_X1 U49 ( .B1(n261), .B2(A[4]), .A(n218), .ZN(n260) );
  OAI21_X1 U50 ( .B1(n341), .B2(n244), .A(n342), .ZN(n339) );
  OAI21_X1 U51 ( .B1(A[13]), .B2(n226), .A(n218), .ZN(n342) );
  INV_X1 U52 ( .A(n341), .ZN(n226) );
  AOI22_X1 U53 ( .A1(n218), .A2(n351), .B1(A[10]), .B2(n224), .ZN(n350) );
  NAND2_X1 U54 ( .A1(n352), .A2(n245), .ZN(n351) );
  INV_X1 U55 ( .A(n352), .ZN(n224) );
  INV_X1 U56 ( .A(A[30]), .ZN(n361) );
  NAND4_X1 U57 ( .A1(n281), .A2(n282), .A3(n283), .A4(n284), .ZN(n278) );
  OAI21_X1 U58 ( .B1(n285), .B2(n217), .A(A[27]), .ZN(n281) );
  NAND2_X1 U59 ( .A1(A[21]), .A2(n217), .ZN(n298) );
  NAND2_X1 U60 ( .A1(A[26]), .A2(n217), .ZN(n282) );
  NAND4_X1 U61 ( .A1(n296), .A2(n297), .A3(n298), .A4(n299), .ZN(n286) );
  OAI21_X1 U62 ( .B1(n300), .B2(n217), .A(A[23]), .ZN(n296) );
  OAI21_X1 U63 ( .B1(n307), .B2(n308), .A(n298), .ZN(n304) );
  NOR2_X1 U64 ( .A1(A[21]), .A2(n217), .ZN(n308) );
  NAND2_X1 U65 ( .A1(A[25]), .A2(n218), .ZN(n283) );
  NAND2_X1 U66 ( .A1(A[2]), .A2(n217), .ZN(n267) );
  AOI21_X1 U67 ( .B1(n319), .B2(A[18]), .A(n228), .ZN(n317) );
  INV_X1 U68 ( .A(n320), .ZN(n228) );
  OAI21_X1 U69 ( .B1(A[18]), .B2(n319), .A(n218), .ZN(n320) );
  NOR2_X1 U70 ( .A1(A[6]), .A2(n218), .ZN(n253) );
  NAND2_X1 U71 ( .A1(A[22]), .A2(n217), .ZN(n297) );
  NAND4_X1 U72 ( .A1(A[3]), .A2(A[1]), .A3(A[2]), .A4(A[0]), .ZN(n333) );
  OAI21_X1 U73 ( .B1(n225), .B2(n360), .A(n338), .ZN(n336) );
  OAI21_X1 U74 ( .B1(A[14]), .B2(n339), .A(n217), .ZN(n338) );
  NAND2_X1 U75 ( .A1(A[5]), .A2(n218), .ZN(n259) );
  INV_X1 U76 ( .A(A[8]), .ZN(n239) );
  INV_X1 U77 ( .A(A[10]), .ZN(n245) );
  OR4_X1 U78 ( .A1(A[15]), .A2(A[1]), .A3(A[2]), .A4(A[3]), .ZN(n334) );
  INV_X1 U79 ( .A(A[14]), .ZN(n360) );
  XNOR2_X1 U80 ( .A(n225), .B(n340), .ZN(SUM[14]) );
  XNOR2_X1 U81 ( .A(n341), .B(n343), .ZN(SUM[13]) );
  INV_X1 U82 ( .A(A[13]), .ZN(n244) );
  XNOR2_X1 U83 ( .A(n290), .B(n291), .ZN(SUM[26]) );
  NOR2_X1 U84 ( .A1(n289), .A2(n234), .ZN(n291) );
  XNOR2_X1 U85 ( .A(n293), .B(n294), .ZN(SUM[25]) );
  OAI21_X1 U86 ( .B1(A[25]), .B2(n217), .A(n283), .ZN(n294) );
  NOR2_X1 U87 ( .A1(n305), .A2(n233), .ZN(n306) );
  XNOR2_X1 U88 ( .A(n317), .B(n318), .ZN(SUM[19]) );
  OAI21_X1 U89 ( .B1(n218), .B2(A[21]), .A(n298), .ZN(n309) );
  XNOR2_X1 U90 ( .A(n247), .B(n248), .ZN(SUM[9]) );
  XNOR2_X1 U91 ( .A(n322), .B(n324), .ZN(SUM[17]) );
  INV_X1 U92 ( .A(A[9]), .ZN(n241) );
  INV_X1 U93 ( .A(A[11]), .ZN(n246) );
  AND3_X1 U94 ( .A1(n259), .A2(n254), .A3(n357), .ZN(n326) );
  OAI21_X1 U95 ( .B1(A[4]), .B2(A[7]), .A(n218), .ZN(n357) );
  AND2_X1 U96 ( .A1(n283), .A2(n292), .ZN(n290) );
  OAI21_X1 U97 ( .B1(A[25]), .B2(n217), .A(n293), .ZN(n292) );
  AND2_X1 U98 ( .A1(n359), .A2(n219), .ZN(n332) );
  NAND4_X1 U99 ( .A1(A[7]), .A2(A[4]), .A3(A[5]), .A4(A[6]), .ZN(n359) );
  INV_X1 U100 ( .A(n277), .ZN(n222) );
  OAI21_X1 U101 ( .B1(A[28]), .B2(n278), .A(n223), .ZN(n277) );
  INV_X1 U102 ( .A(n279), .ZN(n223) );
  AOI21_X1 U103 ( .B1(n278), .B2(A[28]), .A(n218), .ZN(n279) );
  INV_X1 U104 ( .A(A[0]), .ZN(SUM[0]) );
  INV_X1 U105 ( .A(A[12]), .ZN(n242) );
  OR2_X1 U106 ( .A1(n313), .A2(A[16]), .ZN(n315) );
  OR2_X1 U107 ( .A1(A[1]), .A2(A[0]), .ZN(n275) );
  AOI22_X1 U108 ( .A1(A[0]), .A2(A[1]), .B1(n275), .B2(n218), .ZN(n265) );
  NOR2_X1 U109 ( .A1(n217), .A2(A[22]), .ZN(n305) );
  NOR2_X1 U110 ( .A1(n217), .A2(A[26]), .ZN(n289) );
  OAI21_X1 U111 ( .B1(n265), .B2(n266), .A(n267), .ZN(n263) );
  NOR2_X1 U112 ( .A1(A[2]), .A2(n217), .ZN(n266) );
  OAI21_X1 U113 ( .B1(n218), .B2(A[2]), .A(n267), .ZN(n274) );
  XNOR2_X1 U114 ( .A(n310), .B(n301), .ZN(SUM[20]) );
  XNOR2_X1 U115 ( .A(n271), .B(n272), .ZN(SUM[30]) );
  OAI21_X1 U116 ( .B1(n252), .B2(n253), .A(n254), .ZN(n250) );
  OAI21_X1 U117 ( .B1(n218), .B2(A[6]), .A(n254), .ZN(n255) );
  AOI22_X1 U118 ( .A1(n270), .A2(n219), .B1(n271), .B2(n361), .ZN(n268) );
  OR2_X1 U119 ( .A1(n361), .A2(n271), .ZN(n270) );
  AOI21_X1 U120 ( .B1(n301), .B2(A[20]), .A(n220), .ZN(n307) );
  INV_X1 U121 ( .A(n286), .ZN(n221) );
  OAI21_X1 U122 ( .B1(A[24]), .B2(n286), .A(n218), .ZN(n284) );
  AND4_X1 U123 ( .A1(n286), .A2(A[25]), .A3(A[26]), .A4(A[24]), .ZN(n285) );
  OAI21_X1 U124 ( .B1(A[20]), .B2(n301), .A(n218), .ZN(n299) );
  AND4_X1 U125 ( .A1(n301), .A2(A[21]), .A3(A[22]), .A4(A[20]), .ZN(n300) );
  NAND2_X1 U126 ( .A1(n218), .A2(n348), .ZN(n329) );
  NAND2_X1 U127 ( .A1(INC_DEC), .A2(A[6]), .ZN(n254) );
  INV_X1 U175 ( .A(n219), .ZN(n217) );
  INV_X1 U176 ( .A(n219), .ZN(n218) );
endmodule


module windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_3 ( A, INC_DEC, SUM
 );
  input [31:0] A;
  output [31:0] SUM;
  input INC_DEC;
  wire   n1, n2, n3, n4, n5, n6, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n36, n37, n38,
         n39, n40, n41, n42, n43, n46, n47, n48, n49, n50, n51, n52, n53, n55,
         n56, n59, n60, n61, n62, n65, n66, n68, n69, n70, n71, n72, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n88, n90, n92,
         n93, n94, n95, n96, n98, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n114, n116, n118, n119, n120,
         n121, n122, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n138, n139, n140, n143, n145, n146, n147,
         n149, n150, n151, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n174, n175, n176, n177, n179, n182, n184, n185, n186, n188,
         n190, n191, n192, n193, n195, n196, n198, n199, n200, n201, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269;

  XOR2_X1 U183 ( .A(INC_DEC), .B(A[31]), .Z(n6) );
  NAND3_X1 U225 ( .A1(n83), .A2(n84), .A3(n85), .ZN(n75) );
  NAND3_X1 U227 ( .A1(n109), .A2(n110), .A3(n111), .ZN(n101) );
  NAND3_X1 U230 ( .A1(n134), .A2(n135), .A3(n136), .ZN(n126) );
  NAND3_X1 U244 ( .A1(n46), .A2(n65), .A3(n50), .ZN(n157) );
  INV_X1 U1 ( .A(n19), .ZN(n226) );
  BUF_X1 U2 ( .A(n221), .Z(n216) );
  BUF_X1 U3 ( .A(n221), .Z(n215) );
  BUF_X1 U4 ( .A(n221), .Z(n217) );
  BUF_X1 U5 ( .A(n221), .Z(n218) );
  BUF_X1 U6 ( .A(n221), .Z(n220) );
  BUF_X1 U7 ( .A(n221), .Z(n219) );
  NAND2_X1 U8 ( .A1(n154), .A2(n155), .ZN(n150) );
  NOR2_X1 U9 ( .A1(n156), .A2(n157), .ZN(n155) );
  AOI21_X1 U10 ( .B1(n158), .B2(n159), .A(n160), .ZN(n154) );
  NAND2_X1 U11 ( .A1(n2), .A2(n1), .ZN(n156) );
  OAI21_X1 U12 ( .B1(n227), .B2(n165), .A(n1), .ZN(n19) );
  INV_X1 U13 ( .A(n39), .ZN(n227) );
  OAI21_X1 U14 ( .B1(n226), .B2(n167), .A(n2), .ZN(n186) );
  INV_X1 U15 ( .A(INC_DEC), .ZN(n221) );
  OAI21_X1 U16 ( .B1(n125), .B2(n126), .A(n127), .ZN(n121) );
  NOR2_X1 U17 ( .A1(n128), .A2(n129), .ZN(n127) );
  NAND2_X1 U18 ( .A1(n132), .A2(n133), .ZN(n128) );
  OAI21_X1 U19 ( .B1(n265), .B2(n59), .A(n60), .ZN(n52) );
  INV_X1 U20 ( .A(n61), .ZN(n265) );
  OAI21_X1 U21 ( .B1(n100), .B2(n101), .A(n102), .ZN(n95) );
  NOR2_X1 U22 ( .A1(n103), .A2(n104), .ZN(n102) );
  NAND2_X1 U23 ( .A1(n107), .A2(n108), .ZN(n103) );
  OAI21_X1 U24 ( .B1(n74), .B2(n75), .A(n76), .ZN(n70) );
  NOR2_X1 U25 ( .A1(n77), .A2(n78), .ZN(n76) );
  NAND2_X1 U26 ( .A1(n81), .A2(n82), .ZN(n77) );
  AOI21_X1 U27 ( .B1(n52), .B2(n53), .A(n269), .ZN(n51) );
  INV_X1 U28 ( .A(n55), .ZN(n269) );
  AOI21_X1 U29 ( .B1(n83), .B2(n88), .A(n241), .ZN(n86) );
  INV_X1 U30 ( .A(n80), .ZN(n241) );
  NAND4_X1 U31 ( .A1(n192), .A2(n193), .A3(n17), .A4(n21), .ZN(n167) );
  NAND4_X1 U32 ( .A1(n40), .A2(n36), .A3(n26), .A4(n29), .ZN(n165) );
  NOR2_X1 U33 ( .A1(n165), .A2(n166), .ZN(n159) );
  NOR2_X1 U34 ( .A1(n167), .A2(n168), .ZN(n158) );
  NAND4_X1 U35 ( .A1(n169), .A2(n170), .A3(n171), .A4(n172), .ZN(n168) );
  NAND4_X1 U36 ( .A1(n161), .A2(n162), .A3(n163), .A4(n164), .ZN(n160) );
  NAND2_X1 U37 ( .A1(n74), .A2(n82), .ZN(n93) );
  NAND2_X1 U38 ( .A1(n92), .A2(n81), .ZN(n88) );
  NAND2_X1 U39 ( .A1(n85), .A2(n93), .ZN(n92) );
  NAND2_X1 U40 ( .A1(n121), .A2(n122), .ZN(n100) );
  NAND2_X1 U41 ( .A1(n150), .A2(n151), .ZN(n125) );
  NAND2_X1 U42 ( .A1(n95), .A2(n96), .ZN(n74) );
  AND2_X1 U43 ( .A1(n68), .A2(n69), .ZN(n59) );
  NAND2_X1 U44 ( .A1(n70), .A2(n71), .ZN(n68) );
  AND4_X1 U45 ( .A1(n28), .A2(n24), .A3(n33), .A4(n38), .ZN(n1) );
  AND4_X1 U46 ( .A1(n190), .A2(n16), .A3(n20), .A4(n191), .ZN(n2) );
  OAI21_X1 U47 ( .B1(n225), .B2(n256), .A(n163), .ZN(n177) );
  INV_X1 U48 ( .A(n170), .ZN(n256) );
  INV_X1 U49 ( .A(n182), .ZN(n225) );
  OAI21_X1 U50 ( .B1(n31), .B2(n232), .A(n33), .ZN(n27) );
  OAI21_X1 U51 ( .B1(n262), .B2(n226), .A(n20), .ZN(n14) );
  INV_X1 U52 ( .A(n21), .ZN(n262) );
  AOI21_X1 U53 ( .B1(n109), .B2(n114), .A(n246), .ZN(n112) );
  INV_X1 U54 ( .A(n106), .ZN(n246) );
  OAI21_X1 U55 ( .B1(n224), .B2(n250), .A(n131), .ZN(n140) );
  INV_X1 U56 ( .A(n134), .ZN(n250) );
  INV_X1 U57 ( .A(n143), .ZN(n224) );
  OAI21_X1 U58 ( .B1(n222), .B2(n237), .A(n46), .ZN(n43) );
  INV_X1 U59 ( .A(n47), .ZN(n237) );
  INV_X1 U60 ( .A(n48), .ZN(n222) );
  NAND2_X1 U61 ( .A1(n229), .A2(n166), .ZN(n39) );
  INV_X1 U62 ( .A(n157), .ZN(n229) );
  NAND2_X1 U63 ( .A1(n125), .A2(n133), .ZN(n147) );
  NAND2_X1 U64 ( .A1(n100), .A2(n108), .ZN(n119) );
  NAND2_X1 U65 ( .A1(n201), .A2(n16), .ZN(n199) );
  NAND2_X1 U66 ( .A1(n14), .A2(n17), .ZN(n201) );
  NAND2_X1 U67 ( .A1(n185), .A2(n164), .ZN(n182) );
  NAND2_X1 U68 ( .A1(n186), .A2(n169), .ZN(n185) );
  NAND2_X1 U69 ( .A1(n146), .A2(n132), .ZN(n143) );
  NAND2_X1 U70 ( .A1(n136), .A2(n147), .ZN(n146) );
  NAND2_X1 U71 ( .A1(n118), .A2(n107), .ZN(n114) );
  NAND2_X1 U72 ( .A1(n111), .A2(n119), .ZN(n118) );
  NAND2_X1 U73 ( .A1(n24), .A2(n25), .ZN(n23) );
  NAND2_X1 U74 ( .A1(n26), .A2(n27), .ZN(n25) );
  NAND2_X1 U75 ( .A1(n162), .A2(n176), .ZN(n175) );
  NAND2_X1 U76 ( .A1(n171), .A2(n177), .ZN(n176) );
  INV_X1 U77 ( .A(n36), .ZN(n232) );
  NAND2_X1 U78 ( .A1(n191), .A2(n198), .ZN(n195) );
  NAND2_X1 U79 ( .A1(n199), .A2(n193), .ZN(n198) );
  NAND2_X1 U80 ( .A1(n105), .A2(n106), .ZN(n104) );
  NAND2_X1 U81 ( .A1(n79), .A2(n80), .ZN(n78) );
  NAND2_X1 U82 ( .A1(n130), .A2(n131), .ZN(n129) );
  INV_X1 U83 ( .A(n33), .ZN(n234) );
  AND2_X1 U84 ( .A1(n37), .A2(n38), .ZN(n31) );
  NAND2_X1 U85 ( .A1(n39), .A2(n40), .ZN(n37) );
  XNOR2_X1 U86 ( .A(n51), .B(n6), .ZN(SUM[31]) );
  XNOR2_X1 U87 ( .A(n86), .B(n4), .ZN(SUM[27]) );
  AND2_X1 U88 ( .A1(n79), .A2(n84), .ZN(n4) );
  NAND4_X1 U89 ( .A1(A[0]), .A2(n66), .A3(n47), .A4(n49), .ZN(n166) );
  NAND2_X1 U90 ( .A1(INC_DEC), .A2(A[8]), .ZN(n20) );
  NAND2_X1 U91 ( .A1(A[5]), .A2(INC_DEC), .ZN(n33) );
  NAND2_X1 U92 ( .A1(A[10]), .A2(INC_DEC), .ZN(n191) );
  NAND2_X1 U93 ( .A1(A[9]), .A2(INC_DEC), .ZN(n16) );
  NAND2_X1 U94 ( .A1(A[6]), .A2(INC_DEC), .ZN(n24) );
  XNOR2_X1 U95 ( .A(n52), .B(n56), .ZN(SUM[30]) );
  NAND2_X1 U96 ( .A1(n55), .A2(n53), .ZN(n56) );
  NAND2_X1 U97 ( .A1(A[4]), .A2(INC_DEC), .ZN(n38) );
  NAND2_X1 U98 ( .A1(n219), .A2(n263), .ZN(n21) );
  INV_X1 U99 ( .A(A[8]), .ZN(n263) );
  NAND2_X1 U100 ( .A1(A[12]), .A2(INC_DEC), .ZN(n164) );
  NAND2_X1 U101 ( .A1(n220), .A2(n261), .ZN(n17) );
  INV_X1 U102 ( .A(A[9]), .ZN(n261) );
  NAND2_X1 U103 ( .A1(n220), .A2(n260), .ZN(n193) );
  INV_X1 U104 ( .A(A[10]), .ZN(n260) );
  NAND2_X1 U105 ( .A1(n220), .A2(n255), .ZN(n171) );
  INV_X1 U106 ( .A(A[14]), .ZN(n255) );
  NAND2_X1 U107 ( .A1(n220), .A2(n258), .ZN(n169) );
  INV_X1 U108 ( .A(A[12]), .ZN(n258) );
  NAND2_X1 U109 ( .A1(n220), .A2(n235), .ZN(n40) );
  INV_X1 U110 ( .A(A[4]), .ZN(n235) );
  NAND2_X1 U111 ( .A1(n219), .A2(n238), .ZN(n47) );
  INV_X1 U112 ( .A(A[2]), .ZN(n238) );
  NAND2_X1 U113 ( .A1(n219), .A2(n231), .ZN(n26) );
  INV_X1 U114 ( .A(A[6]), .ZN(n231) );
  NAND2_X1 U115 ( .A1(n219), .A2(n228), .ZN(n66) );
  INV_X1 U116 ( .A(A[1]), .ZN(n228) );
  NAND2_X1 U117 ( .A1(n219), .A2(n264), .ZN(n29) );
  INV_X1 U118 ( .A(A[7]), .ZN(n264) );
  NAND2_X1 U119 ( .A1(n218), .A2(n254), .ZN(n172) );
  INV_X1 U120 ( .A(A[15]), .ZN(n254) );
  NAND2_X1 U121 ( .A1(n218), .A2(n236), .ZN(n49) );
  INV_X1 U122 ( .A(A[3]), .ZN(n236) );
  NAND2_X1 U123 ( .A1(n218), .A2(n233), .ZN(n36) );
  INV_X1 U124 ( .A(A[5]), .ZN(n233) );
  NAND2_X1 U125 ( .A1(n218), .A2(n259), .ZN(n192) );
  INV_X1 U126 ( .A(A[11]), .ZN(n259) );
  NAND2_X1 U127 ( .A1(A[7]), .A2(INC_DEC), .ZN(n28) );
  NAND2_X1 U128 ( .A1(A[11]), .A2(INC_DEC), .ZN(n190) );
  NAND2_X1 U129 ( .A1(n218), .A2(n257), .ZN(n170) );
  INV_X1 U130 ( .A(A[13]), .ZN(n257) );
  OAI21_X1 U131 ( .B1(n230), .B2(n223), .A(n65), .ZN(n48) );
  INV_X1 U132 ( .A(A[0]), .ZN(n230) );
  INV_X1 U133 ( .A(n66), .ZN(n223) );
  XNOR2_X1 U134 ( .A(n62), .B(n48), .ZN(SUM[2]) );
  NAND2_X1 U135 ( .A1(n47), .A2(n46), .ZN(n62) );
  XNOR2_X1 U136 ( .A(n42), .B(n43), .ZN(SUM[3]) );
  NAND2_X1 U137 ( .A1(n49), .A2(n50), .ZN(n42) );
  XNOR2_X1 U138 ( .A(n41), .B(n39), .ZN(SUM[4]) );
  NAND2_X1 U139 ( .A1(n38), .A2(n40), .ZN(n41) );
  XNOR2_X1 U140 ( .A(n31), .B(n34), .ZN(SUM[5]) );
  NOR2_X1 U141 ( .A1(n234), .A2(n232), .ZN(n34) );
  XNOR2_X1 U142 ( .A(n30), .B(n27), .ZN(SUM[6]) );
  NAND2_X1 U143 ( .A1(n26), .A2(n24), .ZN(n30) );
  XNOR2_X1 U144 ( .A(n22), .B(n23), .ZN(SUM[7]) );
  NAND2_X1 U145 ( .A1(n28), .A2(n29), .ZN(n22) );
  XNOR2_X1 U146 ( .A(n18), .B(n19), .ZN(SUM[8]) );
  NAND2_X1 U147 ( .A1(n20), .A2(n21), .ZN(n18) );
  XNOR2_X1 U148 ( .A(n14), .B(n15), .ZN(SUM[9]) );
  NAND2_X1 U149 ( .A1(n16), .A2(n17), .ZN(n15) );
  XNOR2_X1 U150 ( .A(n188), .B(n186), .ZN(SUM[12]) );
  NAND2_X1 U151 ( .A1(n164), .A2(n169), .ZN(n188) );
  XNOR2_X1 U152 ( .A(n153), .B(n150), .ZN(SUM[16]) );
  NAND2_X1 U153 ( .A1(n133), .A2(n151), .ZN(n153) );
  XNOR2_X1 U154 ( .A(n149), .B(n147), .ZN(SUM[17]) );
  NAND2_X1 U155 ( .A1(n132), .A2(n136), .ZN(n149) );
  XNOR2_X1 U156 ( .A(n139), .B(n140), .ZN(SUM[19]) );
  NAND2_X1 U157 ( .A1(n130), .A2(n135), .ZN(n139) );
  XNOR2_X1 U158 ( .A(n124), .B(n121), .ZN(SUM[20]) );
  NAND2_X1 U159 ( .A1(n108), .A2(n122), .ZN(n124) );
  XNOR2_X1 U160 ( .A(n120), .B(n119), .ZN(SUM[21]) );
  NAND2_X1 U161 ( .A1(n107), .A2(n111), .ZN(n120) );
  XNOR2_X1 U162 ( .A(n112), .B(n5), .ZN(SUM[23]) );
  AND2_X1 U163 ( .A1(n105), .A2(n110), .ZN(n5) );
  XNOR2_X1 U164 ( .A(A[0]), .B(n138), .ZN(SUM[1]) );
  NAND2_X1 U165 ( .A1(n66), .A2(n65), .ZN(n138) );
  XNOR2_X1 U166 ( .A(n174), .B(n175), .ZN(SUM[15]) );
  NAND2_X1 U167 ( .A1(n161), .A2(n172), .ZN(n174) );
  XNOR2_X1 U168 ( .A(n195), .B(n196), .ZN(SUM[11]) );
  NAND2_X1 U169 ( .A1(n190), .A2(n192), .ZN(n196) );
  XNOR2_X1 U170 ( .A(n114), .B(n116), .ZN(SUM[22]) );
  NAND2_X1 U171 ( .A1(n109), .A2(n106), .ZN(n116) );
  XNOR2_X1 U172 ( .A(n95), .B(n98), .ZN(SUM[24]) );
  NAND2_X1 U173 ( .A1(n82), .A2(n96), .ZN(n98) );
  XNOR2_X1 U174 ( .A(n70), .B(n72), .ZN(SUM[28]) );
  NAND2_X1 U175 ( .A1(n69), .A2(n71), .ZN(n72) );
  NAND2_X1 U176 ( .A1(A[22]), .A2(INC_DEC), .ZN(n106) );
  NAND2_X1 U177 ( .A1(A[26]), .A2(INC_DEC), .ZN(n80) );
  NAND2_X1 U178 ( .A1(A[16]), .A2(INC_DEC), .ZN(n133) );
  NAND2_X1 U179 ( .A1(A[20]), .A2(INC_DEC), .ZN(n108) );
  NAND2_X1 U180 ( .A1(A[24]), .A2(INC_DEC), .ZN(n82) );
  NAND2_X1 U181 ( .A1(A[13]), .A2(INC_DEC), .ZN(n163) );
  NAND2_X1 U182 ( .A1(A[18]), .A2(INC_DEC), .ZN(n131) );
  NAND2_X1 U184 ( .A1(A[17]), .A2(INC_DEC), .ZN(n132) );
  NAND2_X1 U185 ( .A1(A[21]), .A2(INC_DEC), .ZN(n107) );
  NAND2_X1 U186 ( .A1(A[25]), .A2(INC_DEC), .ZN(n81) );
  NAND2_X1 U187 ( .A1(A[14]), .A2(INC_DEC), .ZN(n162) );
  NAND2_X1 U188 ( .A1(A[1]), .A2(INC_DEC), .ZN(n65) );
  NAND2_X1 U189 ( .A1(A[2]), .A2(INC_DEC), .ZN(n46) );
  NAND2_X1 U190 ( .A1(n217), .A2(n245), .ZN(n109) );
  INV_X1 U191 ( .A(A[22]), .ZN(n245) );
  NAND2_X1 U192 ( .A1(n217), .A2(n240), .ZN(n83) );
  INV_X1 U193 ( .A(A[26]), .ZN(n240) );
  NAND2_X1 U194 ( .A1(n216), .A2(n268), .ZN(n53) );
  INV_X1 U195 ( .A(A[30]), .ZN(n268) );
  NAND2_X1 U196 ( .A1(n216), .A2(n253), .ZN(n151) );
  INV_X1 U197 ( .A(A[16]), .ZN(n253) );
  NAND2_X1 U198 ( .A1(n217), .A2(n248), .ZN(n122) );
  INV_X1 U199 ( .A(A[20]), .ZN(n248) );
  NAND2_X1 U200 ( .A1(n217), .A2(n243), .ZN(n96) );
  INV_X1 U201 ( .A(A[24]), .ZN(n243) );
  NAND2_X1 U202 ( .A1(n217), .A2(n239), .ZN(n71) );
  INV_X1 U203 ( .A(A[28]), .ZN(n239) );
  NAND2_X1 U204 ( .A1(A[30]), .A2(INC_DEC), .ZN(n55) );
  NAND2_X1 U205 ( .A1(A[19]), .A2(INC_DEC), .ZN(n130) );
  NAND2_X1 U206 ( .A1(A[15]), .A2(INC_DEC), .ZN(n161) );
  NAND2_X1 U207 ( .A1(A[3]), .A2(INC_DEC), .ZN(n50) );
  NAND2_X1 U208 ( .A1(A[29]), .A2(INC_DEC), .ZN(n60) );
  NAND2_X1 U209 ( .A1(A[28]), .A2(INC_DEC), .ZN(n69) );
  NAND2_X1 U210 ( .A1(A[27]), .A2(INC_DEC), .ZN(n79) );
  NAND2_X1 U211 ( .A1(A[23]), .A2(INC_DEC), .ZN(n105) );
  NAND2_X1 U212 ( .A1(n215), .A2(n249), .ZN(n135) );
  INV_X1 U213 ( .A(A[19]), .ZN(n249) );
  NAND2_X1 U214 ( .A1(n216), .A2(n266), .ZN(n61) );
  INV_X1 U215 ( .A(A[29]), .ZN(n266) );
  NAND2_X1 U216 ( .A1(n216), .A2(n267), .ZN(n84) );
  INV_X1 U217 ( .A(A[27]), .ZN(n267) );
  NAND2_X1 U218 ( .A1(n216), .A2(n244), .ZN(n110) );
  INV_X1 U219 ( .A(A[23]), .ZN(n244) );
  XNOR2_X1 U220 ( .A(n179), .B(n177), .ZN(SUM[14]) );
  NAND2_X1 U221 ( .A1(n162), .A2(n171), .ZN(n179) );
  NAND2_X1 U222 ( .A1(n215), .A2(n252), .ZN(n136) );
  INV_X1 U223 ( .A(A[17]), .ZN(n252) );
  NAND2_X1 U224 ( .A1(n215), .A2(n251), .ZN(n134) );
  INV_X1 U226 ( .A(A[18]), .ZN(n251) );
  NAND2_X1 U228 ( .A1(n215), .A2(n247), .ZN(n111) );
  INV_X1 U229 ( .A(A[21]), .ZN(n247) );
  NAND2_X1 U231 ( .A1(n215), .A2(n242), .ZN(n85) );
  INV_X1 U232 ( .A(A[25]), .ZN(n242) );
  XNOR2_X1 U233 ( .A(n94), .B(n93), .ZN(SUM[25]) );
  NAND2_X1 U234 ( .A1(n81), .A2(n85), .ZN(n94) );
  XNOR2_X1 U235 ( .A(n200), .B(n199), .ZN(SUM[10]) );
  NAND2_X1 U236 ( .A1(n191), .A2(n193), .ZN(n200) );
  XNOR2_X1 U237 ( .A(n184), .B(n182), .ZN(SUM[13]) );
  NAND2_X1 U238 ( .A1(n163), .A2(n170), .ZN(n184) );
  XNOR2_X1 U239 ( .A(n145), .B(n143), .ZN(SUM[18]) );
  NAND2_X1 U240 ( .A1(n131), .A2(n134), .ZN(n145) );
  XNOR2_X1 U241 ( .A(n88), .B(n90), .ZN(SUM[26]) );
  NAND2_X1 U242 ( .A1(n83), .A2(n80), .ZN(n90) );
  XNOR2_X1 U243 ( .A(n59), .B(n3), .ZN(SUM[29]) );
  AND2_X1 U245 ( .A1(n60), .A2(n61), .ZN(n3) );
endmodule


module windowed_register_file_M8_N4_N_bit64_W2 ( CALL, RETURN_signal, CLK, 
        RESET, ENABLE, RD_CPU, WR_CPU, Wait_signal, ADDR_WRCPU, ADDR_RDCPU, 
        DATAIN_CPU, DATAOUT_CPU, RD_WR_MEM, DATAIN_MEM, DATAOUT_MEM );
  input [4:0] ADDR_WRCPU;
  input [4:0] ADDR_RDCPU;
  input [63:0] DATAIN_CPU;
  output [63:0] DATAOUT_CPU;
  input [63:0] DATAIN_MEM;
  output [63:0] DATAOUT_MEM;
  input CALL, RETURN_signal, CLK, RESET, ENABLE, RD_CPU, WR_CPU;
  output Wait_signal, RD_WR_MEM;
  wire   full, count_wait, RD_MEM, start, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N212, N213, N264,
         N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N351, N352,
         N353, \U3/U1/Z_0 , n156, n157, n158, n159, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n196, n197, n198, n200,
         n202, n204, n205, n206, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n248, n282, n283, n290, n387, n389, n390, n392, n393,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n431, n565, n566, n567, n568, n570, n571, n572, n573,
         n576, n577, n578, n579, n581, n582, n583, n588, n589, n621, n675,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n912;
  wire   [4:0] ADDRESS_WRITE;
  wire   [4:0] ADDRESS_READ;
  wire   [4:0] ADDRESS_COUNT;
  wire   [63:0] DATA_WRITE;
  wire   [4:0] swp;
  wire   [4:0] cwp;
  wire   [31:0] canrestore;
  wire   [31:0] cansave;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign \U3/U1/Z_0  = CALL;

  DFF_X1 \canrestore_reg[28]  ( .D(n409), .CK(CLK), .Q(canrestore[28]), .QN(
        n815) );
  DFF_X1 \canrestore_reg[29]  ( .D(n408), .CK(CLK), .Q(canrestore[29]), .QN(
        n814) );
  DFF_X1 \canrestore_reg[26]  ( .D(n411), .CK(CLK), .Q(canrestore[26]), .QN(
        n588) );
  DFF_X1 \canrestore_reg[27]  ( .D(n410), .CK(CLK), .Q(canrestore[27]), .QN(
        n573) );
  DFF_X1 \canrestore_reg[30]  ( .D(n406), .CK(CLK), .Q(canrestore[30]), .QN(
        n813) );
  DFF_X1 \canrestore_reg[31]  ( .D(n405), .CK(CLK), .Q(canrestore[31]), .QN(
        n389) );
  XOR2_X1 U667 ( .A(n197), .B(n725), .Z(n772) );
  NAND3_X1 U668 ( .A1(n775), .A2(cansave[0]), .A3(n776), .ZN(n773) );
  XOR2_X1 U669 ( .A(cansave[1]), .B(\U3/U1/Z_0 ), .Z(n776) );
  NAND3_X1 U670 ( .A1(n731), .A2(n771), .A3(n780), .ZN(n779) );
  XOR2_X1 U671 ( .A(n193), .B(n157), .Z(n787) );
  XOR2_X1 U672 ( .A(n192), .B(n158), .Z(n785) );
  XOR2_X1 U673 ( .A(swp[4]), .B(n788), .Z(n783) );
  XOR2_X1 U674 ( .A(n621), .B(cwp[3]), .Z(n789) );
  NAND3_X1 U675 ( .A1(n872), .A2(cwp[3]), .A3(swp[3]), .ZN(n782) );
  NAND3_X1 U676 ( .A1(n794), .A2(n795), .A3(n796), .ZN(n793) );
  NAND3_X1 U677 ( .A1(n775), .A2(cansave[0]), .A3(n196), .ZN(n731) );
  NAND3_X1 U678 ( .A1(n775), .A2(cansave[1]), .A3(n197), .ZN(n780) );
  NAND3_X1 U679 ( .A1(cansave[1]), .A2(cansave[0]), .A3(n775), .ZN(n770) );
  NAND3_X1 U680 ( .A1(n174), .A2(n173), .A3(n175), .ZN(n811) );
  register_file_NBIT64_NREG32 WRF ( .CLK(CLK), .RESET(RESET), .ENABLE(ENABLE), 
        .RD1(RD_CPU), .RD2(RD_MEM), .WR(n875), .ADD_WR(ADDRESS_WRITE), 
        .ADD_RD1(ADDRESS_READ), .ADD_RD2(ADDRESS_COUNT), .DATAIN(DATA_WRITE), 
        .OUT1(DATAOUT_CPU), .OUT2(DATAOUT_MEM) );
  address_conversion_M8_N4_N_bit64_F3 add_con ( .spill_fill_count(full), 
        .wait_count(count_wait), .start_write(start), .clck(CLK), 
        .address_input_1(ADDR_RDCPU), .address_input_3(ADDR_WRCPU), 
        .address_output_1(ADDRESS_READ), .address_output_2(ADDRESS_COUNT), 
        .address_output_3(ADDRESS_WRITE), .swp({swp[4:3], N353, N352, N351}), 
        .cwp({cwp[4:3], N213, N212, cwp[0]}) );
  MUX21_generic_N64 DATA_multiplexer_write ( .A(DATAIN_MEM), .B(DATAIN_CPU), 
        .sel(Wait_signal), .Y(DATA_WRITE) );
  windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_2 r47 ( .A(canrestore), 
        .INC_DEC(n860), .SUM({N295, N294, N293, N292, N291, N290, N289, N288, 
        N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, 
        N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264}) );
  windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_3 r48 ( .A(cansave), 
        .INC_DEC(\U3/U1/Z_0 ), .SUM({N84, N83, N82, N81, N80, N79, N78, N77, 
        N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, 
        N62, N61, N60, N59, N58, N57, N56, N55, N54, SYNOPSYS_UNCONNECTED__0})
         );
  DFFRS_X1 \swp_reg[0]  ( .D(n283), .CK(n675), .RN(n431), .SN(n206), .Q(N351), 
        .QN(n191) );
  DFFRS_X1 \swp_reg[1]  ( .D(n209), .CK(n675), .RN(n395), .SN(n200), .Q(N352), 
        .QN(n192) );
  DFFRS_X1 \swp_reg[2]  ( .D(n208), .CK(n675), .RN(n396), .SN(n198), .Q(N353), 
        .QN(n193) );
  DFFRS_X1 \swp_reg[4]  ( .D(n211), .CK(n675), .RN(n205), .SN(n204), .Q(swp[4]) );
  DFFRS_X1 \swp_reg[3]  ( .D(n210), .CK(n675), .RN(n397), .SN(n202), .Q(swp[3]), .QN(n290) );
  DFF_X1 \cansave_reg[1]  ( .D(n826), .CK(CLK), .Q(cansave[1]), .QN(n196) );
  DFF_X1 \cansave_reg[0]  ( .D(n248), .CK(CLK), .Q(cansave[0]), .QN(n197) );
  DFF_X1 \canrestore_reg[0]  ( .D(n429), .CK(CLK), .Q(canrestore[0]), .QN(n579) );
  DFF_X1 \cansave_reg[6]  ( .D(n856), .CK(CLK), .Q(cansave[6]), .QN(n185) );
  DFF_X1 \cansave_reg[5]  ( .D(n855), .CK(CLK), .Q(cansave[5]), .QN(n186) );
  DFF_X1 \cansave_reg[4]  ( .D(n854), .CK(CLK), .Q(cansave[4]), .QN(n187) );
  DFF_X1 \cansave_reg[3]  ( .D(n853), .CK(CLK), .Q(cansave[3]), .QN(n188) );
  DFF_X1 \cansave_reg[2]  ( .D(n852), .CK(CLK), .Q(cansave[2]), .QN(n189) );
  DFF_X1 \cwp_reg[4]  ( .D(n825), .CK(CLK), .Q(cwp[4]), .QN(n621) );
  DFF_X1 \cansave_reg[20]  ( .D(n828), .CK(CLK), .Q(cansave[20]), .QN(n171) );
  DFF_X1 \cwp_reg[3]  ( .D(n213), .CK(CLK), .Q(cwp[3]), .QN(n156) );
  DFF_X1 \cansave_reg[21]  ( .D(n829), .CK(CLK), .Q(cansave[21]), .QN(n170) );
  DFF_X1 \cansave_reg[18]  ( .D(n850), .CK(CLK), .Q(cansave[18]), .QN(n173) );
  DFF_X1 \cansave_reg[17]  ( .D(n849), .CK(CLK), .Q(cansave[17]), .QN(n174) );
  DFF_X1 \cansave_reg[16]  ( .D(n848), .CK(CLK), .Q(cansave[16]), .QN(n175) );
  DFF_X1 \cansave_reg[12]  ( .D(n844), .CK(CLK), .Q(cansave[12]), .QN(n179) );
  DFF_X1 \cansave_reg[9]  ( .D(n841), .CK(CLK), .Q(cansave[9]), .QN(n182) );
  DFF_X1 \cansave_reg[8]  ( .D(n840), .CK(CLK), .Q(cansave[8]), .QN(n183) );
  DFF_X1 \cansave_reg[7]  ( .D(n839), .CK(CLK), .Q(cansave[7]), .QN(n184) );
  DFF_X1 \cansave_reg[13]  ( .D(n845), .CK(CLK), .Q(cansave[13]), .QN(n178) );
  DFF_X1 \cansave_reg[10]  ( .D(n842), .CK(CLK), .Q(cansave[10]), .QN(n181) );
  DFF_X1 \cwp_reg[2]  ( .D(n214), .CK(CLK), .Q(N213), .QN(n157) );
  DFF_X1 \cwp_reg[1]  ( .D(n215), .CK(CLK), .Q(N212), .QN(n158) );
  DFF_X1 \cwp_reg[0]  ( .D(n216), .CK(CLK), .Q(cwp[0]), .QN(n159) );
  DFF_X1 \cansave_reg[24]  ( .D(n832), .CK(CLK), .Q(cansave[24]), .QN(n167) );
  DFF_X1 \cansave_reg[19]  ( .D(n827), .CK(CLK), .Q(cansave[19]), .QN(n172) );
  DFF_X1 \cansave_reg[11]  ( .D(n843), .CK(CLK), .Q(cansave[11]), .QN(n180) );
  DFF_X1 \cansave_reg[22]  ( .D(n830), .CK(CLK), .Q(cansave[22]), .QN(n169) );
  DFF_X1 \cansave_reg[23]  ( .D(n831), .CK(CLK), .Q(cansave[23]), .QN(n168) );
  DFF_X1 \cansave_reg[14]  ( .D(n846), .CK(CLK), .Q(cansave[14]), .QN(n177) );
  DFF_X1 \cansave_reg[25]  ( .D(n833), .CK(CLK), .Q(cansave[25]), .QN(n166) );
  DFF_X1 \cansave_reg[28]  ( .D(n836), .CK(CLK), .Q(cansave[28]), .QN(n163) );
  DFF_X1 \canrestore_reg[2]  ( .D(n407), .CK(CLK), .Q(canrestore[2]), .QN(n568) );
  DFF_X1 \cansave_reg[15]  ( .D(n847), .CK(CLK), .Q(cansave[15]), .QN(n176) );
  DFF_X1 \canrestore_reg[1]  ( .D(n418), .CK(CLK), .Q(canrestore[1]), .QN(n589) );
  DFF_X1 \canrestore_reg[3]  ( .D(n404), .CK(CLK), .Q(canrestore[3]), .QN(n392) );
  DFF_X1 \canrestore_reg[4]  ( .D(n403), .CK(CLK), .Q(canrestore[4]), .QN(n393) );
  DFF_X1 \cansave_reg[26]  ( .D(n834), .CK(CLK), .Q(cansave[26]), .QN(n165) );
  DFF_X1 \cansave_reg[29]  ( .D(n837), .CK(CLK), .Q(cansave[29]), .QN(n162) );
  DFF_X1 \cansave_reg[27]  ( .D(n835), .CK(CLK), .Q(cansave[27]), .QN(n164) );
  DFF_X1 SPILL_reg ( .D(n212), .CK(CLK), .Q(n859), .QN(n675) );
  DFF_X1 FILL_reg ( .D(n282), .CK(CLK), .Q(n387), .QN(RD_WR_MEM) );
  DFF_X1 \canrestore_reg[5]  ( .D(n402), .CK(CLK), .Q(canrestore[5]), .QN(n572) );
  DFF_X1 \cansave_reg[30]  ( .D(n838), .CK(CLK), .Q(cansave[30]), .QN(n161) );
  DFF_X1 \canrestore_reg[8]  ( .D(n399), .CK(CLK), .Q(canrestore[8]), .QN(n566) );
  DFF_X1 \canrestore_reg[16]  ( .D(n422), .CK(CLK), .Q(canrestore[16]), .QN(
        n823) );
  DFF_X1 \cansave_reg[31]  ( .D(n851), .CK(CLK), .Q(cansave[31]), .QN(n190) );
  DFF_X1 \canrestore_reg[6]  ( .D(n401), .CK(CLK), .Q(canrestore[6]), .QN(n567) );
  DFF_X1 \canrestore_reg[12]  ( .D(n426), .CK(CLK), .Q(canrestore[12]), .QN(
        n581) );
  DFF_X1 \canrestore_reg[9]  ( .D(n398), .CK(CLK), .Q(canrestore[9]), .QN(n390) );
  DFF_X1 \canrestore_reg[7]  ( .D(n400), .CK(CLK), .Q(canrestore[7]), .QN(n565) );
  DFF_X1 \canrestore_reg[17]  ( .D(n421), .CK(CLK), .Q(canrestore[17]), .QN(
        n822) );
  DFF_X1 \canrestore_reg[13]  ( .D(n425), .CK(CLK), .Q(canrestore[13]), .QN(
        n582) );
  DFF_X1 \canrestore_reg[10]  ( .D(n428), .CK(CLK), .Q(canrestore[10]), .QN(
        n577) );
  DFF_X1 \canrestore_reg[20]  ( .D(n417), .CK(CLK), .Q(canrestore[20]), .QN(
        n819) );
  DFF_X1 \canrestore_reg[18]  ( .D(n420), .CK(CLK), .Q(canrestore[18]), .QN(
        n821) );
  DFF_X1 \canrestore_reg[11]  ( .D(n427), .CK(CLK), .Q(canrestore[11]), .QN(
        n578) );
  DFF_X1 \canrestore_reg[14]  ( .D(n424), .CK(CLK), .Q(canrestore[14]), .QN(
        n583) );
  DFF_X1 \canrestore_reg[21]  ( .D(n416), .CK(CLK), .Q(canrestore[21]), .QN(
        n818) );
  DFF_X1 \canrestore_reg[19]  ( .D(n419), .CK(CLK), .Q(canrestore[19]), .QN(
        n820) );
  DFF_X1 \canrestore_reg[24]  ( .D(n413), .CK(CLK), .Q(canrestore[24]), .QN(
        n570) );
  DFF_X1 \canrestore_reg[15]  ( .D(n423), .CK(CLK), .Q(canrestore[15]), .QN(
        n576) );
  DFF_X1 \canrestore_reg[22]  ( .D(n415), .CK(CLK), .Q(canrestore[22]), .QN(
        n817) );
  DFF_X1 \canrestore_reg[23]  ( .D(n414), .CK(CLK), .Q(canrestore[23]), .QN(
        n816) );
  DFF_X1 \canrestore_reg[25]  ( .D(n412), .CK(CLK), .Q(canrestore[25]), .QN(
        n571) );
  AND2_X1 U681 ( .A1(n725), .A2(n863), .ZN(n774) );
  INV_X1 U682 ( .A(n871), .ZN(n865) );
  INV_X1 U683 ( .A(n871), .ZN(n864) );
  INV_X1 U684 ( .A(n871), .ZN(n866) );
  INV_X1 U685 ( .A(n871), .ZN(n867) );
  INV_X1 U686 ( .A(n871), .ZN(n868) );
  INV_X1 U687 ( .A(n871), .ZN(n869) );
  INV_X1 U688 ( .A(n871), .ZN(n870) );
  BUF_X1 U689 ( .A(n732), .Z(n862) );
  BUF_X1 U690 ( .A(n732), .Z(n861) );
  BUF_X1 U691 ( .A(n732), .Z(n863) );
  NOR2_X1 U692 ( .A1(n858), .A2(n878), .ZN(n767) );
  INV_X1 U693 ( .A(n770), .ZN(n878) );
  NAND2_X1 U694 ( .A1(n725), .A2(n773), .ZN(n732) );
  OR2_X1 U695 ( .A1(n777), .A2(\U3/U1/Z_0 ), .ZN(n858) );
  AOI21_X1 U696 ( .B1(n872), .B2(n777), .A(Wait_signal), .ZN(n725) );
  NOR2_X1 U697 ( .A1(n872), .A2(n731), .ZN(n729) );
  NAND2_X1 U698 ( .A1(n778), .A2(n873), .ZN(n212) );
  INV_X1 U699 ( .A(n765), .ZN(n873) );
  OAI211_X1 U700 ( .C1(RD_WR_MEM), .C2(n874), .A(n779), .B(\U3/U1/Z_0 ), .ZN(
        n778) );
  NAND2_X1 U701 ( .A1(n878), .A2(n872), .ZN(n728) );
  NOR2_X1 U702 ( .A1(RD_WR_MEM), .A2(n878), .ZN(n803) );
  INV_X1 U703 ( .A(n780), .ZN(n879) );
  NAND2_X1 U704 ( .A1(n803), .A2(n912), .ZN(n205) );
  INV_X1 U705 ( .A(n802), .ZN(n912) );
  NOR2_X1 U706 ( .A1(n879), .A2(n802), .ZN(n211) );
  NOR4_X1 U707 ( .A1(n808), .A2(n809), .A3(n810), .A4(n811), .ZN(n807) );
  NAND4_X1 U708 ( .A1(n164), .A2(n163), .A3(n162), .A4(n161), .ZN(n808) );
  NAND4_X1 U709 ( .A1(n168), .A2(n167), .A3(n166), .A4(n165), .ZN(n809) );
  AOI22_X1 U710 ( .A1(n767), .A2(n727), .B1(n621), .B2(\U3/U1/Z_0 ), .ZN(n788)
         );
  OAI211_X1 U711 ( .C1(n792), .C2(n793), .A(RETURN_signal), .B(n389), .ZN(n777) );
  NAND4_X1 U712 ( .A1(n798), .A2(n799), .A3(n800), .A4(n801), .ZN(n792) );
  AND4_X1 U713 ( .A1(n577), .A2(n578), .A3(n579), .A4(n581), .ZN(n798) );
  OAI21_X1 U714 ( .B1(n565), .B2(n870), .A(n762), .ZN(n400) );
  NAND2_X1 U715 ( .A1(N271), .A2(n864), .ZN(n762) );
  OAI21_X1 U716 ( .B1(n572), .B2(n870), .A(n760), .ZN(n402) );
  NAND2_X1 U717 ( .A1(N269), .A2(n864), .ZN(n760) );
  XNOR2_X1 U718 ( .A(n789), .B(n767), .ZN(n727) );
  OAI22_X1 U719 ( .A1(n190), .A2(n868), .B1(n863), .B2(n884), .ZN(n851) );
  INV_X1 U720 ( .A(N84), .ZN(n884) );
  OAI22_X1 U721 ( .A1(n164), .A2(n867), .B1(n861), .B2(n887), .ZN(n835) );
  INV_X1 U722 ( .A(N80), .ZN(n887) );
  OAI22_X1 U723 ( .A1(RD_WR_MEM), .A2(n874), .B1(n765), .B2(n766), .ZN(n282)
         );
  AOI21_X1 U724 ( .B1(n876), .B2(n767), .A(n768), .ZN(n766) );
  AND4_X1 U725 ( .A1(n769), .A2(swp[4]), .A3(n191), .A4(n290), .ZN(n768) );
  INV_X1 U726 ( .A(n771), .ZN(n876) );
  NAND4_X1 U727 ( .A1(n781), .A2(n782), .A3(n783), .A4(n784), .ZN(n771) );
  NOR3_X1 U728 ( .A1(n785), .A2(n786), .A3(n787), .ZN(n784) );
  OAI21_X1 U729 ( .B1(n156), .B2(\U3/U1/Z_0 ), .A(n790), .ZN(n781) );
  OAI22_X1 U730 ( .A1(n161), .A2(n867), .B1(n861), .B2(n883), .ZN(n838) );
  INV_X1 U731 ( .A(N83), .ZN(n883) );
  NAND4_X1 U732 ( .A1(n172), .A2(n171), .A3(n170), .A4(n169), .ZN(n810) );
  OAI21_X1 U733 ( .B1(n576), .B2(n869), .A(n739), .ZN(n423) );
  NAND2_X1 U734 ( .A1(N279), .A2(n866), .ZN(n739) );
  OAI21_X1 U735 ( .B1(n583), .B2(n869), .A(n738), .ZN(n424) );
  NAND2_X1 U736 ( .A1(N278), .A2(n866), .ZN(n738) );
  OAI21_X1 U737 ( .B1(n578), .B2(n869), .A(n735), .ZN(n427) );
  NAND2_X1 U738 ( .A1(N275), .A2(n866), .ZN(n735) );
  OAI21_X1 U739 ( .B1(n577), .B2(n869), .A(n734), .ZN(n428) );
  NAND2_X1 U740 ( .A1(N274), .A2(n864), .ZN(n734) );
  OAI21_X1 U741 ( .B1(n582), .B2(n869), .A(n737), .ZN(n425) );
  NAND2_X1 U742 ( .A1(N277), .A2(n865), .ZN(n737) );
  OAI21_X1 U743 ( .B1(n581), .B2(n869), .A(n736), .ZN(n426) );
  NAND2_X1 U744 ( .A1(N276), .A2(n866), .ZN(n736) );
  OAI21_X1 U745 ( .B1(n389), .B2(n870), .A(n757), .ZN(n405) );
  NAND2_X1 U746 ( .A1(N295), .A2(n864), .ZN(n757) );
  OAI21_X1 U747 ( .B1(n813), .B2(n870), .A(n756), .ZN(n406) );
  NAND2_X1 U748 ( .A1(N294), .A2(n865), .ZN(n756) );
  OAI21_X1 U749 ( .B1(n573), .B2(n870), .A(n752), .ZN(n410) );
  NAND2_X1 U750 ( .A1(N291), .A2(n864), .ZN(n752) );
  OAI21_X1 U751 ( .B1(n588), .B2(n870), .A(n751), .ZN(n411) );
  NAND2_X1 U752 ( .A1(N290), .A2(n865), .ZN(n751) );
  OAI21_X1 U753 ( .B1(n814), .B2(n870), .A(n754), .ZN(n408) );
  NAND2_X1 U754 ( .A1(N293), .A2(n865), .ZN(n754) );
  OAI21_X1 U755 ( .B1(n816), .B2(n869), .A(n748), .ZN(n414) );
  NAND2_X1 U756 ( .A1(N287), .A2(n865), .ZN(n748) );
  OAI21_X1 U757 ( .B1(n571), .B2(n867), .A(n750), .ZN(n412) );
  NAND2_X1 U758 ( .A1(N289), .A2(n865), .ZN(n750) );
  OAI21_X1 U759 ( .B1(n815), .B2(n870), .A(n753), .ZN(n409) );
  NAND2_X1 U760 ( .A1(N292), .A2(n865), .ZN(n753) );
  OAI21_X1 U761 ( .B1(n817), .B2(n868), .A(n747), .ZN(n415) );
  NAND2_X1 U762 ( .A1(N286), .A2(n865), .ZN(n747) );
  OAI21_X1 U763 ( .B1(n820), .B2(n870), .A(n743), .ZN(n419) );
  NAND2_X1 U764 ( .A1(N283), .A2(n866), .ZN(n743) );
  OAI21_X1 U765 ( .B1(n818), .B2(n869), .A(n746), .ZN(n416) );
  NAND2_X1 U766 ( .A1(N285), .A2(n865), .ZN(n746) );
  OAI21_X1 U767 ( .B1(n570), .B2(n867), .A(n749), .ZN(n413) );
  NAND2_X1 U768 ( .A1(N288), .A2(n865), .ZN(n749) );
  OAI21_X1 U769 ( .B1(n821), .B2(n868), .A(n742), .ZN(n420) );
  NAND2_X1 U770 ( .A1(N282), .A2(n864), .ZN(n742) );
  OAI21_X1 U771 ( .B1(n390), .B2(n870), .A(n764), .ZN(n398) );
  NAND2_X1 U772 ( .A1(N273), .A2(n864), .ZN(n764) );
  OAI21_X1 U773 ( .B1(n822), .B2(n870), .A(n741), .ZN(n421) );
  NAND2_X1 U774 ( .A1(N281), .A2(n866), .ZN(n741) );
  OAI21_X1 U775 ( .B1(n819), .B2(n869), .A(n745), .ZN(n417) );
  NAND2_X1 U776 ( .A1(N284), .A2(n865), .ZN(n745) );
  OAI21_X1 U777 ( .B1(n567), .B2(n870), .A(n761), .ZN(n401) );
  NAND2_X1 U778 ( .A1(N270), .A2(n864), .ZN(n761) );
  OAI21_X1 U779 ( .B1(n823), .B2(n867), .A(n740), .ZN(n422) );
  NAND2_X1 U780 ( .A1(N280), .A2(n866), .ZN(n740) );
  OAI21_X1 U781 ( .B1(n566), .B2(n866), .A(n763), .ZN(n399) );
  NAND2_X1 U782 ( .A1(N272), .A2(n864), .ZN(n763) );
  AND4_X1 U783 ( .A1(n804), .A2(n805), .A3(n806), .A4(n807), .ZN(n775) );
  AND4_X1 U784 ( .A1(n180), .A2(n181), .A3(n182), .A4(n183), .ZN(n804) );
  AND4_X1 U785 ( .A1(n176), .A2(n177), .A3(n178), .A4(n179), .ZN(n805) );
  AND4_X1 U786 ( .A1(n812), .A2(n190), .A3(n188), .A4(n189), .ZN(n806) );
  AND4_X1 U787 ( .A1(n390), .A2(n392), .A3(n393), .A4(n565), .ZN(n801) );
  AND4_X1 U788 ( .A1(n566), .A2(n567), .A3(n568), .A4(n570), .ZN(n800) );
  AND4_X1 U789 ( .A1(n571), .A2(n572), .A3(n573), .A4(n576), .ZN(n799) );
  AND4_X1 U790 ( .A1(n797), .A2(n813), .A3(n815), .A4(n814), .ZN(n796) );
  AND4_X1 U791 ( .A1(n816), .A2(n817), .A3(n818), .A4(n819), .ZN(n797) );
  AND4_X1 U792 ( .A1(n582), .A2(n583), .A3(n588), .A4(n589), .ZN(n795) );
  AND4_X1 U793 ( .A1(n823), .A2(n822), .A3(n821), .A4(n820), .ZN(n794) );
  NOR4_X1 U794 ( .A1(n770), .A2(n858), .A3(N352), .A4(N353), .ZN(n769) );
  OAI21_X1 U795 ( .B1(n393), .B2(n870), .A(n759), .ZN(n403) );
  NAND2_X1 U796 ( .A1(N268), .A2(n864), .ZN(n759) );
  OAI21_X1 U797 ( .B1(n392), .B2(n870), .A(n758), .ZN(n404) );
  NAND2_X1 U798 ( .A1(N267), .A2(n864), .ZN(n758) );
  OAI22_X1 U799 ( .A1(n189), .A2(n868), .B1(n863), .B2(n882), .ZN(n852) );
  INV_X1 U800 ( .A(N55), .ZN(n882) );
  OAI22_X1 U801 ( .A1(n188), .A2(n868), .B1(n863), .B2(n881), .ZN(n853) );
  INV_X1 U802 ( .A(N56), .ZN(n881) );
  OAI22_X1 U803 ( .A1(n187), .A2(n868), .B1(n863), .B2(n910), .ZN(n854) );
  INV_X1 U804 ( .A(N57), .ZN(n910) );
  OAI22_X1 U805 ( .A1(n186), .A2(n869), .B1(n863), .B2(n909), .ZN(n855) );
  INV_X1 U806 ( .A(N58), .ZN(n909) );
  OAI22_X1 U807 ( .A1(n185), .A2(n869), .B1(n863), .B2(n908), .ZN(n856) );
  INV_X1 U808 ( .A(N59), .ZN(n908) );
  OAI22_X1 U809 ( .A1(n184), .A2(n867), .B1(n862), .B2(n907), .ZN(n839) );
  INV_X1 U810 ( .A(N60), .ZN(n907) );
  OAI22_X1 U811 ( .A1(n183), .A2(n867), .B1(n862), .B2(n906), .ZN(n840) );
  INV_X1 U812 ( .A(N61), .ZN(n906) );
  OAI22_X1 U813 ( .A1(n182), .A2(n867), .B1(n862), .B2(n901), .ZN(n841) );
  INV_X1 U814 ( .A(N62), .ZN(n901) );
  OAI22_X1 U815 ( .A1(n179), .A2(n868), .B1(n862), .B2(n905), .ZN(n844) );
  INV_X1 U816 ( .A(N65), .ZN(n905) );
  OAI22_X1 U817 ( .A1(n175), .A2(n869), .B1(n862), .B2(n898), .ZN(n848) );
  INV_X1 U818 ( .A(N69), .ZN(n898) );
  OAI22_X1 U819 ( .A1(n174), .A2(n868), .B1(n862), .B2(n897), .ZN(n849) );
  INV_X1 U820 ( .A(N70), .ZN(n897) );
  OAI22_X1 U821 ( .A1(n172), .A2(n867), .B1(n862), .B2(n895), .ZN(n827) );
  INV_X1 U822 ( .A(N72), .ZN(n895) );
  OAI22_X1 U823 ( .A1(n171), .A2(n866), .B1(n861), .B2(n894), .ZN(n828) );
  INV_X1 U824 ( .A(N73), .ZN(n894) );
  OAI22_X1 U825 ( .A1(n170), .A2(n867), .B1(n861), .B2(n893), .ZN(n829) );
  INV_X1 U826 ( .A(N74), .ZN(n893) );
  OAI22_X1 U827 ( .A1(n168), .A2(n867), .B1(n861), .B2(n891), .ZN(n831) );
  INV_X1 U828 ( .A(N76), .ZN(n891) );
  OAI22_X1 U829 ( .A1(n621), .A2(n866), .B1(n726), .B2(n871), .ZN(n825) );
  AOI21_X1 U830 ( .B1(n727), .B2(n880), .A(n877), .ZN(n726) );
  INV_X1 U831 ( .A(n729), .ZN(n880) );
  INV_X1 U832 ( .A(n728), .ZN(n877) );
  OAI22_X1 U833 ( .A1(n196), .A2(n866), .B1(n730), .B2(n871), .ZN(n826) );
  AOI21_X1 U834 ( .B1(N54), .B2(n728), .A(n729), .ZN(n730) );
  OAI22_X1 U835 ( .A1(n156), .A2(n869), .B1(cwp[3]), .B2(n861), .ZN(n213) );
  NOR2_X1 U836 ( .A1(n874), .A2(n675), .ZN(n765) );
  NAND2_X1 U837 ( .A1(n675), .A2(RD_WR_MEM), .ZN(full) );
  XNOR2_X1 U838 ( .A(N351), .B(n159), .ZN(n786) );
  XNOR2_X1 U839 ( .A(swp[3]), .B(n791), .ZN(n790) );
  NOR2_X1 U840 ( .A1(n767), .A2(cwp[3]), .ZN(n791) );
  OAI22_X1 U841 ( .A1(n176), .A2(n868), .B1(n862), .B2(n902), .ZN(n847) );
  INV_X1 U842 ( .A(N68), .ZN(n902) );
  OAI22_X1 U843 ( .A1(n180), .A2(n869), .B1(n862), .B2(n899), .ZN(n843) );
  INV_X1 U844 ( .A(N64), .ZN(n899) );
  OAI22_X1 U845 ( .A1(n169), .A2(n866), .B1(n861), .B2(n892), .ZN(n830) );
  INV_X1 U846 ( .A(N75), .ZN(n892) );
  OAI22_X1 U847 ( .A1(n167), .A2(n867), .B1(n861), .B2(n890), .ZN(n832) );
  INV_X1 U848 ( .A(N77), .ZN(n890) );
  OAI22_X1 U849 ( .A1(n163), .A2(n867), .B1(n861), .B2(n886), .ZN(n836) );
  INV_X1 U850 ( .A(N81), .ZN(n886) );
  INV_X1 U851 ( .A(n724), .ZN(n875) );
  AOI21_X1 U852 ( .B1(start), .B2(n387), .A(WR_CPU), .ZN(n724) );
  AND2_X1 U853 ( .A1(count_wait), .A2(full), .ZN(Wait_signal) );
  OAI21_X1 U854 ( .B1(n579), .B2(n869), .A(n733), .ZN(n429) );
  NAND2_X1 U855 ( .A1(N264), .A2(n864), .ZN(n733) );
  OAI21_X1 U856 ( .B1(n568), .B2(n870), .A(n755), .ZN(n407) );
  NAND2_X1 U857 ( .A1(N266), .A2(n865), .ZN(n755) );
  OAI21_X1 U858 ( .B1(n589), .B2(n868), .A(n744), .ZN(n418) );
  NAND2_X1 U859 ( .A1(N265), .A2(n866), .ZN(n744) );
  NOR2_X1 U860 ( .A1(n158), .A2(n774), .ZN(n215) );
  NOR2_X1 U861 ( .A1(n159), .A2(n774), .ZN(n216) );
  NOR2_X1 U862 ( .A1(n157), .A2(n774), .ZN(n214) );
  NAND2_X1 U863 ( .A1(n772), .A2(n773), .ZN(n248) );
  AND2_X1 U864 ( .A1(n859), .A2(start), .ZN(RD_MEM) );
  AND4_X1 U865 ( .A1(n187), .A2(n186), .A3(n185), .A4(n184), .ZN(n812) );
  OAI22_X1 U866 ( .A1(n177), .A2(n868), .B1(n862), .B2(n903), .ZN(n846) );
  INV_X1 U867 ( .A(N67), .ZN(n903) );
  OAI22_X1 U868 ( .A1(n166), .A2(n867), .B1(n861), .B2(n889), .ZN(n833) );
  INV_X1 U869 ( .A(N78), .ZN(n889) );
  OAI22_X1 U870 ( .A1(n181), .A2(n868), .B1(n862), .B2(n900), .ZN(n842) );
  INV_X1 U871 ( .A(N63), .ZN(n900) );
  OAI22_X1 U872 ( .A1(n178), .A2(n868), .B1(n862), .B2(n904), .ZN(n845) );
  INV_X1 U873 ( .A(N66), .ZN(n904) );
  OAI22_X1 U874 ( .A1(n173), .A2(n868), .B1(n862), .B2(n896), .ZN(n850) );
  INV_X1 U875 ( .A(N71), .ZN(n896) );
  OAI22_X1 U876 ( .A1(n165), .A2(n867), .B1(n861), .B2(n888), .ZN(n834) );
  INV_X1 U877 ( .A(N79), .ZN(n888) );
  OAI22_X1 U878 ( .A1(n162), .A2(n868), .B1(n861), .B2(n885), .ZN(n837) );
  INV_X1 U879 ( .A(N82), .ZN(n885) );
  XNOR2_X1 U880 ( .A(swp[4]), .B(swp[3]), .ZN(n802) );
  INV_X1 U881 ( .A(count_wait), .ZN(n874) );
  OAI21_X1 U882 ( .B1(n878), .B2(n802), .A(n387), .ZN(n204) );
  OAI21_X1 U883 ( .B1(swp[3]), .B2(n878), .A(n387), .ZN(n397) );
  OAI21_X1 U884 ( .B1(n193), .B2(n878), .A(n387), .ZN(n396) );
  OAI21_X1 U885 ( .B1(n192), .B2(n878), .A(n387), .ZN(n395) );
  OAI21_X1 U886 ( .B1(n191), .B2(n878), .A(n387), .ZN(n431) );
  NAND2_X1 U887 ( .A1(n803), .A2(n290), .ZN(n202) );
  NAND2_X1 U888 ( .A1(n803), .A2(N351), .ZN(n206) );
  NOR2_X1 U889 ( .A1(swp[3]), .A2(n879), .ZN(n210) );
  NOR2_X1 U890 ( .A1(n191), .A2(n879), .ZN(n283) );
  NOR2_X1 U891 ( .A1(n193), .A2(n879), .ZN(n208) );
  NOR2_X1 U892 ( .A1(n192), .A2(n879), .ZN(n209) );
  NAND2_X1 U893 ( .A1(N353), .A2(n803), .ZN(n198) );
  NAND2_X1 U894 ( .A1(N352), .A2(n803), .ZN(n200) );
  INV_X1 U895 ( .A(n858), .ZN(n860) );
  INV_X1 U896 ( .A(n725), .ZN(n871) );
  INV_X1 U897 ( .A(\U3/U1/Z_0 ), .ZN(n872) );
endmodule

