
module register_file_NBIT64_NREG32 ( CLK, RESET, ENABLE, RD1, RD2, WR, ADD_WR, 
        ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [63:0] DATAIN;
  output [63:0] OUT1;
  output [63:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n17148, n17149, n17156,
         n17157, n17161, n17163, n17169, n17170, n17177, n17178, n17182,
         n17184, n17190, n17191, n17198, n17199, n17203, n17205, n17211,
         n17212, n17219, n17220, n17224, n17226, n17232, n17233, n17240,
         n17241, n17245, n17247, n17253, n17254, n17261, n17262, n17266,
         n17268, n17274, n17275, n17282, n17283, n17287, n17289, n17295,
         n17296, n17303, n17304, n17308, n17310, n17316, n17317, n17324,
         n17325, n17329, n17331, n17337, n17338, n17345, n17346, n17350,
         n17352, n17358, n17359, n17366, n17367, n17371, n17373, n17379,
         n17380, n17387, n17388, n17392, n17394, n17400, n17401, n17408,
         n17409, n17413, n17415, n17421, n17422, n17429, n17430, n17434,
         n17436, n17442, n17443, n17450, n17451, n17455, n17457, n17463,
         n17464, n17471, n17472, n17476, n17478, n17484, n17485, n17492,
         n17493, n17497, n17499, n17505, n17506, n17513, n17514, n17518,
         n17520, n17526, n17527, n17534, n17535, n17539, n17541, n17547,
         n17548, n17555, n17556, n17560, n17562, n17568, n17569, n17576,
         n17577, n17581, n17583, n17589, n17590, n17597, n17598, n17602,
         n17604, n17610, n17611, n17618, n17619, n17623, n17625, n17631,
         n17632, n17639, n17640, n17644, n17646, n17652, n17653, n17660,
         n17661, n17665, n17667, n17673, n17674, n17681, n17682, n17686,
         n17688, n17694, n17695, n17702, n17703, n17707, n17709, n17715,
         n17716, n17723, n17724, n17728, n17730, n17736, n17737, n17744,
         n17745, n17749, n17751, n17757, n17758, n17765, n17766, n17770,
         n17772, n17778, n17779, n17786, n17787, n17791, n17793, n17799,
         n17800, n17807, n17808, n17812, n17814, n17820, n17821, n17828,
         n17829, n17833, n17835, n17841, n17842, n17849, n17850, n17854,
         n17856, n17862, n17863, n17870, n17871, n17875, n17877, n17883,
         n17884, n17891, n17892, n17896, n17898, n17904, n17905, n17912,
         n17913, n17917, n17919, n17925, n17926, n17933, n17934, n17938,
         n17940, n17946, n17947, n17954, n17955, n17959, n17961, n17967,
         n17968, n17975, n17976, n17980, n17982, n17988, n17989, n17996,
         n17997, n18001, n18003, n18009, n18010, n18017, n18018, n18022,
         n18024, n18030, n18031, n18038, n18039, n18043, n18045, n18051,
         n18052, n18059, n18060, n18064, n18066, n18072, n18073, n18080,
         n18081, n18085, n18087, n18093, n18094, n18101, n18102, n18106,
         n18108, n18114, n18115, n18122, n18123, n18127, n18129, n18135,
         n18136, n18143, n18144, n18148, n18150, n18156, n18157, n18164,
         n18165, n18169, n18171, n18177, n18178, n18185, n18186, n18190,
         n18192, n18198, n18199, n18206, n18207, n18211, n18213, n18219,
         n18220, n18227, n18228, n18232, n18234, n18240, n18241, n18248,
         n18249, n18253, n18255, n18261, n18262, n18269, n18270, n18274,
         n18276, n18282, n18283, n18290, n18291, n18295, n18297, n18303,
         n18304, n18311, n18312, n18316, n18318, n18324, n18325, n18332,
         n18333, n18337, n18339, n18345, n18346, n18353, n18354, n18358,
         n18360, n18366, n18367, n18374, n18375, n18379, n18381, n18387,
         n18388, n18395, n18396, n18400, n18402, n18408, n18409, n18416,
         n18417, n18421, n18423, n18429, n18430, n18437, n18438, n18442,
         n18444, n18450, n18451, n18458, n18459, n18463, n18465, n18471,
         n18472, n18479, n18480, n18484, n18486, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,
         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,
         n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
         n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
         n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168,
         n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176,
         n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
         n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192,
         n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200,
         n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
         n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216,
         n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224,
         n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232,
         n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240,
         n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
         n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256,
         n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264,
         n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
         n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
         n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288,
         n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296,
         n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304,
         n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
         n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,
         n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
         n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336,
         n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,
         n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
         n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360,
         n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368,
         n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
         n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
         n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,
         n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,
         n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408,
         n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,
         n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
         n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432,
         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,
         n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480,
         n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,
         n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
         n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504,
         n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512,
         n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520,
         n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528,
         n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536,
         n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544,
         n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552,
         n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560,
         n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
         n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576,
         n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584,
         n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592,
         n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600,
         n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608,
         n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616,
         n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624,
         n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
         n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
         n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648,
         n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656,
         n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664,
         n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672,
         n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680,
         n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688,
         n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696,
         n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,
         n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,
         n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720,
         n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728,
         n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736,
         n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744,
         n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752,
         n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,
         n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768,
         n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,
         n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
         n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792,
         n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800,
         n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808,
         n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,
         n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,
         n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
         n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840,
         n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,
         n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
         n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864,
         n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872,
         n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,
         n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888,
         n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,
         n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904,
         n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912,
         n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920,
         n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,
         n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936,
         n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944,
         n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
         n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960,
         n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,
         n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976,
         n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984,
         n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992,
         n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,
         n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008,
         n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016,
         n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
         n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032,
         n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040,
         n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048,
         n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056,
         n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,
         n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,
         n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080,
         n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088,
         n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
         n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104,
         n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,
         n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120,
         n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128,
         n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,
         n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
         n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152,
         n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160,
         n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
         n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176,
         n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184,
         n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192,
         n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200,
         n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208,
         n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
         n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224,
         n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232,
         n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
         n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248,
         n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256,
         n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,
         n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,
         n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280,
         n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
         n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296,
         n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304,
         n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
         n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320,
         n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
         n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,
         n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
         n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,
         n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
         n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368,
         n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
         n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,
         n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392,
         n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,
         n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,
         n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,
         n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424,
         n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432,
         n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440,
         n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448,
         n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456,
         n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464,
         n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472,
         n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480,
         n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488,
         n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496,
         n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504,
         n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512,
         n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520,
         n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528,
         n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536,
         n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544,
         n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552,
         n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560,
         n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568,
         n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576,
         n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584,
         n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592,
         n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600,
         n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608,
         n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616,
         n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624,
         n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632,
         n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640,
         n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648,
         n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656,
         n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664,
         n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672,
         n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680,
         n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688,
         n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696,
         n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704,
         n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712,
         n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,
         n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728,
         n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,
         n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744,
         n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752,
         n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760,
         n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768,
         n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776,
         n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784,
         n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792,
         n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800,
         n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808,
         n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816,
         n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824,
         n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832,
         n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840,
         n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848,
         n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856,
         n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864,
         n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872,
         n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880,
         n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888,
         n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896,
         n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904,
         n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912,
         n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920,
         n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928,
         n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936,
         n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944,
         n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952,
         n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960,
         n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968,
         n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976,
         n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984,
         n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992,
         n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000,
         n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008,
         n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016,
         n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024,
         n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032,
         n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040,
         n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048,
         n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056,
         n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064,
         n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072,
         n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,
         n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088,
         n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096,
         n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104,
         n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112,
         n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120,
         n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128,
         n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136,
         n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144,
         n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152,
         n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160,
         n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168,
         n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176,
         n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184,
         n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192,
         n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200,
         n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208,
         n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216,
         n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224,
         n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232,
         n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240,
         n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248,
         n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256,
         n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264,
         n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272,
         n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280,
         n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288,
         n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296,
         n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304,
         n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312,
         n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320,
         n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328,
         n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336,
         n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344,
         n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352,
         n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360,
         n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368,
         n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376,
         n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384,
         n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392,
         n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400,
         n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408,
         n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416,
         n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424,
         n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432,
         n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440,
         n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448,
         n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456,
         n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464,
         n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472,
         n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480,
         n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488,
         n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496,
         n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504,
         n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512,
         n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520,
         n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528,
         n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536,
         n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544,
         n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552,
         n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560,
         n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568,
         n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576,
         n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584,
         n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592,
         n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600,
         n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608,
         n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616,
         n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624,
         n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632,
         n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640,
         n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648,
         n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656,
         n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664,
         n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672,
         n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680,
         n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688,
         n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696,
         n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704,
         n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712,
         n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720,
         n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728,
         n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736,
         n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744,
         n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752,
         n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760,
         n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768,
         n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776,
         n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784,
         n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792,
         n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800,
         n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808,
         n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816,
         n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824,
         n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832,
         n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840,
         n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848,
         n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856,
         n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864,
         n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872,
         n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880,
         n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888,
         n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896,
         n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904,
         n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912,
         n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920,
         n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928,
         n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936,
         n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944,
         n23945, n23946, n23947, n23948, n23949, n23954, n23955, n23956,
         n23957, n24018, n24019, n24020, n24021, n24022, n24023, n24024,
         n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032,
         n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040,
         n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048,
         n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056,
         n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064,
         n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072,
         n24073, n24074, n24075, n24076, n24077, n24079, n24081, n24083,
         n24085, n24087, n24089, n24091, n24093, n24095, n24097, n24099,
         n24101, n24103, n24105, n24107, n24109, n24111, n24113, n24115,
         n24117, n24119, n24121, n24123, n24125, n24127, n24129, n24131,
         n24133, n24135, n24137, n24139, n24141, n24143, n24145, n24147,
         n24149, n24151, n24153, n24155, n24157, n24159, n24161, n24163,
         n24165, n24167, n24169, n24171, n24173, n24175, n24177, n24179,
         n24181, n24183, n24185, n24187, n24189, n24191, n24193, n24195,
         n24197, n24199, n24201, n24203, n24205, n24206, n24208, n24210,
         n24212, n24214, n24216, n24218, n24220, n24222, n24224, n24226,
         n24228, n24230, n24232, n24234, n24236, n24238, n24240, n24242,
         n24244, n24246, n24248, n24250, n24252, n24254, n24256, n24258,
         n24260, n24262, n24264, n24266, n24268, n24270, n24272, n24274,
         n24276, n24278, n24280, n24282, n24284, n24286, n24288, n24290,
         n24292, n24294, n24296, n24298, n24300, n24302, n24305, n24308,
         n24311, n24314, n24316, n24318, n24320, n24322, n24324, n24326,
         n24328, n24330, n24332, n24334, n24336, n24339, n24341, n24343,
         n24345, n24347, n24349, n24351, n24353, n24355, n24357, n24359,
         n24361, n24363, n24365, n24367, n24369, n24371, n24373, n24375,
         n24377, n24379, n24381, n24383, n24385, n24387, n24389, n24391,
         n24393, n24395, n24397, n24399, n24401, n24403, n24405, n24407,
         n24409, n24411, n24413, n24415, n24417, n24419, n24421, n24423,
         n24425, n24427, n24429, n24431, n24433, n24435, n24437, n24439,
         n24441, n24443, n24445, n24447, n24449, n24451, n24453, n24455,
         n24457, n24459, n24461, n24463, n24465, n24474, n24475, n24476,
         n24477, n24478, n24479, n24480, n24481, n24607, n24609, n24611,
         n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620,
         n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628,
         n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636,
         n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644,
         n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652,
         n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660,
         n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668,
         n24669, n24670, n24671, n24672, n24673, n24794, n24795, n24796,
         n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804,
         n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812,
         n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820,
         n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828,
         n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836,
         n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844,
         n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852,
         n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860,
         n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868,
         n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876,
         n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884,
         n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892,
         n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900,
         n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908,
         n24909, n24910, n24911, n24912, n24913, n24974, n24975, n24976,
         n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984,
         n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992,
         n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000,
         n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008,
         n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016,
         n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024,
         n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032,
         n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040,
         n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048,
         n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056,
         n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064,
         n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072,
         n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080,
         n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088,
         n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
         n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104,
         n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112,
         n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120,
         n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128,
         n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136,
         n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,
         n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152,
         n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160,
         n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,
         n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176,
         n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184,
         n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,
         n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200,
         n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208,
         n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216,
         n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224,
         n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232,
         n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240,
         n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248,
         n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256,
         n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264,
         n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272,
         n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280,
         n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288,
         n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296,
         n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304,
         n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312,
         n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320,
         n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328,
         n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336,
         n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344,
         n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352,
         n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360,
         n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368,
         n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376,
         n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,
         n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392,
         n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400,
         n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408,
         n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416,
         n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
         n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432,
         n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440,
         n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448,
         n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456,
         n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464,
         n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472,
         n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480,
         n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488,
         n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496,
         n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504,
         n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512,
         n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520,
         n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528,
         n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536,
         n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544,
         n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552,
         n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560,
         n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568,
         n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576,
         n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584,
         n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592,
         n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600,
         n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608,
         n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616,
         n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624,
         n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632,
         n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640,
         n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648,
         n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656,
         n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664,
         n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672,
         n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680,
         n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688,
         n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696,
         n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704,
         n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712,
         n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720,
         n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728,
         n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736,
         n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744,
         n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752,
         n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760,
         n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768,
         n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776,
         n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784,
         n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792,
         n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800,
         n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808,
         n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816,
         n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824,
         n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832,
         n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840,
         n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848,
         n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,
         n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864,
         n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872,
         n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880,
         n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888,
         n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896,
         n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904,
         n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912,
         n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920,
         n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928,
         n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936,
         n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944,
         n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952,
         n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960,
         n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968,
         n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976,
         n25977, n25978;

  DFF_X1 \OUT1_reg[63]  ( .D(n5438), .CK(CLK), .Q(OUT1[63]) );
  DFF_X1 \OUT1_reg[62]  ( .D(n5437), .CK(CLK), .Q(OUT1[62]) );
  DFF_X1 \OUT1_reg[61]  ( .D(n5436), .CK(CLK), .Q(OUT1[61]) );
  DFF_X1 \OUT1_reg[60]  ( .D(n5435), .CK(CLK), .Q(OUT1[60]) );
  DFF_X1 \OUT1_reg[59]  ( .D(n5434), .CK(CLK), .Q(OUT1[59]) );
  DFF_X1 \OUT1_reg[58]  ( .D(n5433), .CK(CLK), .Q(OUT1[58]) );
  DFF_X1 \OUT1_reg[57]  ( .D(n5432), .CK(CLK), .Q(OUT1[57]) );
  DFF_X1 \OUT1_reg[56]  ( .D(n5431), .CK(CLK), .Q(OUT1[56]) );
  DFF_X1 \OUT1_reg[55]  ( .D(n5430), .CK(CLK), .Q(OUT1[55]) );
  DFF_X1 \OUT1_reg[54]  ( .D(n5429), .CK(CLK), .Q(OUT1[54]) );
  DFF_X1 \OUT1_reg[53]  ( .D(n5428), .CK(CLK), .Q(OUT1[53]) );
  DFF_X1 \OUT1_reg[52]  ( .D(n5427), .CK(CLK), .Q(OUT1[52]) );
  DFF_X1 \OUT1_reg[51]  ( .D(n5426), .CK(CLK), .Q(OUT1[51]) );
  DFF_X1 \OUT1_reg[50]  ( .D(n5425), .CK(CLK), .Q(OUT1[50]) );
  DFF_X1 \OUT1_reg[49]  ( .D(n5424), .CK(CLK), .Q(OUT1[49]) );
  DFF_X1 \OUT1_reg[48]  ( .D(n5423), .CK(CLK), .Q(OUT1[48]) );
  DFF_X1 \OUT1_reg[47]  ( .D(n5422), .CK(CLK), .Q(OUT1[47]) );
  DFF_X1 \OUT1_reg[46]  ( .D(n5421), .CK(CLK), .Q(OUT1[46]) );
  DFF_X1 \OUT1_reg[45]  ( .D(n5420), .CK(CLK), .Q(OUT1[45]) );
  DFF_X1 \OUT1_reg[44]  ( .D(n5419), .CK(CLK), .Q(OUT1[44]) );
  DFF_X1 \OUT1_reg[43]  ( .D(n5418), .CK(CLK), .Q(OUT1[43]) );
  DFF_X1 \OUT1_reg[42]  ( .D(n5417), .CK(CLK), .Q(OUT1[42]) );
  DFF_X1 \OUT1_reg[41]  ( .D(n5416), .CK(CLK), .Q(OUT1[41]) );
  DFF_X1 \OUT1_reg[40]  ( .D(n5415), .CK(CLK), .Q(OUT1[40]) );
  DFF_X1 \OUT1_reg[39]  ( .D(n5414), .CK(CLK), .Q(OUT1[39]) );
  DFF_X1 \OUT1_reg[38]  ( .D(n5413), .CK(CLK), .Q(OUT1[38]) );
  DFF_X1 \OUT1_reg[37]  ( .D(n5412), .CK(CLK), .Q(OUT1[37]) );
  DFF_X1 \OUT1_reg[36]  ( .D(n5411), .CK(CLK), .Q(OUT1[36]) );
  DFF_X1 \OUT1_reg[35]  ( .D(n5410), .CK(CLK), .Q(OUT1[35]) );
  DFF_X1 \OUT1_reg[34]  ( .D(n5409), .CK(CLK), .Q(OUT1[34]) );
  DFF_X1 \OUT1_reg[33]  ( .D(n5408), .CK(CLK), .Q(OUT1[33]) );
  DFF_X1 \OUT1_reg[32]  ( .D(n5407), .CK(CLK), .Q(OUT1[32]) );
  DFF_X1 \OUT1_reg[31]  ( .D(n5406), .CK(CLK), .Q(OUT1[31]) );
  DFF_X1 \OUT1_reg[30]  ( .D(n5405), .CK(CLK), .Q(OUT1[30]) );
  DFF_X1 \OUT1_reg[29]  ( .D(n5404), .CK(CLK), .Q(OUT1[29]) );
  DFF_X1 \OUT1_reg[28]  ( .D(n5403), .CK(CLK), .Q(OUT1[28]) );
  DFF_X1 \OUT1_reg[27]  ( .D(n5402), .CK(CLK), .Q(OUT1[27]) );
  DFF_X1 \OUT1_reg[26]  ( .D(n5401), .CK(CLK), .Q(OUT1[26]) );
  DFF_X1 \OUT1_reg[25]  ( .D(n5400), .CK(CLK), .Q(OUT1[25]) );
  DFF_X1 \OUT1_reg[24]  ( .D(n5399), .CK(CLK), .Q(OUT1[24]) );
  DFF_X1 \OUT1_reg[23]  ( .D(n5398), .CK(CLK), .Q(OUT1[23]) );
  DFF_X1 \OUT1_reg[22]  ( .D(n5397), .CK(CLK), .Q(OUT1[22]) );
  DFF_X1 \OUT1_reg[21]  ( .D(n5396), .CK(CLK), .Q(OUT1[21]) );
  DFF_X1 \OUT1_reg[20]  ( .D(n5395), .CK(CLK), .Q(OUT1[20]) );
  DFF_X1 \OUT1_reg[19]  ( .D(n5394), .CK(CLK), .Q(OUT1[19]) );
  DFF_X1 \OUT1_reg[18]  ( .D(n5393), .CK(CLK), .Q(OUT1[18]) );
  DFF_X1 \OUT1_reg[17]  ( .D(n5392), .CK(CLK), .Q(OUT1[17]) );
  DFF_X1 \OUT1_reg[16]  ( .D(n5391), .CK(CLK), .Q(OUT1[16]) );
  DFF_X1 \OUT1_reg[15]  ( .D(n5390), .CK(CLK), .Q(OUT1[15]) );
  DFF_X1 \OUT1_reg[14]  ( .D(n5389), .CK(CLK), .Q(OUT1[14]) );
  DFF_X1 \OUT1_reg[13]  ( .D(n5388), .CK(CLK), .Q(OUT1[13]) );
  DFF_X1 \OUT1_reg[12]  ( .D(n5387), .CK(CLK), .Q(OUT1[12]) );
  DFF_X1 \OUT1_reg[11]  ( .D(n5386), .CK(CLK), .Q(OUT1[11]) );
  DFF_X1 \OUT1_reg[10]  ( .D(n5385), .CK(CLK), .Q(OUT1[10]) );
  DFF_X1 \OUT1_reg[9]  ( .D(n5384), .CK(CLK), .Q(OUT1[9]) );
  DFF_X1 \OUT1_reg[8]  ( .D(n5383), .CK(CLK), .Q(OUT1[8]) );
  DFF_X1 \OUT1_reg[7]  ( .D(n5382), .CK(CLK), .Q(OUT1[7]) );
  DFF_X1 \OUT1_reg[6]  ( .D(n5381), .CK(CLK), .Q(OUT1[6]) );
  DFF_X1 \OUT1_reg[5]  ( .D(n5380), .CK(CLK), .Q(OUT1[5]) );
  DFF_X1 \OUT1_reg[4]  ( .D(n5379), .CK(CLK), .Q(OUT1[4]) );
  DFF_X1 \OUT1_reg[3]  ( .D(n5378), .CK(CLK), .Q(OUT1[3]) );
  DFF_X1 \OUT1_reg[2]  ( .D(n5377), .CK(CLK), .Q(OUT1[2]) );
  DFF_X1 \OUT1_reg[1]  ( .D(n5376), .CK(CLK), .Q(OUT1[1]) );
  DFF_X1 \OUT1_reg[0]  ( .D(n5375), .CK(CLK), .Q(OUT1[0]) );
  DFF_X1 \OUT2_reg[62]  ( .D(n5373), .CK(CLK), .Q(OUT2[62]) );
  DFF_X1 \OUT2_reg[61]  ( .D(n5372), .CK(CLK), .Q(OUT2[61]) );
  DFF_X1 \OUT2_reg[60]  ( .D(n5371), .CK(CLK), .Q(OUT2[60]) );
  DFF_X1 \OUT2_reg[59]  ( .D(n5370), .CK(CLK), .Q(OUT2[59]) );
  DFF_X1 \OUT2_reg[58]  ( .D(n5369), .CK(CLK), .Q(OUT2[58]) );
  DFF_X1 \OUT2_reg[57]  ( .D(n5368), .CK(CLK), .Q(OUT2[57]) );
  DFF_X1 \OUT2_reg[56]  ( .D(n5367), .CK(CLK), .Q(OUT2[56]) );
  DFF_X1 \OUT2_reg[55]  ( .D(n5366), .CK(CLK), .Q(OUT2[55]) );
  DFF_X1 \OUT2_reg[54]  ( .D(n5365), .CK(CLK), .Q(OUT2[54]) );
  DFF_X1 \OUT2_reg[53]  ( .D(n5364), .CK(CLK), .Q(OUT2[53]) );
  DFF_X1 \OUT2_reg[52]  ( .D(n5363), .CK(CLK), .Q(OUT2[52]) );
  DFF_X1 \OUT2_reg[51]  ( .D(n5362), .CK(CLK), .Q(OUT2[51]) );
  DFF_X1 \OUT2_reg[50]  ( .D(n5361), .CK(CLK), .Q(OUT2[50]) );
  DFF_X1 \OUT2_reg[49]  ( .D(n5360), .CK(CLK), .Q(OUT2[49]) );
  DFF_X1 \OUT2_reg[48]  ( .D(n5359), .CK(CLK), .Q(OUT2[48]) );
  DFF_X1 \OUT2_reg[47]  ( .D(n5358), .CK(CLK), .Q(OUT2[47]) );
  DFF_X1 \OUT2_reg[46]  ( .D(n5357), .CK(CLK), .Q(OUT2[46]) );
  DFF_X1 \OUT2_reg[45]  ( .D(n5356), .CK(CLK), .Q(OUT2[45]) );
  DFF_X1 \OUT2_reg[44]  ( .D(n5355), .CK(CLK), .Q(OUT2[44]) );
  DFF_X1 \OUT2_reg[43]  ( .D(n5354), .CK(CLK), .Q(OUT2[43]) );
  DFF_X1 \OUT2_reg[42]  ( .D(n5353), .CK(CLK), .Q(OUT2[42]) );
  DFF_X1 \OUT2_reg[41]  ( .D(n5352), .CK(CLK), .Q(OUT2[41]) );
  DFF_X1 \OUT2_reg[40]  ( .D(n5351), .CK(CLK), .Q(OUT2[40]) );
  DFF_X1 \OUT2_reg[39]  ( .D(n5350), .CK(CLK), .Q(OUT2[39]) );
  DFF_X1 \OUT2_reg[38]  ( .D(n5349), .CK(CLK), .Q(OUT2[38]) );
  DFF_X1 \OUT2_reg[37]  ( .D(n5348), .CK(CLK), .Q(OUT2[37]) );
  DFF_X1 \OUT2_reg[36]  ( .D(n5347), .CK(CLK), .Q(OUT2[36]) );
  DFF_X1 \OUT2_reg[35]  ( .D(n5346), .CK(CLK), .Q(OUT2[35]) );
  DFF_X1 \OUT2_reg[34]  ( .D(n5345), .CK(CLK), .Q(OUT2[34]) );
  DFF_X1 \OUT2_reg[33]  ( .D(n5344), .CK(CLK), .Q(OUT2[33]) );
  DFF_X1 \OUT2_reg[32]  ( .D(n5343), .CK(CLK), .Q(OUT2[32]) );
  DFF_X1 \OUT2_reg[31]  ( .D(n5342), .CK(CLK), .Q(OUT2[31]) );
  DFF_X1 \OUT2_reg[30]  ( .D(n5341), .CK(CLK), .Q(OUT2[30]) );
  DFF_X1 \OUT2_reg[29]  ( .D(n5340), .CK(CLK), .Q(OUT2[29]) );
  DFF_X1 \OUT2_reg[28]  ( .D(n5339), .CK(CLK), .Q(OUT2[28]) );
  DFF_X1 \OUT2_reg[27]  ( .D(n5338), .CK(CLK), .Q(OUT2[27]) );
  DFF_X1 \OUT2_reg[26]  ( .D(n5337), .CK(CLK), .Q(OUT2[26]) );
  DFF_X1 \OUT2_reg[25]  ( .D(n5336), .CK(CLK), .Q(OUT2[25]) );
  DFF_X1 \OUT2_reg[24]  ( .D(n5335), .CK(CLK), .Q(OUT2[24]) );
  DFF_X1 \OUT2_reg[23]  ( .D(n5334), .CK(CLK), .Q(OUT2[23]) );
  DFF_X1 \OUT2_reg[22]  ( .D(n5333), .CK(CLK), .Q(OUT2[22]) );
  DFF_X1 \OUT2_reg[21]  ( .D(n5332), .CK(CLK), .Q(OUT2[21]) );
  DFF_X1 \OUT2_reg[20]  ( .D(n5331), .CK(CLK), .Q(OUT2[20]) );
  DFF_X1 \OUT2_reg[19]  ( .D(n5330), .CK(CLK), .Q(OUT2[19]) );
  DFF_X1 \OUT2_reg[18]  ( .D(n5329), .CK(CLK), .Q(OUT2[18]) );
  DFF_X1 \OUT2_reg[17]  ( .D(n5328), .CK(CLK), .Q(OUT2[17]) );
  DFF_X1 \OUT2_reg[16]  ( .D(n5327), .CK(CLK), .Q(OUT2[16]) );
  DFF_X1 \OUT2_reg[15]  ( .D(n5326), .CK(CLK), .Q(OUT2[15]) );
  DFF_X1 \OUT2_reg[14]  ( .D(n5325), .CK(CLK), .Q(OUT2[14]) );
  DFF_X1 \OUT2_reg[13]  ( .D(n5324), .CK(CLK), .Q(OUT2[13]) );
  DFF_X1 \OUT2_reg[12]  ( .D(n5323), .CK(CLK), .Q(OUT2[12]) );
  DFF_X1 \OUT2_reg[11]  ( .D(n5322), .CK(CLK), .Q(OUT2[11]) );
  DFF_X1 \OUT2_reg[10]  ( .D(n5321), .CK(CLK), .Q(OUT2[10]) );
  DFF_X1 \OUT2_reg[9]  ( .D(n5320), .CK(CLK), .Q(OUT2[9]) );
  DFF_X1 \OUT2_reg[8]  ( .D(n5319), .CK(CLK), .Q(OUT2[8]) );
  DFF_X1 \OUT2_reg[7]  ( .D(n5318), .CK(CLK), .Q(OUT2[7]) );
  DFF_X1 \OUT2_reg[6]  ( .D(n5317), .CK(CLK), .Q(OUT2[6]) );
  DFF_X1 \OUT2_reg[5]  ( .D(n5316), .CK(CLK), .Q(OUT2[5]) );
  DFF_X1 \OUT2_reg[4]  ( .D(n5315), .CK(CLK), .Q(OUT2[4]) );
  DFF_X1 \OUT2_reg[3]  ( .D(n5314), .CK(CLK), .Q(OUT2[3]) );
  DFF_X1 \OUT2_reg[2]  ( .D(n5313), .CK(CLK), .Q(OUT2[2]) );
  DFF_X1 \OUT2_reg[1]  ( .D(n5312), .CK(CLK), .Q(OUT2[1]) );
  DFF_X1 \OUT2_reg[0]  ( .D(n5311), .CK(CLK), .Q(OUT2[0]) );
  DFF_X1 \REGISTERS_reg[0][63]  ( .D(n7486), .CK(CLK), .QN(n9415) );
  DFF_X1 \REGISTERS_reg[0][62]  ( .D(n7485), .CK(CLK), .QN(n9416) );
  DFF_X1 \REGISTERS_reg[0][61]  ( .D(n7484), .CK(CLK), .QN(n9417) );
  DFF_X1 \REGISTERS_reg[0][60]  ( .D(n7483), .CK(CLK), .QN(n9418) );
  DFF_X1 \REGISTERS_reg[0][59]  ( .D(n7482), .CK(CLK), .QN(n9419) );
  DFF_X1 \REGISTERS_reg[0][58]  ( .D(n7481), .CK(CLK), .QN(n9420) );
  DFF_X1 \REGISTERS_reg[0][57]  ( .D(n7480), .CK(CLK), .QN(n9421) );
  DFF_X1 \REGISTERS_reg[0][56]  ( .D(n7479), .CK(CLK), .QN(n9422) );
  DFF_X1 \REGISTERS_reg[0][55]  ( .D(n7478), .CK(CLK), .QN(n9423) );
  DFF_X1 \REGISTERS_reg[0][54]  ( .D(n7477), .CK(CLK), .QN(n9424) );
  DFF_X1 \REGISTERS_reg[0][53]  ( .D(n7476), .CK(CLK), .QN(n9425) );
  DFF_X1 \REGISTERS_reg[0][52]  ( .D(n7475), .CK(CLK), .QN(n9426) );
  DFF_X1 \REGISTERS_reg[0][51]  ( .D(n7474), .CK(CLK), .QN(n9427) );
  DFF_X1 \REGISTERS_reg[0][50]  ( .D(n7473), .CK(CLK), .QN(n9428) );
  DFF_X1 \REGISTERS_reg[0][49]  ( .D(n7472), .CK(CLK), .QN(n9429) );
  DFF_X1 \REGISTERS_reg[0][48]  ( .D(n7471), .CK(CLK), .QN(n9430) );
  DFF_X1 \REGISTERS_reg[0][47]  ( .D(n7470), .CK(CLK), .QN(n9431) );
  DFF_X1 \REGISTERS_reg[0][46]  ( .D(n7469), .CK(CLK), .QN(n9432) );
  DFF_X1 \REGISTERS_reg[0][45]  ( .D(n7468), .CK(CLK), .QN(n9433) );
  DFF_X1 \REGISTERS_reg[0][44]  ( .D(n7467), .CK(CLK), .QN(n9434) );
  DFF_X1 \REGISTERS_reg[0][43]  ( .D(n7466), .CK(CLK), .QN(n9435) );
  DFF_X1 \REGISTERS_reg[0][42]  ( .D(n7465), .CK(CLK), .QN(n9436) );
  DFF_X1 \REGISTERS_reg[0][41]  ( .D(n7464), .CK(CLK), .QN(n9437) );
  DFF_X1 \REGISTERS_reg[0][40]  ( .D(n7463), .CK(CLK), .QN(n9438) );
  DFF_X1 \REGISTERS_reg[0][39]  ( .D(n7462), .CK(CLK), .QN(n9439) );
  DFF_X1 \REGISTERS_reg[0][38]  ( .D(n7461), .CK(CLK), .QN(n9440) );
  DFF_X1 \REGISTERS_reg[0][37]  ( .D(n7460), .CK(CLK), .QN(n9441) );
  DFF_X1 \REGISTERS_reg[0][36]  ( .D(n7459), .CK(CLK), .QN(n9442) );
  DFF_X1 \REGISTERS_reg[0][35]  ( .D(n7458), .CK(CLK), .QN(n9443) );
  DFF_X1 \REGISTERS_reg[0][34]  ( .D(n7457), .CK(CLK), .QN(n9444) );
  DFF_X1 \REGISTERS_reg[0][33]  ( .D(n7456), .CK(CLK), .QN(n9445) );
  DFF_X1 \REGISTERS_reg[0][32]  ( .D(n7455), .CK(CLK), .QN(n9446) );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n7454), .CK(CLK), .QN(n9447) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n7453), .CK(CLK), .QN(n9448) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n7452), .CK(CLK), .QN(n9449) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n7451), .CK(CLK), .QN(n9450) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n7450), .CK(CLK), .QN(n9451) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n7449), .CK(CLK), .QN(n9452) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n7448), .CK(CLK), .QN(n9453) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n7447), .CK(CLK), .QN(n9454) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n7446), .CK(CLK), .QN(n9455) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n7445), .CK(CLK), .QN(n9456) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n7444), .CK(CLK), .QN(n9457) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n7443), .CK(CLK), .QN(n9458) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n7442), .CK(CLK), .QN(n9459) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n7441), .CK(CLK), .QN(n9460) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n7440), .CK(CLK), .QN(n9461) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n7439), .CK(CLK), .QN(n9462) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n7438), .CK(CLK), .QN(n9463) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n7437), .CK(CLK), .QN(n9464) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n7436), .CK(CLK), .QN(n9465) );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n7435), .CK(CLK), .QN(n9466) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n7434), .CK(CLK), .QN(n9467) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n7433), .CK(CLK), .QN(n9468) );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n7432), .CK(CLK), .QN(n9469) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n7431), .CK(CLK), .QN(n9470) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n7430), .CK(CLK), .QN(n9471) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n7429), .CK(CLK), .QN(n9472) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n7428), .CK(CLK), .QN(n9473) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n7427), .CK(CLK), .QN(n9474) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n7426), .CK(CLK), .QN(n9475) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n7425), .CK(CLK), .QN(n9476) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n7424), .CK(CLK), .QN(n9477) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n7423), .CK(CLK), .QN(n9478) );
  DFF_X1 \REGISTERS_reg[21][62]  ( .D(n6141), .CK(CLK), .QN(n8968) );
  DFF_X1 \REGISTERS_reg[21][61]  ( .D(n6140), .CK(CLK), .QN(n8969) );
  DFF_X1 \REGISTERS_reg[21][60]  ( .D(n6139), .CK(CLK), .QN(n8970) );
  DFF_X1 \REGISTERS_reg[21][59]  ( .D(n6138), .CK(CLK), .QN(n8971) );
  DFF_X1 \REGISTERS_reg[21][58]  ( .D(n6137), .CK(CLK), .QN(n8972) );
  DFF_X1 \REGISTERS_reg[21][57]  ( .D(n6136), .CK(CLK), .QN(n8973) );
  DFF_X1 \REGISTERS_reg[21][56]  ( .D(n6135), .CK(CLK), .QN(n8974) );
  DFF_X1 \REGISTERS_reg[21][55]  ( .D(n6134), .CK(CLK), .QN(n8975) );
  DFF_X1 \REGISTERS_reg[21][54]  ( .D(n6133), .CK(CLK), .QN(n8976) );
  DFF_X1 \REGISTERS_reg[21][53]  ( .D(n6132), .CK(CLK), .QN(n8977) );
  DFF_X1 \REGISTERS_reg[21][52]  ( .D(n6131), .CK(CLK), .QN(n8978) );
  DFF_X1 \REGISTERS_reg[21][51]  ( .D(n6130), .CK(CLK), .QN(n8979) );
  DFF_X1 \REGISTERS_reg[21][50]  ( .D(n6129), .CK(CLK), .QN(n8980) );
  DFF_X1 \REGISTERS_reg[21][49]  ( .D(n6128), .CK(CLK), .QN(n8981) );
  DFF_X1 \REGISTERS_reg[21][48]  ( .D(n6127), .CK(CLK), .QN(n8982) );
  DFF_X1 \REGISTERS_reg[21][47]  ( .D(n6126), .CK(CLK), .QN(n8983) );
  DFF_X1 \REGISTERS_reg[21][46]  ( .D(n6125), .CK(CLK), .QN(n8984) );
  DFF_X1 \REGISTERS_reg[21][45]  ( .D(n6124), .CK(CLK), .QN(n8985) );
  DFF_X1 \REGISTERS_reg[21][44]  ( .D(n6123), .CK(CLK), .QN(n8986) );
  DFF_X1 \REGISTERS_reg[21][43]  ( .D(n6122), .CK(CLK), .QN(n8987) );
  DFF_X1 \REGISTERS_reg[21][42]  ( .D(n6121), .CK(CLK), .QN(n8988) );
  DFF_X1 \REGISTERS_reg[21][41]  ( .D(n6120), .CK(CLK), .QN(n8989) );
  DFF_X1 \REGISTERS_reg[21][40]  ( .D(n6119), .CK(CLK), .QN(n8990) );
  DFF_X1 \REGISTERS_reg[21][39]  ( .D(n6118), .CK(CLK), .QN(n8991) );
  DFF_X1 \REGISTERS_reg[21][38]  ( .D(n6117), .CK(CLK), .QN(n8992) );
  DFF_X1 \REGISTERS_reg[21][37]  ( .D(n6116), .CK(CLK), .QN(n8993) );
  DFF_X1 \REGISTERS_reg[21][36]  ( .D(n6115), .CK(CLK), .QN(n8994) );
  DFF_X1 \REGISTERS_reg[21][35]  ( .D(n6114), .CK(CLK), .QN(n8995) );
  DFF_X1 \REGISTERS_reg[21][34]  ( .D(n6113), .CK(CLK), .QN(n8996) );
  DFF_X1 \REGISTERS_reg[21][33]  ( .D(n6112), .CK(CLK), .QN(n8997) );
  DFF_X1 \REGISTERS_reg[21][32]  ( .D(n6111), .CK(CLK), .QN(n8998) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n6110), .CK(CLK), .QN(n8999) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n6109), .CK(CLK), .QN(n9000) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n6108), .CK(CLK), .QN(n9001) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n6107), .CK(CLK), .QN(n9002) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n6106), .CK(CLK), .QN(n9003) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n6105), .CK(CLK), .QN(n9004) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n6104), .CK(CLK), .QN(n9005) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n6103), .CK(CLK), .QN(n9006) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n6102), .CK(CLK), .QN(n9007) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n6101), .CK(CLK), .QN(n9008) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n6100), .CK(CLK), .QN(n9009) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n6099), .CK(CLK), .QN(n9010) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n6098), .CK(CLK), .QN(n9011) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n6097), .CK(CLK), .QN(n9012) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n6096), .CK(CLK), .QN(n9013) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n6095), .CK(CLK), .QN(n9014) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n6094), .CK(CLK), .QN(n9015) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n6093), .CK(CLK), .QN(n9016) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n6092), .CK(CLK), .QN(n9017) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n6091), .CK(CLK), .QN(n9018) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n6090), .CK(CLK), .QN(n9019) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n6089), .CK(CLK), .QN(n9020) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n6088), .CK(CLK), .QN(n9021) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n6087), .CK(CLK), .QN(n9022) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n6086), .CK(CLK), .QN(n9023) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n6085), .CK(CLK), .QN(n9024) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n6084), .CK(CLK), .QN(n9025) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n6083), .CK(CLK), .QN(n9026) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n6082), .CK(CLK), .QN(n9027) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n6081), .CK(CLK), .QN(n9028) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n6080), .CK(CLK), .QN(n9029) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n6079), .CK(CLK), .QN(n9030) );
  NOR3_X2 U15207 ( .A1(n25244), .A2(ADD_RD1[1]), .A3(n19486), .ZN(n22733) );
  NOR3_X2 U16467 ( .A1(n25046), .A2(ADD_RD2[1]), .A3(n19491), .ZN(n23930) );
  NAND3_X1 U18471 ( .A1(n19481), .A2(n19480), .A3(n21491), .ZN(n21480) );
  NAND3_X1 U18472 ( .A1(n21491), .A2(n19480), .A3(ADD_WR[2]), .ZN(n21494) );
  NAND3_X1 U18473 ( .A1(n21491), .A2(n19481), .A3(ADD_WR[3]), .ZN(n21503) );
  NAND3_X1 U18474 ( .A1(ADD_WR[2]), .A2(n21491), .A3(ADD_WR[3]), .ZN(n21512)
         );
  NAND3_X1 U18475 ( .A1(n19481), .A2(n19480), .A3(n21528), .ZN(n21521) );
  NAND3_X1 U18476 ( .A1(ADD_WR[2]), .A2(n19480), .A3(n21528), .ZN(n21531) );
  NAND3_X1 U18477 ( .A1(ADD_WR[3]), .A2(n19481), .A3(n21528), .ZN(n21540) );
  NAND3_X1 U18478 ( .A1(ADD_WR[3]), .A2(ADD_WR[2]), .A3(n21528), .ZN(n21549)
         );
  NAND3_X1 U18479 ( .A1(ENABLE), .A2(n25978), .A3(RD1), .ZN(n21591) );
  NAND3_X1 U18480 ( .A1(ENABLE), .A2(n25978), .A3(RD2), .ZN(n22788) );
  DFF_X1 \REGISTERS_reg[7][63]  ( .D(n7038), .CK(CLK), .Q(n19941), .QN(n9287)
         );
  DFF_X1 \REGISTERS_reg[7][62]  ( .D(n7037), .CK(CLK), .Q(n19942), .QN(n9288)
         );
  DFF_X1 \REGISTERS_reg[7][61]  ( .D(n7036), .CK(CLK), .Q(n19943), .QN(n9289)
         );
  DFF_X1 \REGISTERS_reg[7][60]  ( .D(n7035), .CK(CLK), .Q(n19944), .QN(n9290)
         );
  DFF_X1 \REGISTERS_reg[7][59]  ( .D(n7034), .CK(CLK), .Q(n19945), .QN(n9291)
         );
  DFF_X1 \REGISTERS_reg[7][58]  ( .D(n7033), .CK(CLK), .Q(n19946), .QN(n9292)
         );
  DFF_X1 \REGISTERS_reg[7][57]  ( .D(n7032), .CK(CLK), .Q(n19947), .QN(n9293)
         );
  DFF_X1 \REGISTERS_reg[7][56]  ( .D(n7031), .CK(CLK), .Q(n19948), .QN(n9294)
         );
  DFF_X1 \REGISTERS_reg[7][55]  ( .D(n7030), .CK(CLK), .Q(n19949), .QN(n9295)
         );
  DFF_X1 \REGISTERS_reg[7][54]  ( .D(n7029), .CK(CLK), .Q(n19950), .QN(n9296)
         );
  DFF_X1 \REGISTERS_reg[7][53]  ( .D(n7028), .CK(CLK), .Q(n19951), .QN(n9297)
         );
  DFF_X1 \REGISTERS_reg[7][52]  ( .D(n7027), .CK(CLK), .Q(n19952), .QN(n9298)
         );
  DFF_X1 \REGISTERS_reg[7][51]  ( .D(n7026), .CK(CLK), .Q(n19953), .QN(n9299)
         );
  DFF_X1 \REGISTERS_reg[7][50]  ( .D(n7025), .CK(CLK), .Q(n19954), .QN(n9300)
         );
  DFF_X1 \REGISTERS_reg[7][49]  ( .D(n7024), .CK(CLK), .Q(n19955), .QN(n9301)
         );
  DFF_X1 \REGISTERS_reg[7][48]  ( .D(n7023), .CK(CLK), .Q(n19956), .QN(n9302)
         );
  DFF_X1 \REGISTERS_reg[7][47]  ( .D(n7022), .CK(CLK), .Q(n19957), .QN(n9303)
         );
  DFF_X1 \REGISTERS_reg[7][46]  ( .D(n7021), .CK(CLK), .Q(n19958), .QN(n9304)
         );
  DFF_X1 \REGISTERS_reg[7][45]  ( .D(n7020), .CK(CLK), .Q(n19959), .QN(n9305)
         );
  DFF_X1 \REGISTERS_reg[7][44]  ( .D(n7019), .CK(CLK), .Q(n19960), .QN(n9306)
         );
  DFF_X1 \REGISTERS_reg[7][43]  ( .D(n7018), .CK(CLK), .Q(n19961), .QN(n9307)
         );
  DFF_X1 \REGISTERS_reg[7][42]  ( .D(n7017), .CK(CLK), .Q(n19962), .QN(n9308)
         );
  DFF_X1 \REGISTERS_reg[7][41]  ( .D(n7016), .CK(CLK), .Q(n19963), .QN(n9309)
         );
  DFF_X1 \REGISTERS_reg[7][40]  ( .D(n7015), .CK(CLK), .Q(n19964), .QN(n9310)
         );
  DFF_X1 \REGISTERS_reg[7][39]  ( .D(n7014), .CK(CLK), .Q(n19965), .QN(n9311)
         );
  DFF_X1 \REGISTERS_reg[7][38]  ( .D(n7013), .CK(CLK), .Q(n19966), .QN(n9312)
         );
  DFF_X1 \REGISTERS_reg[7][37]  ( .D(n7012), .CK(CLK), .Q(n19967), .QN(n9313)
         );
  DFF_X1 \REGISTERS_reg[7][36]  ( .D(n7011), .CK(CLK), .Q(n19968), .QN(n9314)
         );
  DFF_X1 \REGISTERS_reg[7][35]  ( .D(n7010), .CK(CLK), .Q(n19969), .QN(n9315)
         );
  DFF_X1 \REGISTERS_reg[7][34]  ( .D(n7009), .CK(CLK), .Q(n19970), .QN(n9316)
         );
  DFF_X1 \REGISTERS_reg[7][33]  ( .D(n7008), .CK(CLK), .Q(n19971), .QN(n9317)
         );
  DFF_X1 \REGISTERS_reg[7][32]  ( .D(n7007), .CK(CLK), .Q(n19972), .QN(n9318)
         );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n7006), .CK(CLK), .Q(n19973), .QN(n9319)
         );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n7005), .CK(CLK), .Q(n19974), .QN(n9320)
         );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n7004), .CK(CLK), .Q(n19975), .QN(n9321)
         );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n7003), .CK(CLK), .Q(n19976), .QN(n9322)
         );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n7002), .CK(CLK), .Q(n19977), .QN(n9323)
         );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n7001), .CK(CLK), .Q(n19978), .QN(n9324)
         );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n7000), .CK(CLK), .Q(n19979), .QN(n9325)
         );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n6999), .CK(CLK), .Q(n19980), .QN(n9326)
         );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n6998), .CK(CLK), .Q(n19981), .QN(n9327)
         );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n6997), .CK(CLK), .Q(n19982), .QN(n9328)
         );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n6996), .CK(CLK), .Q(n19983), .QN(n9329)
         );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n6995), .CK(CLK), .Q(n19984), .QN(n9330)
         );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n6994), .CK(CLK), .Q(n19985), .QN(n9331)
         );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n6993), .CK(CLK), .Q(n19986), .QN(n9332)
         );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n6992), .CK(CLK), .Q(n19987), .QN(n9333)
         );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n6991), .CK(CLK), .Q(n19988), .QN(n9334)
         );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n6990), .CK(CLK), .Q(n19989), .QN(n9335)
         );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n6989), .CK(CLK), .Q(n19990), .QN(n9336)
         );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n6988), .CK(CLK), .Q(n19991), .QN(n9337)
         );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n6987), .CK(CLK), .Q(n19992), .QN(n9338)
         );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n6986), .CK(CLK), .Q(n19993), .QN(n9339)
         );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n6985), .CK(CLK), .Q(n19994), .QN(n9340)
         );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n6984), .CK(CLK), .Q(n19995), .QN(n9341)
         );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n6983), .CK(CLK), .Q(n19996), .QN(n9342)
         );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n6982), .CK(CLK), .Q(n19997), .QN(n9343)
         );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n6981), .CK(CLK), .Q(n19998), .QN(n9344)
         );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n6980), .CK(CLK), .Q(n19999), .QN(n9345)
         );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n6979), .CK(CLK), .Q(n20000), .QN(n9346)
         );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n6978), .CK(CLK), .Q(n20001), .QN(n9347)
         );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n6977), .CK(CLK), .Q(n20002), .QN(n9348)
         );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n6976), .CK(CLK), .Q(n20003), .QN(n9349)
         );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n6975), .CK(CLK), .Q(n20004), .QN(n9350)
         );
  DFF_X1 \REGISTERS_reg[2][63]  ( .D(n7358), .CK(CLK), .Q(n20005), .QN(n9031)
         );
  DFF_X1 \REGISTERS_reg[2][62]  ( .D(n7357), .CK(CLK), .Q(n20006), .QN(n9032)
         );
  DFF_X1 \REGISTERS_reg[2][61]  ( .D(n7356), .CK(CLK), .Q(n20007), .QN(n9033)
         );
  DFF_X1 \REGISTERS_reg[2][60]  ( .D(n7355), .CK(CLK), .Q(n20008), .QN(n9034)
         );
  DFF_X1 \REGISTERS_reg[2][59]  ( .D(n7354), .CK(CLK), .Q(n20009), .QN(n9035)
         );
  DFF_X1 \REGISTERS_reg[2][58]  ( .D(n7353), .CK(CLK), .Q(n20010), .QN(n9036)
         );
  DFF_X1 \REGISTERS_reg[2][57]  ( .D(n7352), .CK(CLK), .Q(n20011), .QN(n9037)
         );
  DFF_X1 \REGISTERS_reg[2][56]  ( .D(n7351), .CK(CLK), .Q(n20012), .QN(n9038)
         );
  DFF_X1 \REGISTERS_reg[2][55]  ( .D(n7350), .CK(CLK), .Q(n20013), .QN(n9039)
         );
  DFF_X1 \REGISTERS_reg[2][54]  ( .D(n7349), .CK(CLK), .Q(n20014), .QN(n9040)
         );
  DFF_X1 \REGISTERS_reg[2][53]  ( .D(n7348), .CK(CLK), .Q(n20015), .QN(n9041)
         );
  DFF_X1 \REGISTERS_reg[2][52]  ( .D(n7347), .CK(CLK), .Q(n20016), .QN(n9042)
         );
  DFF_X1 \REGISTERS_reg[2][51]  ( .D(n7346), .CK(CLK), .Q(n20017), .QN(n9043)
         );
  DFF_X1 \REGISTERS_reg[2][50]  ( .D(n7345), .CK(CLK), .Q(n20018), .QN(n9044)
         );
  DFF_X1 \REGISTERS_reg[2][49]  ( .D(n7344), .CK(CLK), .Q(n20019), .QN(n9045)
         );
  DFF_X1 \REGISTERS_reg[2][48]  ( .D(n7343), .CK(CLK), .Q(n20020), .QN(n9046)
         );
  DFF_X1 \REGISTERS_reg[2][47]  ( .D(n7342), .CK(CLK), .Q(n20021), .QN(n9047)
         );
  DFF_X1 \REGISTERS_reg[2][46]  ( .D(n7341), .CK(CLK), .Q(n20022), .QN(n9048)
         );
  DFF_X1 \REGISTERS_reg[2][45]  ( .D(n7340), .CK(CLK), .Q(n20023), .QN(n9049)
         );
  DFF_X1 \REGISTERS_reg[2][44]  ( .D(n7339), .CK(CLK), .Q(n20024), .QN(n9050)
         );
  DFF_X1 \REGISTERS_reg[2][43]  ( .D(n7338), .CK(CLK), .Q(n20025), .QN(n9051)
         );
  DFF_X1 \REGISTERS_reg[2][42]  ( .D(n7337), .CK(CLK), .Q(n20026), .QN(n9052)
         );
  DFF_X1 \REGISTERS_reg[2][41]  ( .D(n7336), .CK(CLK), .Q(n20027), .QN(n9053)
         );
  DFF_X1 \REGISTERS_reg[2][40]  ( .D(n7335), .CK(CLK), .Q(n20028), .QN(n9054)
         );
  DFF_X1 \REGISTERS_reg[2][39]  ( .D(n7334), .CK(CLK), .Q(n20029), .QN(n9055)
         );
  DFF_X1 \REGISTERS_reg[2][38]  ( .D(n7333), .CK(CLK), .Q(n20030), .QN(n9056)
         );
  DFF_X1 \REGISTERS_reg[2][37]  ( .D(n7332), .CK(CLK), .Q(n20031), .QN(n9057)
         );
  DFF_X1 \REGISTERS_reg[2][36]  ( .D(n7331), .CK(CLK), .Q(n20032), .QN(n9058)
         );
  DFF_X1 \REGISTERS_reg[2][35]  ( .D(n7330), .CK(CLK), .Q(n20033), .QN(n9059)
         );
  DFF_X1 \REGISTERS_reg[2][34]  ( .D(n7329), .CK(CLK), .Q(n20034), .QN(n9060)
         );
  DFF_X1 \REGISTERS_reg[2][33]  ( .D(n7328), .CK(CLK), .Q(n20035), .QN(n9061)
         );
  DFF_X1 \REGISTERS_reg[2][32]  ( .D(n7327), .CK(CLK), .Q(n20036), .QN(n9062)
         );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n7326), .CK(CLK), .Q(n20037), .QN(n9063)
         );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n7325), .CK(CLK), .Q(n20038), .QN(n9064)
         );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n7324), .CK(CLK), .Q(n20039), .QN(n9065)
         );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n7323), .CK(CLK), .Q(n20040), .QN(n9066)
         );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n7322), .CK(CLK), .Q(n20041), .QN(n9067)
         );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n7321), .CK(CLK), .Q(n20042), .QN(n9068)
         );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n7320), .CK(CLK), .Q(n20043), .QN(n9069)
         );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n7319), .CK(CLK), .Q(n20044), .QN(n9070)
         );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n7318), .CK(CLK), .Q(n20045), .QN(n9071)
         );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n7317), .CK(CLK), .Q(n20046), .QN(n9072)
         );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n7316), .CK(CLK), .Q(n20047), .QN(n9073)
         );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n7315), .CK(CLK), .Q(n20048), .QN(n9074)
         );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n7314), .CK(CLK), .Q(n20049), .QN(n9075)
         );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n7313), .CK(CLK), .Q(n20050), .QN(n9076)
         );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n7312), .CK(CLK), .Q(n20051), .QN(n9077)
         );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n7311), .CK(CLK), .Q(n20052), .QN(n9078)
         );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n7310), .CK(CLK), .Q(n20053), .QN(n9079)
         );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n7309), .CK(CLK), .Q(n20054), .QN(n9080)
         );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n7308), .CK(CLK), .Q(n20055), .QN(n9081)
         );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n7307), .CK(CLK), .Q(n20056), .QN(n9082)
         );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n7306), .CK(CLK), .Q(n20057), .QN(n9083)
         );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n7305), .CK(CLK), .Q(n20058), .QN(n9084)
         );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n7304), .CK(CLK), .Q(n20059), .QN(n9085)
         );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n7303), .CK(CLK), .Q(n20060), .QN(n9086)
         );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n7302), .CK(CLK), .Q(n20061), .QN(n9087)
         );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n7301), .CK(CLK), .Q(n20062), .QN(n9088)
         );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n7300), .CK(CLK), .Q(n20063), .QN(n9089)
         );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n7299), .CK(CLK), .Q(n20064), .QN(n9090)
         );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n7298), .CK(CLK), .Q(n20065), .QN(n9091)
         );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n7297), .CK(CLK), .Q(n20066), .QN(n9092)
         );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n7296), .CK(CLK), .Q(n20067), .QN(n9093)
         );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n7295), .CK(CLK), .Q(n20068), .QN(n9094)
         );
  DFF_X1 \REGISTERS_reg[15][63]  ( .D(n6526), .CK(CLK), .Q(n20069), .QN(n9223)
         );
  DFF_X1 \REGISTERS_reg[15][62]  ( .D(n6525), .CK(CLK), .Q(n20070), .QN(n9224)
         );
  DFF_X1 \REGISTERS_reg[15][61]  ( .D(n6524), .CK(CLK), .Q(n20071), .QN(n9225)
         );
  DFF_X1 \REGISTERS_reg[15][60]  ( .D(n6523), .CK(CLK), .Q(n20072), .QN(n9226)
         );
  DFF_X1 \REGISTERS_reg[15][59]  ( .D(n6522), .CK(CLK), .Q(n20073), .QN(n9227)
         );
  DFF_X1 \REGISTERS_reg[15][58]  ( .D(n6521), .CK(CLK), .Q(n20074), .QN(n9228)
         );
  DFF_X1 \REGISTERS_reg[15][57]  ( .D(n6520), .CK(CLK), .Q(n20075), .QN(n9229)
         );
  DFF_X1 \REGISTERS_reg[15][56]  ( .D(n6519), .CK(CLK), .Q(n20076), .QN(n9230)
         );
  DFF_X1 \REGISTERS_reg[15][55]  ( .D(n6518), .CK(CLK), .Q(n20077), .QN(n9231)
         );
  DFF_X1 \REGISTERS_reg[15][54]  ( .D(n6517), .CK(CLK), .Q(n20078), .QN(n9232)
         );
  DFF_X1 \REGISTERS_reg[15][53]  ( .D(n6516), .CK(CLK), .Q(n20079), .QN(n9233)
         );
  DFF_X1 \REGISTERS_reg[15][52]  ( .D(n6515), .CK(CLK), .Q(n20080), .QN(n9234)
         );
  DFF_X1 \REGISTERS_reg[15][51]  ( .D(n6514), .CK(CLK), .Q(n20081), .QN(n9235)
         );
  DFF_X1 \REGISTERS_reg[15][50]  ( .D(n6513), .CK(CLK), .Q(n20082), .QN(n9236)
         );
  DFF_X1 \REGISTERS_reg[15][49]  ( .D(n6512), .CK(CLK), .Q(n20083), .QN(n9237)
         );
  DFF_X1 \REGISTERS_reg[15][48]  ( .D(n6511), .CK(CLK), .Q(n20084), .QN(n9238)
         );
  DFF_X1 \REGISTERS_reg[15][47]  ( .D(n6510), .CK(CLK), .Q(n20085), .QN(n9239)
         );
  DFF_X1 \REGISTERS_reg[15][46]  ( .D(n6509), .CK(CLK), .Q(n20086), .QN(n9240)
         );
  DFF_X1 \REGISTERS_reg[15][45]  ( .D(n6508), .CK(CLK), .Q(n20087), .QN(n9241)
         );
  DFF_X1 \REGISTERS_reg[15][44]  ( .D(n6507), .CK(CLK), .Q(n20088), .QN(n9242)
         );
  DFF_X1 \REGISTERS_reg[15][43]  ( .D(n6506), .CK(CLK), .Q(n20089), .QN(n9243)
         );
  DFF_X1 \REGISTERS_reg[15][42]  ( .D(n6505), .CK(CLK), .Q(n20090), .QN(n9244)
         );
  DFF_X1 \REGISTERS_reg[15][41]  ( .D(n6504), .CK(CLK), .Q(n20091), .QN(n9245)
         );
  DFF_X1 \REGISTERS_reg[15][40]  ( .D(n6503), .CK(CLK), .Q(n20092), .QN(n9246)
         );
  DFF_X1 \REGISTERS_reg[15][39]  ( .D(n6502), .CK(CLK), .Q(n20093), .QN(n9247)
         );
  DFF_X1 \REGISTERS_reg[15][38]  ( .D(n6501), .CK(CLK), .Q(n20094), .QN(n9248)
         );
  DFF_X1 \REGISTERS_reg[15][37]  ( .D(n6500), .CK(CLK), .Q(n20095), .QN(n9249)
         );
  DFF_X1 \REGISTERS_reg[15][36]  ( .D(n6499), .CK(CLK), .Q(n20096), .QN(n9250)
         );
  DFF_X1 \REGISTERS_reg[15][35]  ( .D(n6498), .CK(CLK), .Q(n20097), .QN(n9251)
         );
  DFF_X1 \REGISTERS_reg[15][34]  ( .D(n6497), .CK(CLK), .Q(n20098), .QN(n9252)
         );
  DFF_X1 \REGISTERS_reg[15][33]  ( .D(n6496), .CK(CLK), .Q(n20099), .QN(n9253)
         );
  DFF_X1 \REGISTERS_reg[15][32]  ( .D(n6495), .CK(CLK), .Q(n20100), .QN(n9254)
         );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n6494), .CK(CLK), .Q(n20101), .QN(n9255)
         );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n6493), .CK(CLK), .Q(n20102), .QN(n9256)
         );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n6492), .CK(CLK), .Q(n20103), .QN(n9257)
         );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n6491), .CK(CLK), .Q(n20104), .QN(n9258)
         );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n6490), .CK(CLK), .Q(n20105), .QN(n9259)
         );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n6489), .CK(CLK), .Q(n20106), .QN(n9260)
         );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n6488), .CK(CLK), .Q(n20107), .QN(n9261)
         );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n6487), .CK(CLK), .Q(n20108), .QN(n9262)
         );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n6486), .CK(CLK), .Q(n20109), .QN(n9263)
         );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n6485), .CK(CLK), .Q(n20110), .QN(n9264)
         );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n6484), .CK(CLK), .Q(n20111), .QN(n9265)
         );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n6483), .CK(CLK), .Q(n20112), .QN(n9266)
         );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n6482), .CK(CLK), .Q(n20113), .QN(n9267)
         );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n6481), .CK(CLK), .Q(n20114), .QN(n9268)
         );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n6480), .CK(CLK), .Q(n20115), .QN(n9269)
         );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n6479), .CK(CLK), .Q(n20116), .QN(n9270)
         );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n6478), .CK(CLK), .Q(n20117), .QN(n9271)
         );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n6477), .CK(CLK), .Q(n20118), .QN(n9272)
         );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n6476), .CK(CLK), .Q(n20119), .QN(n9273)
         );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n6475), .CK(CLK), .Q(n20120), .QN(n9274)
         );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n6474), .CK(CLK), .Q(n20121), .QN(n9275)
         );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n6473), .CK(CLK), .Q(n20122), .QN(n9276)
         );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n6472), .CK(CLK), .Q(n20123), .QN(n9277)
         );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n6471), .CK(CLK), .Q(n20124), .QN(n9278)
         );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n6470), .CK(CLK), .Q(n20125), .QN(n9279)
         );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n6469), .CK(CLK), .Q(n20126), .QN(n9280)
         );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n6468), .CK(CLK), .Q(n20127), .QN(n9281)
         );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n6467), .CK(CLK), .Q(n20128), .QN(n9282)
         );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n6466), .CK(CLK), .Q(n20129), .QN(n9283)
         );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n6465), .CK(CLK), .Q(n20130), .QN(n9284)
         );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n6464), .CK(CLK), .Q(n20131), .QN(n9285)
         );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n6463), .CK(CLK), .Q(n20132), .QN(n9286)
         );
  DFF_X1 \REGISTERS_reg[21][63]  ( .D(n6142), .CK(CLK), .QN(n8967) );
  DFF_X1 \REGISTERS_reg[27][63]  ( .D(n5758), .CK(CLK), .QN(n20134) );
  DFF_X1 \REGISTERS_reg[27][62]  ( .D(n5757), .CK(CLK), .QN(n20135) );
  DFF_X1 \REGISTERS_reg[27][61]  ( .D(n5756), .CK(CLK), .QN(n20136) );
  DFF_X1 \REGISTERS_reg[27][60]  ( .D(n5755), .CK(CLK), .QN(n20137) );
  DFF_X1 \REGISTERS_reg[27][59]  ( .D(n5754), .CK(CLK), .QN(n20138) );
  DFF_X1 \REGISTERS_reg[27][58]  ( .D(n5753), .CK(CLK), .QN(n20139) );
  DFF_X1 \REGISTERS_reg[27][57]  ( .D(n5752), .CK(CLK), .QN(n20140) );
  DFF_X1 \REGISTERS_reg[27][56]  ( .D(n5751), .CK(CLK), .QN(n20141) );
  DFF_X1 \REGISTERS_reg[27][55]  ( .D(n5750), .CK(CLK), .QN(n20142) );
  DFF_X1 \REGISTERS_reg[27][54]  ( .D(n5749), .CK(CLK), .QN(n20143) );
  DFF_X1 \REGISTERS_reg[27][53]  ( .D(n5748), .CK(CLK), .QN(n20144) );
  DFF_X1 \REGISTERS_reg[27][52]  ( .D(n5747), .CK(CLK), .QN(n20145) );
  DFF_X1 \REGISTERS_reg[27][51]  ( .D(n5746), .CK(CLK), .QN(n20146) );
  DFF_X1 \REGISTERS_reg[27][50]  ( .D(n5745), .CK(CLK), .QN(n20147) );
  DFF_X1 \REGISTERS_reg[27][49]  ( .D(n5744), .CK(CLK), .QN(n20148) );
  DFF_X1 \REGISTERS_reg[27][48]  ( .D(n5743), .CK(CLK), .QN(n20149) );
  DFF_X1 \REGISTERS_reg[27][47]  ( .D(n5742), .CK(CLK), .QN(n20150) );
  DFF_X1 \REGISTERS_reg[27][46]  ( .D(n5741), .CK(CLK), .QN(n20151) );
  DFF_X1 \REGISTERS_reg[27][45]  ( .D(n5740), .CK(CLK), .QN(n20152) );
  DFF_X1 \REGISTERS_reg[27][44]  ( .D(n5739), .CK(CLK), .QN(n20153) );
  DFF_X1 \REGISTERS_reg[27][43]  ( .D(n5738), .CK(CLK), .QN(n20154) );
  DFF_X1 \REGISTERS_reg[27][42]  ( .D(n5737), .CK(CLK), .QN(n20155) );
  DFF_X1 \REGISTERS_reg[27][41]  ( .D(n5736), .CK(CLK), .QN(n20156) );
  DFF_X1 \REGISTERS_reg[27][40]  ( .D(n5735), .CK(CLK), .QN(n20157) );
  DFF_X1 \REGISTERS_reg[27][39]  ( .D(n5734), .CK(CLK), .QN(n20158) );
  DFF_X1 \REGISTERS_reg[27][38]  ( .D(n5733), .CK(CLK), .QN(n20159) );
  DFF_X1 \REGISTERS_reg[27][37]  ( .D(n5732), .CK(CLK), .QN(n20160) );
  DFF_X1 \REGISTERS_reg[27][36]  ( .D(n5731), .CK(CLK), .QN(n20161) );
  DFF_X1 \REGISTERS_reg[27][35]  ( .D(n5730), .CK(CLK), .QN(n20162) );
  DFF_X1 \REGISTERS_reg[27][34]  ( .D(n5729), .CK(CLK), .QN(n20163) );
  DFF_X1 \REGISTERS_reg[27][33]  ( .D(n5728), .CK(CLK), .QN(n20164) );
  DFF_X1 \REGISTERS_reg[27][32]  ( .D(n5727), .CK(CLK), .QN(n20165) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n5726), .CK(CLK), .QN(n20166) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n5725), .CK(CLK), .QN(n20167) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n5724), .CK(CLK), .QN(n20168) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n5723), .CK(CLK), .QN(n20169) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n5722), .CK(CLK), .QN(n20170) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n5721), .CK(CLK), .QN(n20171) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n5720), .CK(CLK), .QN(n20172) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n5719), .CK(CLK), .QN(n20173) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n5718), .CK(CLK), .QN(n20174) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n5717), .CK(CLK), .QN(n20175) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n5716), .CK(CLK), .QN(n20176) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n5715), .CK(CLK), .QN(n20177) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n5714), .CK(CLK), .QN(n20178) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n5713), .CK(CLK), .QN(n20179) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n5712), .CK(CLK), .QN(n20180) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n5711), .CK(CLK), .QN(n20181) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n5710), .CK(CLK), .QN(n20182) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n5709), .CK(CLK), .QN(n20183) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n5708), .CK(CLK), .QN(n20184) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n5707), .CK(CLK), .QN(n20185) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n5706), .CK(CLK), .QN(n20186) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n5705), .CK(CLK), .QN(n20187) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n5704), .CK(CLK), .QN(n20188) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n5703), .CK(CLK), .QN(n20189) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n5702), .CK(CLK), .QN(n20190) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n5701), .CK(CLK), .QN(n20191) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n5700), .CK(CLK), .QN(n20192) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n5699), .CK(CLK), .QN(n20193) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n5698), .CK(CLK), .QN(n20194) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n5697), .CK(CLK), .QN(n20195) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n5696), .CK(CLK), .QN(n20196) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n5695), .CK(CLK), .QN(n20197) );
  DFF_X1 \REGISTERS_reg[5][63]  ( .D(n7166), .CK(CLK), .QN(n19558) );
  DFF_X1 \REGISTERS_reg[5][62]  ( .D(n7165), .CK(CLK), .QN(n19559) );
  DFF_X1 \REGISTERS_reg[5][61]  ( .D(n7164), .CK(CLK), .QN(n19560) );
  DFF_X1 \REGISTERS_reg[5][60]  ( .D(n7163), .CK(CLK), .QN(n19561) );
  DFF_X1 \REGISTERS_reg[5][59]  ( .D(n7162), .CK(CLK), .QN(n19562) );
  DFF_X1 \REGISTERS_reg[5][58]  ( .D(n7161), .CK(CLK), .QN(n19563) );
  DFF_X1 \REGISTERS_reg[5][57]  ( .D(n7160), .CK(CLK), .QN(n19564) );
  DFF_X1 \REGISTERS_reg[5][56]  ( .D(n7159), .CK(CLK), .QN(n19565) );
  DFF_X1 \REGISTERS_reg[5][55]  ( .D(n7158), .CK(CLK), .QN(n19566) );
  DFF_X1 \REGISTERS_reg[5][54]  ( .D(n7157), .CK(CLK), .QN(n19567) );
  DFF_X1 \REGISTERS_reg[5][53]  ( .D(n7156), .CK(CLK), .QN(n19568) );
  DFF_X1 \REGISTERS_reg[5][52]  ( .D(n7155), .CK(CLK), .QN(n19569) );
  DFF_X1 \REGISTERS_reg[5][51]  ( .D(n7154), .CK(CLK), .QN(n19570) );
  DFF_X1 \REGISTERS_reg[5][50]  ( .D(n7153), .CK(CLK), .QN(n19571) );
  DFF_X1 \REGISTERS_reg[5][49]  ( .D(n7152), .CK(CLK), .QN(n19572) );
  DFF_X1 \REGISTERS_reg[5][48]  ( .D(n7151), .CK(CLK), .QN(n19573) );
  DFF_X1 \REGISTERS_reg[5][47]  ( .D(n7150), .CK(CLK), .QN(n19574) );
  DFF_X1 \REGISTERS_reg[5][46]  ( .D(n7149), .CK(CLK), .QN(n19575) );
  DFF_X1 \REGISTERS_reg[5][45]  ( .D(n7148), .CK(CLK), .QN(n19576) );
  DFF_X1 \REGISTERS_reg[5][44]  ( .D(n7147), .CK(CLK), .QN(n19577) );
  DFF_X1 \REGISTERS_reg[5][43]  ( .D(n7146), .CK(CLK), .QN(n19578) );
  DFF_X1 \REGISTERS_reg[5][42]  ( .D(n7145), .CK(CLK), .QN(n19579) );
  DFF_X1 \REGISTERS_reg[5][41]  ( .D(n7144), .CK(CLK), .QN(n19580) );
  DFF_X1 \REGISTERS_reg[5][40]  ( .D(n7143), .CK(CLK), .QN(n19581) );
  DFF_X1 \REGISTERS_reg[5][39]  ( .D(n7142), .CK(CLK), .QN(n19582) );
  DFF_X1 \REGISTERS_reg[5][38]  ( .D(n7141), .CK(CLK), .QN(n19583) );
  DFF_X1 \REGISTERS_reg[5][37]  ( .D(n7140), .CK(CLK), .QN(n19584) );
  DFF_X1 \REGISTERS_reg[5][36]  ( .D(n7139), .CK(CLK), .QN(n19585) );
  DFF_X1 \REGISTERS_reg[5][35]  ( .D(n7138), .CK(CLK), .QN(n19586) );
  DFF_X1 \REGISTERS_reg[5][34]  ( .D(n7137), .CK(CLK), .QN(n19587) );
  DFF_X1 \REGISTERS_reg[5][33]  ( .D(n7136), .CK(CLK), .QN(n19588) );
  DFF_X1 \REGISTERS_reg[5][32]  ( .D(n7135), .CK(CLK), .QN(n19589) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n7134), .CK(CLK), .QN(n19590) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n7133), .CK(CLK), .QN(n19591) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n7132), .CK(CLK), .QN(n19592) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n7131), .CK(CLK), .QN(n19593) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n7130), .CK(CLK), .QN(n19594) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n7129), .CK(CLK), .QN(n19595) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n7128), .CK(CLK), .QN(n19596) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n7127), .CK(CLK), .QN(n19597) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n7126), .CK(CLK), .QN(n19598) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n7125), .CK(CLK), .QN(n19599) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n7124), .CK(CLK), .QN(n19600) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n7123), .CK(CLK), .QN(n19601) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n7122), .CK(CLK), .QN(n19602) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n7121), .CK(CLK), .QN(n19603) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n7120), .CK(CLK), .QN(n19604) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n7119), .CK(CLK), .QN(n19605) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n7118), .CK(CLK), .QN(n19606) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n7117), .CK(CLK), .QN(n19607) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n7116), .CK(CLK), .QN(n19608) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n7115), .CK(CLK), .QN(n19609) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n7114), .CK(CLK), .QN(n19610) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n7113), .CK(CLK), .QN(n19611) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n7112), .CK(CLK), .QN(n19612) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n7111), .CK(CLK), .QN(n19613) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n7110), .CK(CLK), .QN(n19614) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n7109), .CK(CLK), .QN(n19615) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n7108), .CK(CLK), .QN(n19616) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n7107), .CK(CLK), .QN(n19617) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n7106), .CK(CLK), .QN(n19618) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n7105), .CK(CLK), .QN(n19619) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n7104), .CK(CLK), .QN(n19620) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n7103), .CK(CLK), .QN(n19621) );
  DFF_X1 \REGISTERS_reg[1][63]  ( .D(n7422), .CK(CLK), .QN(n20966) );
  DFF_X1 \REGISTERS_reg[1][62]  ( .D(n7421), .CK(CLK), .QN(n20967) );
  DFF_X1 \REGISTERS_reg[1][61]  ( .D(n7420), .CK(CLK), .QN(n20968) );
  DFF_X1 \REGISTERS_reg[1][60]  ( .D(n7419), .CK(CLK), .QN(n20969) );
  DFF_X1 \REGISTERS_reg[1][59]  ( .D(n7418), .CK(CLK), .QN(n20970) );
  DFF_X1 \REGISTERS_reg[1][58]  ( .D(n7417), .CK(CLK), .QN(n20971) );
  DFF_X1 \REGISTERS_reg[1][57]  ( .D(n7416), .CK(CLK), .QN(n20972) );
  DFF_X1 \REGISTERS_reg[1][56]  ( .D(n7415), .CK(CLK), .QN(n20973) );
  DFF_X1 \REGISTERS_reg[1][55]  ( .D(n7414), .CK(CLK), .QN(n20974) );
  DFF_X1 \REGISTERS_reg[1][54]  ( .D(n7413), .CK(CLK), .QN(n20975) );
  DFF_X1 \REGISTERS_reg[1][53]  ( .D(n7412), .CK(CLK), .QN(n20976) );
  DFF_X1 \REGISTERS_reg[1][52]  ( .D(n7411), .CK(CLK), .QN(n20977) );
  DFF_X1 \REGISTERS_reg[1][51]  ( .D(n7410), .CK(CLK), .QN(n20978) );
  DFF_X1 \REGISTERS_reg[1][50]  ( .D(n7409), .CK(CLK), .QN(n20979) );
  DFF_X1 \REGISTERS_reg[1][49]  ( .D(n7408), .CK(CLK), .QN(n20980) );
  DFF_X1 \REGISTERS_reg[1][48]  ( .D(n7407), .CK(CLK), .QN(n20981) );
  DFF_X1 \REGISTERS_reg[1][47]  ( .D(n7406), .CK(CLK), .QN(n20982) );
  DFF_X1 \REGISTERS_reg[1][46]  ( .D(n7405), .CK(CLK), .QN(n20983) );
  DFF_X1 \REGISTERS_reg[1][45]  ( .D(n7404), .CK(CLK), .QN(n20984) );
  DFF_X1 \REGISTERS_reg[1][44]  ( .D(n7403), .CK(CLK), .QN(n20985) );
  DFF_X1 \REGISTERS_reg[1][43]  ( .D(n7402), .CK(CLK), .QN(n20986) );
  DFF_X1 \REGISTERS_reg[1][42]  ( .D(n7401), .CK(CLK), .QN(n20987) );
  DFF_X1 \REGISTERS_reg[1][41]  ( .D(n7400), .CK(CLK), .QN(n20988) );
  DFF_X1 \REGISTERS_reg[1][40]  ( .D(n7399), .CK(CLK), .QN(n20989) );
  DFF_X1 \REGISTERS_reg[1][39]  ( .D(n7398), .CK(CLK), .QN(n20990) );
  DFF_X1 \REGISTERS_reg[1][38]  ( .D(n7397), .CK(CLK), .QN(n20991) );
  DFF_X1 \REGISTERS_reg[1][37]  ( .D(n7396), .CK(CLK), .QN(n20992) );
  DFF_X1 \REGISTERS_reg[1][36]  ( .D(n7395), .CK(CLK), .QN(n20993) );
  DFF_X1 \REGISTERS_reg[1][35]  ( .D(n7394), .CK(CLK), .QN(n20994) );
  DFF_X1 \REGISTERS_reg[1][34]  ( .D(n7393), .CK(CLK), .QN(n20995) );
  DFF_X1 \REGISTERS_reg[1][33]  ( .D(n7392), .CK(CLK), .QN(n20996) );
  DFF_X1 \REGISTERS_reg[1][32]  ( .D(n7391), .CK(CLK), .QN(n20997) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n7390), .CK(CLK), .QN(n20998) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n7389), .CK(CLK), .QN(n20999) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n7388), .CK(CLK), .QN(n21000) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n7387), .CK(CLK), .QN(n21001) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n7386), .CK(CLK), .QN(n21002) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n7385), .CK(CLK), .QN(n21003) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n7384), .CK(CLK), .QN(n21004) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n7383), .CK(CLK), .QN(n21005) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n7382), .CK(CLK), .QN(n21006) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n7381), .CK(CLK), .QN(n21007) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n7380), .CK(CLK), .QN(n21008) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n7379), .CK(CLK), .QN(n21009) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n7378), .CK(CLK), .QN(n21010) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n7377), .CK(CLK), .QN(n21011) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n7376), .CK(CLK), .QN(n21012) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n7375), .CK(CLK), .QN(n21013) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n7374), .CK(CLK), .QN(n21014) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n7373), .CK(CLK), .QN(n21015) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n7372), .CK(CLK), .QN(n21016) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n7371), .CK(CLK), .QN(n21017) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n7370), .CK(CLK), .QN(n21018) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n7369), .CK(CLK), .QN(n21019) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n7368), .CK(CLK), .QN(n21020) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n7367), .CK(CLK), .QN(n21021) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n7366), .CK(CLK), .QN(n21022) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n7365), .CK(CLK), .QN(n21023) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n7364), .CK(CLK), .QN(n21024) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n7363), .CK(CLK), .QN(n21025) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n7362), .CK(CLK), .QN(n21026) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n7361), .CK(CLK), .QN(n21027) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n7360), .CK(CLK), .QN(n21028) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n7359), .CK(CLK), .QN(n21029) );
  DFF_X1 \REGISTERS_reg[20][63]  ( .D(n6206), .CK(CLK), .QN(n20270) );
  DFF_X1 \REGISTERS_reg[20][62]  ( .D(n6205), .CK(CLK), .QN(n20271) );
  DFF_X1 \REGISTERS_reg[20][61]  ( .D(n6204), .CK(CLK), .QN(n20272) );
  DFF_X1 \REGISTERS_reg[20][60]  ( .D(n6203), .CK(CLK), .QN(n20273) );
  DFF_X1 \REGISTERS_reg[20][59]  ( .D(n6202), .CK(CLK), .QN(n20274) );
  DFF_X1 \REGISTERS_reg[20][58]  ( .D(n6201), .CK(CLK), .QN(n20275) );
  DFF_X1 \REGISTERS_reg[20][57]  ( .D(n6200), .CK(CLK), .QN(n20276) );
  DFF_X1 \REGISTERS_reg[20][56]  ( .D(n6199), .CK(CLK), .QN(n20277) );
  DFF_X1 \REGISTERS_reg[20][55]  ( .D(n6198), .CK(CLK), .QN(n20278) );
  DFF_X1 \REGISTERS_reg[20][54]  ( .D(n6197), .CK(CLK), .QN(n20279) );
  DFF_X1 \REGISTERS_reg[20][53]  ( .D(n6196), .CK(CLK), .QN(n20280) );
  DFF_X1 \REGISTERS_reg[20][52]  ( .D(n6195), .CK(CLK), .QN(n20281) );
  DFF_X1 \REGISTERS_reg[20][51]  ( .D(n6194), .CK(CLK), .QN(n20282) );
  DFF_X1 \REGISTERS_reg[20][50]  ( .D(n6193), .CK(CLK), .QN(n20283) );
  DFF_X1 \REGISTERS_reg[20][49]  ( .D(n6192), .CK(CLK), .QN(n20284) );
  DFF_X1 \REGISTERS_reg[20][48]  ( .D(n6191), .CK(CLK), .QN(n20285) );
  DFF_X1 \REGISTERS_reg[20][47]  ( .D(n6190), .CK(CLK), .QN(n20286) );
  DFF_X1 \REGISTERS_reg[20][46]  ( .D(n6189), .CK(CLK), .QN(n20287) );
  DFF_X1 \REGISTERS_reg[20][45]  ( .D(n6188), .CK(CLK), .QN(n20288) );
  DFF_X1 \REGISTERS_reg[20][44]  ( .D(n6187), .CK(CLK), .QN(n20289) );
  DFF_X1 \REGISTERS_reg[20][43]  ( .D(n6186), .CK(CLK), .QN(n20290) );
  DFF_X1 \REGISTERS_reg[20][42]  ( .D(n6185), .CK(CLK), .QN(n20291) );
  DFF_X1 \REGISTERS_reg[20][41]  ( .D(n6184), .CK(CLK), .QN(n20292) );
  DFF_X1 \REGISTERS_reg[20][40]  ( .D(n6183), .CK(CLK), .QN(n20293) );
  DFF_X1 \REGISTERS_reg[20][39]  ( .D(n6182), .CK(CLK), .QN(n20294) );
  DFF_X1 \REGISTERS_reg[20][38]  ( .D(n6181), .CK(CLK), .QN(n20295) );
  DFF_X1 \REGISTERS_reg[20][37]  ( .D(n6180), .CK(CLK), .QN(n20296) );
  DFF_X1 \REGISTERS_reg[20][36]  ( .D(n6179), .CK(CLK), .QN(n20297) );
  DFF_X1 \REGISTERS_reg[20][35]  ( .D(n6178), .CK(CLK), .QN(n20298) );
  DFF_X1 \REGISTERS_reg[20][34]  ( .D(n6177), .CK(CLK), .QN(n20299) );
  DFF_X1 \REGISTERS_reg[20][33]  ( .D(n6176), .CK(CLK), .QN(n20300) );
  DFF_X1 \REGISTERS_reg[20][32]  ( .D(n6175), .CK(CLK), .QN(n20301) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n6174), .CK(CLK), .QN(n20302) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n6173), .CK(CLK), .QN(n20303) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n6172), .CK(CLK), .QN(n20304) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n6171), .CK(CLK), .QN(n20305) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n6170), .CK(CLK), .QN(n20306) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n6169), .CK(CLK), .QN(n20307) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n6168), .CK(CLK), .QN(n20308) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n6167), .CK(CLK), .QN(n20309) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n6166), .CK(CLK), .QN(n20310) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n6165), .CK(CLK), .QN(n20311) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n6164), .CK(CLK), .QN(n20312) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n6163), .CK(CLK), .QN(n20313) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n6162), .CK(CLK), .QN(n20314) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n6161), .CK(CLK), .QN(n20315) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n6160), .CK(CLK), .QN(n20316) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n6159), .CK(CLK), .QN(n20317) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n6158), .CK(CLK), .QN(n20318) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n6157), .CK(CLK), .QN(n20319) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n6156), .CK(CLK), .QN(n20320) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n6155), .CK(CLK), .QN(n20321) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n6154), .CK(CLK), .QN(n20322) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n6153), .CK(CLK), .QN(n20323) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n6152), .CK(CLK), .QN(n20324) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n6151), .CK(CLK), .QN(n20325) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n6150), .CK(CLK), .QN(n20326) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n6149), .CK(CLK), .QN(n20327) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n6148), .CK(CLK), .QN(n20328) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n6147), .CK(CLK), .QN(n20329) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n6146), .CK(CLK), .QN(n20330) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n6145), .CK(CLK), .QN(n20331) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n6144), .CK(CLK), .QN(n20332) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n6143), .CK(CLK), .QN(n20333) );
  DFF_X1 \REGISTERS_reg[18][63]  ( .D(n6334), .CK(CLK), .QN(n20334) );
  DFF_X1 \REGISTERS_reg[18][62]  ( .D(n6333), .CK(CLK), .QN(n20335) );
  DFF_X1 \REGISTERS_reg[18][61]  ( .D(n6332), .CK(CLK), .QN(n20336) );
  DFF_X1 \REGISTERS_reg[18][60]  ( .D(n6331), .CK(CLK), .QN(n20337) );
  DFF_X1 \REGISTERS_reg[18][59]  ( .D(n6330), .CK(CLK), .QN(n20338) );
  DFF_X1 \REGISTERS_reg[18][58]  ( .D(n6329), .CK(CLK), .QN(n20339) );
  DFF_X1 \REGISTERS_reg[18][57]  ( .D(n6328), .CK(CLK), .QN(n20340) );
  DFF_X1 \REGISTERS_reg[18][56]  ( .D(n6327), .CK(CLK), .QN(n20341) );
  DFF_X1 \REGISTERS_reg[18][55]  ( .D(n6326), .CK(CLK), .QN(n20342) );
  DFF_X1 \REGISTERS_reg[18][54]  ( .D(n6325), .CK(CLK), .QN(n20343) );
  DFF_X1 \REGISTERS_reg[18][53]  ( .D(n6324), .CK(CLK), .QN(n20344) );
  DFF_X1 \REGISTERS_reg[18][52]  ( .D(n6323), .CK(CLK), .QN(n20345) );
  DFF_X1 \REGISTERS_reg[18][51]  ( .D(n6322), .CK(CLK), .QN(n20346) );
  DFF_X1 \REGISTERS_reg[18][50]  ( .D(n6321), .CK(CLK), .QN(n20347) );
  DFF_X1 \REGISTERS_reg[18][49]  ( .D(n6320), .CK(CLK), .QN(n20348) );
  DFF_X1 \REGISTERS_reg[18][48]  ( .D(n6319), .CK(CLK), .QN(n20349) );
  DFF_X1 \REGISTERS_reg[18][47]  ( .D(n6318), .CK(CLK), .QN(n20350) );
  DFF_X1 \REGISTERS_reg[18][46]  ( .D(n6317), .CK(CLK), .QN(n20351) );
  DFF_X1 \REGISTERS_reg[18][45]  ( .D(n6316), .CK(CLK), .QN(n20352) );
  DFF_X1 \REGISTERS_reg[18][44]  ( .D(n6315), .CK(CLK), .QN(n20353) );
  DFF_X1 \REGISTERS_reg[18][43]  ( .D(n6314), .CK(CLK), .QN(n20354) );
  DFF_X1 \REGISTERS_reg[18][42]  ( .D(n6313), .CK(CLK), .QN(n20355) );
  DFF_X1 \REGISTERS_reg[18][41]  ( .D(n6312), .CK(CLK), .QN(n20356) );
  DFF_X1 \REGISTERS_reg[18][40]  ( .D(n6311), .CK(CLK), .QN(n20357) );
  DFF_X1 \REGISTERS_reg[18][39]  ( .D(n6310), .CK(CLK), .QN(n20358) );
  DFF_X1 \REGISTERS_reg[18][38]  ( .D(n6309), .CK(CLK), .QN(n20359) );
  DFF_X1 \REGISTERS_reg[18][37]  ( .D(n6308), .CK(CLK), .QN(n20360) );
  DFF_X1 \REGISTERS_reg[18][36]  ( .D(n6307), .CK(CLK), .QN(n20361) );
  DFF_X1 \REGISTERS_reg[18][35]  ( .D(n6306), .CK(CLK), .QN(n20362) );
  DFF_X1 \REGISTERS_reg[18][34]  ( .D(n6305), .CK(CLK), .QN(n20363) );
  DFF_X1 \REGISTERS_reg[18][33]  ( .D(n6304), .CK(CLK), .QN(n20364) );
  DFF_X1 \REGISTERS_reg[18][32]  ( .D(n6303), .CK(CLK), .QN(n20365) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n6302), .CK(CLK), .QN(n20366) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n6301), .CK(CLK), .QN(n20367) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n6300), .CK(CLK), .QN(n20368) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n6299), .CK(CLK), .QN(n20369) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n6298), .CK(CLK), .QN(n20370) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n6297), .CK(CLK), .QN(n20371) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n6296), .CK(CLK), .QN(n20372) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n6295), .CK(CLK), .QN(n20373) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n6294), .CK(CLK), .QN(n20374) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n6293), .CK(CLK), .QN(n20375) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n6292), .CK(CLK), .QN(n20376) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n6291), .CK(CLK), .QN(n20377) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n6290), .CK(CLK), .QN(n20378) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n6289), .CK(CLK), .QN(n20379) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n6288), .CK(CLK), .QN(n20380) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n6287), .CK(CLK), .QN(n20381) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n6286), .CK(CLK), .QN(n20382) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n6285), .CK(CLK), .QN(n20383) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n6284), .CK(CLK), .QN(n20384) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n6283), .CK(CLK), .QN(n20385) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n6282), .CK(CLK), .QN(n20386) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n6281), .CK(CLK), .QN(n20387) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n6280), .CK(CLK), .QN(n20388) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n6279), .CK(CLK), .QN(n20389) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n6278), .CK(CLK), .QN(n20390) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n6277), .CK(CLK), .QN(n20391) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n6276), .CK(CLK), .QN(n20392) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n6275), .CK(CLK), .QN(n20393) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n6274), .CK(CLK), .QN(n20394) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n6273), .CK(CLK), .QN(n20395) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n6272), .CK(CLK), .QN(n20396) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n6271), .CK(CLK), .QN(n20397) );
  DFF_X1 \REGISTERS_reg[13][63]  ( .D(n6654), .CK(CLK), .QN(n19813) );
  DFF_X1 \REGISTERS_reg[13][62]  ( .D(n6653), .CK(CLK), .QN(n19814) );
  DFF_X1 \REGISTERS_reg[13][61]  ( .D(n6652), .CK(CLK), .QN(n19815) );
  DFF_X1 \REGISTERS_reg[13][60]  ( .D(n6651), .CK(CLK), .QN(n19816) );
  DFF_X1 \REGISTERS_reg[13][59]  ( .D(n6650), .CK(CLK), .QN(n19817) );
  DFF_X1 \REGISTERS_reg[13][58]  ( .D(n6649), .CK(CLK), .QN(n19818) );
  DFF_X1 \REGISTERS_reg[13][57]  ( .D(n6648), .CK(CLK), .QN(n19819) );
  DFF_X1 \REGISTERS_reg[13][56]  ( .D(n6647), .CK(CLK), .QN(n19820) );
  DFF_X1 \REGISTERS_reg[13][55]  ( .D(n6646), .CK(CLK), .QN(n19821) );
  DFF_X1 \REGISTERS_reg[13][54]  ( .D(n6645), .CK(CLK), .QN(n19822) );
  DFF_X1 \REGISTERS_reg[13][53]  ( .D(n6644), .CK(CLK), .QN(n19823) );
  DFF_X1 \REGISTERS_reg[13][52]  ( .D(n6643), .CK(CLK), .QN(n19824) );
  DFF_X1 \REGISTERS_reg[13][51]  ( .D(n6642), .CK(CLK), .QN(n19825) );
  DFF_X1 \REGISTERS_reg[13][50]  ( .D(n6641), .CK(CLK), .QN(n19826) );
  DFF_X1 \REGISTERS_reg[13][49]  ( .D(n6640), .CK(CLK), .QN(n19827) );
  DFF_X1 \REGISTERS_reg[13][48]  ( .D(n6639), .CK(CLK), .QN(n19828) );
  DFF_X1 \REGISTERS_reg[13][47]  ( .D(n6638), .CK(CLK), .QN(n19829) );
  DFF_X1 \REGISTERS_reg[13][46]  ( .D(n6637), .CK(CLK), .QN(n19830) );
  DFF_X1 \REGISTERS_reg[13][45]  ( .D(n6636), .CK(CLK), .QN(n19831) );
  DFF_X1 \REGISTERS_reg[13][44]  ( .D(n6635), .CK(CLK), .QN(n19832) );
  DFF_X1 \REGISTERS_reg[13][43]  ( .D(n6634), .CK(CLK), .QN(n19833) );
  DFF_X1 \REGISTERS_reg[13][42]  ( .D(n6633), .CK(CLK), .QN(n19834) );
  DFF_X1 \REGISTERS_reg[13][41]  ( .D(n6632), .CK(CLK), .QN(n19835) );
  DFF_X1 \REGISTERS_reg[13][40]  ( .D(n6631), .CK(CLK), .QN(n19836) );
  DFF_X1 \REGISTERS_reg[13][39]  ( .D(n6630), .CK(CLK), .QN(n19837) );
  DFF_X1 \REGISTERS_reg[13][38]  ( .D(n6629), .CK(CLK), .QN(n19838) );
  DFF_X1 \REGISTERS_reg[13][37]  ( .D(n6628), .CK(CLK), .QN(n19839) );
  DFF_X1 \REGISTERS_reg[13][36]  ( .D(n6627), .CK(CLK), .QN(n19840) );
  DFF_X1 \REGISTERS_reg[13][35]  ( .D(n6626), .CK(CLK), .QN(n19841) );
  DFF_X1 \REGISTERS_reg[13][34]  ( .D(n6625), .CK(CLK), .QN(n19842) );
  DFF_X1 \REGISTERS_reg[13][33]  ( .D(n6624), .CK(CLK), .QN(n19843) );
  DFF_X1 \REGISTERS_reg[13][32]  ( .D(n6623), .CK(CLK), .QN(n19844) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n6622), .CK(CLK), .QN(n19845) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n6621), .CK(CLK), .QN(n19846) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n6620), .CK(CLK), .QN(n19847) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n6619), .CK(CLK), .QN(n19848) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n6618), .CK(CLK), .QN(n19849) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n6617), .CK(CLK), .QN(n19850) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n6616), .CK(CLK), .QN(n19851) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n6615), .CK(CLK), .QN(n19852) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n6614), .CK(CLK), .QN(n19853) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n6613), .CK(CLK), .QN(n19854) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n6612), .CK(CLK), .QN(n19855) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n6611), .CK(CLK), .QN(n19856) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n6610), .CK(CLK), .QN(n19857) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n6609), .CK(CLK), .QN(n19858) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n6608), .CK(CLK), .QN(n19859) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n6607), .CK(CLK), .QN(n19860) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n6606), .CK(CLK), .QN(n19861) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n6605), .CK(CLK), .QN(n19862) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n6604), .CK(CLK), .QN(n19863) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n6603), .CK(CLK), .QN(n19864) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n6602), .CK(CLK), .QN(n19865) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n6601), .CK(CLK), .QN(n19866) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n6600), .CK(CLK), .QN(n19867) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n6599), .CK(CLK), .QN(n19868) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n6598), .CK(CLK), .QN(n19869) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n6597), .CK(CLK), .QN(n19870) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n6596), .CK(CLK), .QN(n19871) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n6595), .CK(CLK), .QN(n19872) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n6594), .CK(CLK), .QN(n19873) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n6593), .CK(CLK), .QN(n19874) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n6592), .CK(CLK), .QN(n19875) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n6591), .CK(CLK), .QN(n19876) );
  DFF_X1 \REGISTERS_reg[12][63]  ( .D(n6718), .CK(CLK), .QN(n20398) );
  DFF_X1 \REGISTERS_reg[12][62]  ( .D(n6717), .CK(CLK), .QN(n20399) );
  DFF_X1 \REGISTERS_reg[12][61]  ( .D(n6716), .CK(CLK), .QN(n20400) );
  DFF_X1 \REGISTERS_reg[12][60]  ( .D(n6715), .CK(CLK), .QN(n20401) );
  DFF_X1 \REGISTERS_reg[12][59]  ( .D(n6714), .CK(CLK), .QN(n20402) );
  DFF_X1 \REGISTERS_reg[12][58]  ( .D(n6713), .CK(CLK), .QN(n20403) );
  DFF_X1 \REGISTERS_reg[12][57]  ( .D(n6712), .CK(CLK), .QN(n20404) );
  DFF_X1 \REGISTERS_reg[12][56]  ( .D(n6711), .CK(CLK), .QN(n20405) );
  DFF_X1 \REGISTERS_reg[12][55]  ( .D(n6710), .CK(CLK), .QN(n20406) );
  DFF_X1 \REGISTERS_reg[12][54]  ( .D(n6709), .CK(CLK), .QN(n20407) );
  DFF_X1 \REGISTERS_reg[12][53]  ( .D(n6708), .CK(CLK), .QN(n20408) );
  DFF_X1 \REGISTERS_reg[12][52]  ( .D(n6707), .CK(CLK), .QN(n20409) );
  DFF_X1 \REGISTERS_reg[12][51]  ( .D(n6706), .CK(CLK), .QN(n20410) );
  DFF_X1 \REGISTERS_reg[12][50]  ( .D(n6705), .CK(CLK), .QN(n20411) );
  DFF_X1 \REGISTERS_reg[12][49]  ( .D(n6704), .CK(CLK), .QN(n20412) );
  DFF_X1 \REGISTERS_reg[12][48]  ( .D(n6703), .CK(CLK), .QN(n20413) );
  DFF_X1 \REGISTERS_reg[12][47]  ( .D(n6702), .CK(CLK), .QN(n20414) );
  DFF_X1 \REGISTERS_reg[12][46]  ( .D(n6701), .CK(CLK), .QN(n20415) );
  DFF_X1 \REGISTERS_reg[12][45]  ( .D(n6700), .CK(CLK), .QN(n20416) );
  DFF_X1 \REGISTERS_reg[12][44]  ( .D(n6699), .CK(CLK), .QN(n20417) );
  DFF_X1 \REGISTERS_reg[12][43]  ( .D(n6698), .CK(CLK), .QN(n20418) );
  DFF_X1 \REGISTERS_reg[12][42]  ( .D(n6697), .CK(CLK), .QN(n20419) );
  DFF_X1 \REGISTERS_reg[12][41]  ( .D(n6696), .CK(CLK), .QN(n20420) );
  DFF_X1 \REGISTERS_reg[12][40]  ( .D(n6695), .CK(CLK), .QN(n20421) );
  DFF_X1 \REGISTERS_reg[12][39]  ( .D(n6694), .CK(CLK), .QN(n20422) );
  DFF_X1 \REGISTERS_reg[12][38]  ( .D(n6693), .CK(CLK), .QN(n20423) );
  DFF_X1 \REGISTERS_reg[12][37]  ( .D(n6692), .CK(CLK), .QN(n20424) );
  DFF_X1 \REGISTERS_reg[12][36]  ( .D(n6691), .CK(CLK), .QN(n20425) );
  DFF_X1 \REGISTERS_reg[12][35]  ( .D(n6690), .CK(CLK), .QN(n20426) );
  DFF_X1 \REGISTERS_reg[12][34]  ( .D(n6689), .CK(CLK), .QN(n20427) );
  DFF_X1 \REGISTERS_reg[12][33]  ( .D(n6688), .CK(CLK), .QN(n20428) );
  DFF_X1 \REGISTERS_reg[12][32]  ( .D(n6687), .CK(CLK), .QN(n20429) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n6686), .CK(CLK), .QN(n20430) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n6685), .CK(CLK), .QN(n20431) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n6684), .CK(CLK), .QN(n20432) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n6683), .CK(CLK), .QN(n20433) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n6682), .CK(CLK), .QN(n20434) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n6681), .CK(CLK), .QN(n20435) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n6680), .CK(CLK), .QN(n20436) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n6679), .CK(CLK), .QN(n20437) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n6678), .CK(CLK), .QN(n20438) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n6677), .CK(CLK), .QN(n20439) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n6676), .CK(CLK), .QN(n20440) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n6675), .CK(CLK), .QN(n20441) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n6674), .CK(CLK), .QN(n20442) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n6673), .CK(CLK), .QN(n20443) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n6672), .CK(CLK), .QN(n20444) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n6671), .CK(CLK), .QN(n20445) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n6670), .CK(CLK), .QN(n20446) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n6669), .CK(CLK), .QN(n20447) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n6668), .CK(CLK), .QN(n20448) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n6667), .CK(CLK), .QN(n20449) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n6666), .CK(CLK), .QN(n20450) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n6665), .CK(CLK), .QN(n20451) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n6664), .CK(CLK), .QN(n20452) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n6663), .CK(CLK), .QN(n20453) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n6662), .CK(CLK), .QN(n20454) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n6661), .CK(CLK), .QN(n20455) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n6660), .CK(CLK), .QN(n20456) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n6659), .CK(CLK), .QN(n20457) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n6658), .CK(CLK), .QN(n20458) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n6657), .CK(CLK), .QN(n20459) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n6656), .CK(CLK), .QN(n20460) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n6655), .CK(CLK), .QN(n20461) );
  DFF_X1 \REGISTERS_reg[29][63]  ( .D(n5630), .CK(CLK), .QN(n21094) );
  DFF_X1 \REGISTERS_reg[29][62]  ( .D(n5629), .CK(CLK), .QN(n21095) );
  DFF_X1 \REGISTERS_reg[29][61]  ( .D(n5628), .CK(CLK), .QN(n21096) );
  DFF_X1 \REGISTERS_reg[29][60]  ( .D(n5627), .CK(CLK), .QN(n21097) );
  DFF_X1 \REGISTERS_reg[26][63]  ( .D(n5822), .CK(CLK), .QN(n21098) );
  DFF_X1 \REGISTERS_reg[26][62]  ( .D(n5821), .CK(CLK), .QN(n21099) );
  DFF_X1 \REGISTERS_reg[26][61]  ( .D(n5820), .CK(CLK), .QN(n21100) );
  DFF_X1 \REGISTERS_reg[26][60]  ( .D(n5819), .CK(CLK), .QN(n21101) );
  DFF_X1 \REGISTERS_reg[29][59]  ( .D(n5626), .CK(CLK), .QN(n21102) );
  DFF_X1 \REGISTERS_reg[29][58]  ( .D(n5625), .CK(CLK), .QN(n21103) );
  DFF_X1 \REGISTERS_reg[29][57]  ( .D(n5624), .CK(CLK), .QN(n21104) );
  DFF_X1 \REGISTERS_reg[29][56]  ( .D(n5623), .CK(CLK), .QN(n21105) );
  DFF_X1 \REGISTERS_reg[29][55]  ( .D(n5622), .CK(CLK), .QN(n21106) );
  DFF_X1 \REGISTERS_reg[29][54]  ( .D(n5621), .CK(CLK), .QN(n21107) );
  DFF_X1 \REGISTERS_reg[29][53]  ( .D(n5620), .CK(CLK), .QN(n21108) );
  DFF_X1 \REGISTERS_reg[29][52]  ( .D(n5619), .CK(CLK), .QN(n21109) );
  DFF_X1 \REGISTERS_reg[29][51]  ( .D(n5618), .CK(CLK), .QN(n21110) );
  DFF_X1 \REGISTERS_reg[29][50]  ( .D(n5617), .CK(CLK), .QN(n21111) );
  DFF_X1 \REGISTERS_reg[29][49]  ( .D(n5616), .CK(CLK), .QN(n21112) );
  DFF_X1 \REGISTERS_reg[29][48]  ( .D(n5615), .CK(CLK), .QN(n21113) );
  DFF_X1 \REGISTERS_reg[29][47]  ( .D(n5614), .CK(CLK), .QN(n21114) );
  DFF_X1 \REGISTERS_reg[29][46]  ( .D(n5613), .CK(CLK), .QN(n21115) );
  DFF_X1 \REGISTERS_reg[29][45]  ( .D(n5612), .CK(CLK), .QN(n21116) );
  DFF_X1 \REGISTERS_reg[29][44]  ( .D(n5611), .CK(CLK), .QN(n21117) );
  DFF_X1 \REGISTERS_reg[29][43]  ( .D(n5610), .CK(CLK), .QN(n21118) );
  DFF_X1 \REGISTERS_reg[29][42]  ( .D(n5609), .CK(CLK), .QN(n21119) );
  DFF_X1 \REGISTERS_reg[29][41]  ( .D(n5608), .CK(CLK), .QN(n21120) );
  DFF_X1 \REGISTERS_reg[29][40]  ( .D(n5607), .CK(CLK), .QN(n21121) );
  DFF_X1 \REGISTERS_reg[29][39]  ( .D(n5606), .CK(CLK), .QN(n21122) );
  DFF_X1 \REGISTERS_reg[29][38]  ( .D(n5605), .CK(CLK), .QN(n21123) );
  DFF_X1 \REGISTERS_reg[29][37]  ( .D(n5604), .CK(CLK), .QN(n21124) );
  DFF_X1 \REGISTERS_reg[29][36]  ( .D(n5603), .CK(CLK), .QN(n21125) );
  DFF_X1 \REGISTERS_reg[29][35]  ( .D(n5602), .CK(CLK), .QN(n21126) );
  DFF_X1 \REGISTERS_reg[29][34]  ( .D(n5601), .CK(CLK), .QN(n21127) );
  DFF_X1 \REGISTERS_reg[29][33]  ( .D(n5600), .CK(CLK), .QN(n21128) );
  DFF_X1 \REGISTERS_reg[29][32]  ( .D(n5599), .CK(CLK), .QN(n21129) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n5598), .CK(CLK), .QN(n21130) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n5597), .CK(CLK), .QN(n21131) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n5596), .CK(CLK), .QN(n21132) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n5595), .CK(CLK), .QN(n21133) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n5594), .CK(CLK), .QN(n21134) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n5593), .CK(CLK), .QN(n21135) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n5592), .CK(CLK), .QN(n21136) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n5591), .CK(CLK), .QN(n21137) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n5590), .CK(CLK), .QN(n21138) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n5589), .CK(CLK), .QN(n21139) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n5588), .CK(CLK), .QN(n21140) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n5587), .CK(CLK), .QN(n21141) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n5586), .CK(CLK), .QN(n21142) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n5585), .CK(CLK), .QN(n21143) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n5584), .CK(CLK), .QN(n21144) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n5583), .CK(CLK), .QN(n21145) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n5582), .CK(CLK), .QN(n21146) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n5581), .CK(CLK), .QN(n21147) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n5580), .CK(CLK), .QN(n21148) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n5579), .CK(CLK), .QN(n21149) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n5578), .CK(CLK), .QN(n21150) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n5577), .CK(CLK), .QN(n21151) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n5576), .CK(CLK), .QN(n21152) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n5575), .CK(CLK), .QN(n21153) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n5574), .CK(CLK), .QN(n21154) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n5573), .CK(CLK), .QN(n21155) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n5572), .CK(CLK), .QN(n21156) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n5571), .CK(CLK), .QN(n21157) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n5570), .CK(CLK), .QN(n21158) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n5569), .CK(CLK), .QN(n21159) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n5568), .CK(CLK), .QN(n21160) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n5567), .CK(CLK), .QN(n21161) );
  DFF_X1 \REGISTERS_reg[26][59]  ( .D(n5818), .CK(CLK), .QN(n21162) );
  DFF_X1 \REGISTERS_reg[26][58]  ( .D(n5817), .CK(CLK), .QN(n21163) );
  DFF_X1 \REGISTERS_reg[26][57]  ( .D(n5816), .CK(CLK), .QN(n21164) );
  DFF_X1 \REGISTERS_reg[26][56]  ( .D(n5815), .CK(CLK), .QN(n21165) );
  DFF_X1 \REGISTERS_reg[26][55]  ( .D(n5814), .CK(CLK), .QN(n21166) );
  DFF_X1 \REGISTERS_reg[26][54]  ( .D(n5813), .CK(CLK), .QN(n21167) );
  DFF_X1 \REGISTERS_reg[26][53]  ( .D(n5812), .CK(CLK), .QN(n21168) );
  DFF_X1 \REGISTERS_reg[26][52]  ( .D(n5811), .CK(CLK), .QN(n21169) );
  DFF_X1 \REGISTERS_reg[26][51]  ( .D(n5810), .CK(CLK), .QN(n21170) );
  DFF_X1 \REGISTERS_reg[26][50]  ( .D(n5809), .CK(CLK), .QN(n21171) );
  DFF_X1 \REGISTERS_reg[26][49]  ( .D(n5808), .CK(CLK), .QN(n21172) );
  DFF_X1 \REGISTERS_reg[26][48]  ( .D(n5807), .CK(CLK), .QN(n21173) );
  DFF_X1 \REGISTERS_reg[26][47]  ( .D(n5806), .CK(CLK), .QN(n21174) );
  DFF_X1 \REGISTERS_reg[26][46]  ( .D(n5805), .CK(CLK), .QN(n21175) );
  DFF_X1 \REGISTERS_reg[26][45]  ( .D(n5804), .CK(CLK), .QN(n21176) );
  DFF_X1 \REGISTERS_reg[26][44]  ( .D(n5803), .CK(CLK), .QN(n21177) );
  DFF_X1 \REGISTERS_reg[26][43]  ( .D(n5802), .CK(CLK), .QN(n21178) );
  DFF_X1 \REGISTERS_reg[26][42]  ( .D(n5801), .CK(CLK), .QN(n21179) );
  DFF_X1 \REGISTERS_reg[26][41]  ( .D(n5800), .CK(CLK), .QN(n21180) );
  DFF_X1 \REGISTERS_reg[26][40]  ( .D(n5799), .CK(CLK), .QN(n21181) );
  DFF_X1 \REGISTERS_reg[26][39]  ( .D(n5798), .CK(CLK), .QN(n21182) );
  DFF_X1 \REGISTERS_reg[26][38]  ( .D(n5797), .CK(CLK), .QN(n21183) );
  DFF_X1 \REGISTERS_reg[26][37]  ( .D(n5796), .CK(CLK), .QN(n21184) );
  DFF_X1 \REGISTERS_reg[26][36]  ( .D(n5795), .CK(CLK), .QN(n21185) );
  DFF_X1 \REGISTERS_reg[26][35]  ( .D(n5794), .CK(CLK), .QN(n21186) );
  DFF_X1 \REGISTERS_reg[26][34]  ( .D(n5793), .CK(CLK), .QN(n21187) );
  DFF_X1 \REGISTERS_reg[26][33]  ( .D(n5792), .CK(CLK), .QN(n21188) );
  DFF_X1 \REGISTERS_reg[26][32]  ( .D(n5791), .CK(CLK), .QN(n21189) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n5790), .CK(CLK), .QN(n21190) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n5789), .CK(CLK), .QN(n21191) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n5788), .CK(CLK), .QN(n21192) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n5787), .CK(CLK), .QN(n21193) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n5786), .CK(CLK), .QN(n21194) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n5785), .CK(CLK), .QN(n21195) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n5784), .CK(CLK), .QN(n21196) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n5783), .CK(CLK), .QN(n21197) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n5782), .CK(CLK), .QN(n21198) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n5781), .CK(CLK), .QN(n21199) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n5780), .CK(CLK), .QN(n21200) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n5779), .CK(CLK), .QN(n21201) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n5778), .CK(CLK), .QN(n21202) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n5777), .CK(CLK), .QN(n21203) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n5776), .CK(CLK), .QN(n21204) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n5775), .CK(CLK), .QN(n21205) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n5774), .CK(CLK), .QN(n21206) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n5773), .CK(CLK), .QN(n21207) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n5772), .CK(CLK), .QN(n21208) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n5771), .CK(CLK), .QN(n21209) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n5770), .CK(CLK), .QN(n21210) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n5769), .CK(CLK), .QN(n21211) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n5768), .CK(CLK), .QN(n21212) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n5767), .CK(CLK), .QN(n21213) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n5766), .CK(CLK), .QN(n21214) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n5765), .CK(CLK), .QN(n21215) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n5764), .CK(CLK), .QN(n21216) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n5763), .CK(CLK), .QN(n21217) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n5762), .CK(CLK), .QN(n21218) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n5761), .CK(CLK), .QN(n21219) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n5760), .CK(CLK), .QN(n21220) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n5759), .CK(CLK), .QN(n21221) );
  DFF_X1 \REGISTERS_reg[11][63]  ( .D(n6782), .CK(CLK), .QN(n21222) );
  DFF_X1 \REGISTERS_reg[11][62]  ( .D(n6781), .CK(CLK), .QN(n21223) );
  DFF_X1 \REGISTERS_reg[11][61]  ( .D(n6780), .CK(CLK), .QN(n21224) );
  DFF_X1 \REGISTERS_reg[11][60]  ( .D(n6779), .CK(CLK), .QN(n21225) );
  DFF_X1 \REGISTERS_reg[11][59]  ( .D(n6778), .CK(CLK), .QN(n21226) );
  DFF_X1 \REGISTERS_reg[11][58]  ( .D(n6777), .CK(CLK), .QN(n21227) );
  DFF_X1 \REGISTERS_reg[11][57]  ( .D(n6776), .CK(CLK), .QN(n21228) );
  DFF_X1 \REGISTERS_reg[11][56]  ( .D(n6775), .CK(CLK), .QN(n21229) );
  DFF_X1 \REGISTERS_reg[11][55]  ( .D(n6774), .CK(CLK), .QN(n21230) );
  DFF_X1 \REGISTERS_reg[11][54]  ( .D(n6773), .CK(CLK), .QN(n21231) );
  DFF_X1 \REGISTERS_reg[11][53]  ( .D(n6772), .CK(CLK), .QN(n21232) );
  DFF_X1 \REGISTERS_reg[11][52]  ( .D(n6771), .CK(CLK), .QN(n21233) );
  DFF_X1 \REGISTERS_reg[11][51]  ( .D(n6770), .CK(CLK), .QN(n21234) );
  DFF_X1 \REGISTERS_reg[11][50]  ( .D(n6769), .CK(CLK), .QN(n21235) );
  DFF_X1 \REGISTERS_reg[11][49]  ( .D(n6768), .CK(CLK), .QN(n21236) );
  DFF_X1 \REGISTERS_reg[11][48]  ( .D(n6767), .CK(CLK), .QN(n21237) );
  DFF_X1 \REGISTERS_reg[11][47]  ( .D(n6766), .CK(CLK), .QN(n21238) );
  DFF_X1 \REGISTERS_reg[11][46]  ( .D(n6765), .CK(CLK), .QN(n21239) );
  DFF_X1 \REGISTERS_reg[11][45]  ( .D(n6764), .CK(CLK), .QN(n21240) );
  DFF_X1 \REGISTERS_reg[11][44]  ( .D(n6763), .CK(CLK), .QN(n21241) );
  DFF_X1 \REGISTERS_reg[11][43]  ( .D(n6762), .CK(CLK), .QN(n21242) );
  DFF_X1 \REGISTERS_reg[11][42]  ( .D(n6761), .CK(CLK), .QN(n21243) );
  DFF_X1 \REGISTERS_reg[11][41]  ( .D(n6760), .CK(CLK), .QN(n21244) );
  DFF_X1 \REGISTERS_reg[11][40]  ( .D(n6759), .CK(CLK), .QN(n21245) );
  DFF_X1 \REGISTERS_reg[11][39]  ( .D(n6758), .CK(CLK), .QN(n21246) );
  DFF_X1 \REGISTERS_reg[11][38]  ( .D(n6757), .CK(CLK), .QN(n21247) );
  DFF_X1 \REGISTERS_reg[11][37]  ( .D(n6756), .CK(CLK), .QN(n21248) );
  DFF_X1 \REGISTERS_reg[11][36]  ( .D(n6755), .CK(CLK), .QN(n21249) );
  DFF_X1 \REGISTERS_reg[11][35]  ( .D(n6754), .CK(CLK), .QN(n21250) );
  DFF_X1 \REGISTERS_reg[11][34]  ( .D(n6753), .CK(CLK), .QN(n21251) );
  DFF_X1 \REGISTERS_reg[11][33]  ( .D(n6752), .CK(CLK), .QN(n21252) );
  DFF_X1 \REGISTERS_reg[11][32]  ( .D(n6751), .CK(CLK), .QN(n21253) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n6750), .CK(CLK), .QN(n21254) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n6749), .CK(CLK), .QN(n21255) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n6748), .CK(CLK), .QN(n21256) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n6747), .CK(CLK), .QN(n21257) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n6746), .CK(CLK), .QN(n21258) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n6745), .CK(CLK), .QN(n21259) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n6744), .CK(CLK), .QN(n21260) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n6743), .CK(CLK), .QN(n21261) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n6742), .CK(CLK), .QN(n21262) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n6741), .CK(CLK), .QN(n21263) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n6740), .CK(CLK), .QN(n21264) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n6739), .CK(CLK), .QN(n21265) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n6738), .CK(CLK), .QN(n21266) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n6737), .CK(CLK), .QN(n21267) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n6736), .CK(CLK), .QN(n21268) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n6735), .CK(CLK), .QN(n21269) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n6734), .CK(CLK), .QN(n21270) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n6733), .CK(CLK), .QN(n21271) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n6732), .CK(CLK), .QN(n21272) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n6731), .CK(CLK), .QN(n21273) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n6730), .CK(CLK), .QN(n21274) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n6729), .CK(CLK), .QN(n21275) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n6728), .CK(CLK), .QN(n21276) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n6727), .CK(CLK), .QN(n21277) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n6726), .CK(CLK), .QN(n21278) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n6725), .CK(CLK), .QN(n21279) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n6724), .CK(CLK), .QN(n21280) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n6723), .CK(CLK), .QN(n21281) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n6722), .CK(CLK), .QN(n21282) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n6721), .CK(CLK), .QN(n21283) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n6720), .CK(CLK), .QN(n21284) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n6719), .CK(CLK), .QN(n21285) );
  DFF_X1 \REGISTERS_reg[9][63]  ( .D(n6910), .CK(CLK), .QN(n20133) );
  DFF_X1 \REGISTERS_reg[9][62]  ( .D(n6909), .CK(CLK), .QN(n19750) );
  DFF_X1 \REGISTERS_reg[9][61]  ( .D(n6908), .CK(CLK), .QN(n19751) );
  DFF_X1 \REGISTERS_reg[9][60]  ( .D(n6907), .CK(CLK), .QN(n19752) );
  DFF_X1 \REGISTERS_reg[9][59]  ( .D(n6906), .CK(CLK), .QN(n19753) );
  DFF_X1 \REGISTERS_reg[9][58]  ( .D(n6905), .CK(CLK), .QN(n19754) );
  DFF_X1 \REGISTERS_reg[9][57]  ( .D(n6904), .CK(CLK), .QN(n19755) );
  DFF_X1 \REGISTERS_reg[9][56]  ( .D(n6903), .CK(CLK), .QN(n19756) );
  DFF_X1 \REGISTERS_reg[9][55]  ( .D(n6902), .CK(CLK), .QN(n19757) );
  DFF_X1 \REGISTERS_reg[9][54]  ( .D(n6901), .CK(CLK), .QN(n19758) );
  DFF_X1 \REGISTERS_reg[9][53]  ( .D(n6900), .CK(CLK), .QN(n19759) );
  DFF_X1 \REGISTERS_reg[9][52]  ( .D(n6899), .CK(CLK), .QN(n19760) );
  DFF_X1 \REGISTERS_reg[9][51]  ( .D(n6898), .CK(CLK), .QN(n19761) );
  DFF_X1 \REGISTERS_reg[9][50]  ( .D(n6897), .CK(CLK), .QN(n19762) );
  DFF_X1 \REGISTERS_reg[9][49]  ( .D(n6896), .CK(CLK), .QN(n19763) );
  DFF_X1 \REGISTERS_reg[9][48]  ( .D(n6895), .CK(CLK), .QN(n19764) );
  DFF_X1 \REGISTERS_reg[9][47]  ( .D(n6894), .CK(CLK), .QN(n19765) );
  DFF_X1 \REGISTERS_reg[9][46]  ( .D(n6893), .CK(CLK), .QN(n19766) );
  DFF_X1 \REGISTERS_reg[9][45]  ( .D(n6892), .CK(CLK), .QN(n19767) );
  DFF_X1 \REGISTERS_reg[9][44]  ( .D(n6891), .CK(CLK), .QN(n19768) );
  DFF_X1 \REGISTERS_reg[9][43]  ( .D(n6890), .CK(CLK), .QN(n19769) );
  DFF_X1 \REGISTERS_reg[9][42]  ( .D(n6889), .CK(CLK), .QN(n19770) );
  DFF_X1 \REGISTERS_reg[9][41]  ( .D(n6888), .CK(CLK), .QN(n19771) );
  DFF_X1 \REGISTERS_reg[9][40]  ( .D(n6887), .CK(CLK), .QN(n19772) );
  DFF_X1 \REGISTERS_reg[9][39]  ( .D(n6886), .CK(CLK), .QN(n19773) );
  DFF_X1 \REGISTERS_reg[9][38]  ( .D(n6885), .CK(CLK), .QN(n19774) );
  DFF_X1 \REGISTERS_reg[9][37]  ( .D(n6884), .CK(CLK), .QN(n19775) );
  DFF_X1 \REGISTERS_reg[9][36]  ( .D(n6883), .CK(CLK), .QN(n19776) );
  DFF_X1 \REGISTERS_reg[9][35]  ( .D(n6882), .CK(CLK), .QN(n19777) );
  DFF_X1 \REGISTERS_reg[9][34]  ( .D(n6881), .CK(CLK), .QN(n19778) );
  DFF_X1 \REGISTERS_reg[9][33]  ( .D(n6880), .CK(CLK), .QN(n19779) );
  DFF_X1 \REGISTERS_reg[9][32]  ( .D(n6879), .CK(CLK), .QN(n19780) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n6878), .CK(CLK), .QN(n19781) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n6877), .CK(CLK), .QN(n19782) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n6876), .CK(CLK), .QN(n19783) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n6875), .CK(CLK), .QN(n19784) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n6874), .CK(CLK), .QN(n19785) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n6873), .CK(CLK), .QN(n19786) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n6872), .CK(CLK), .QN(n19787) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n6871), .CK(CLK), .QN(n19788) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n6870), .CK(CLK), .QN(n19789) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n6869), .CK(CLK), .QN(n19790) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n6868), .CK(CLK), .QN(n19791) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n6867), .CK(CLK), .QN(n19792) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n6866), .CK(CLK), .QN(n19793) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n6865), .CK(CLK), .QN(n19794) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n6864), .CK(CLK), .QN(n19795) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n6863), .CK(CLK), .QN(n19796) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n6862), .CK(CLK), .QN(n19797) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n6861), .CK(CLK), .QN(n19798) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n6860), .CK(CLK), .QN(n19799) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n6859), .CK(CLK), .QN(n19800) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n6858), .CK(CLK), .QN(n19801) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n6857), .CK(CLK), .QN(n19802) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n6856), .CK(CLK), .QN(n19803) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n6855), .CK(CLK), .QN(n19804) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n6854), .CK(CLK), .QN(n19805) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n6853), .CK(CLK), .QN(n19806) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n6852), .CK(CLK), .QN(n19807) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n6851), .CK(CLK), .QN(n19808) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n6850), .CK(CLK), .QN(n19809) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n6849), .CK(CLK), .QN(n19810) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n6848), .CK(CLK), .QN(n19811) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n6847), .CK(CLK), .QN(n19812) );
  DFF_X1 \REGISTERS_reg[4][63]  ( .D(n7230), .CK(CLK), .QN(n20646) );
  DFF_X1 \REGISTERS_reg[4][62]  ( .D(n7229), .CK(CLK), .QN(n20647) );
  DFF_X1 \REGISTERS_reg[4][61]  ( .D(n7228), .CK(CLK), .QN(n20648) );
  DFF_X1 \REGISTERS_reg[4][60]  ( .D(n7227), .CK(CLK), .QN(n20649) );
  DFF_X1 \REGISTERS_reg[4][59]  ( .D(n7226), .CK(CLK), .QN(n20650) );
  DFF_X1 \REGISTERS_reg[4][58]  ( .D(n7225), .CK(CLK), .QN(n20651) );
  DFF_X1 \REGISTERS_reg[4][57]  ( .D(n7224), .CK(CLK), .QN(n20652) );
  DFF_X1 \REGISTERS_reg[4][56]  ( .D(n7223), .CK(CLK), .QN(n20653) );
  DFF_X1 \REGISTERS_reg[4][55]  ( .D(n7222), .CK(CLK), .QN(n20654) );
  DFF_X1 \REGISTERS_reg[4][54]  ( .D(n7221), .CK(CLK), .QN(n20655) );
  DFF_X1 \REGISTERS_reg[4][53]  ( .D(n7220), .CK(CLK), .QN(n20656) );
  DFF_X1 \REGISTERS_reg[4][52]  ( .D(n7219), .CK(CLK), .QN(n20657) );
  DFF_X1 \REGISTERS_reg[4][51]  ( .D(n7218), .CK(CLK), .QN(n20658) );
  DFF_X1 \REGISTERS_reg[4][50]  ( .D(n7217), .CK(CLK), .QN(n20659) );
  DFF_X1 \REGISTERS_reg[4][49]  ( .D(n7216), .CK(CLK), .QN(n20660) );
  DFF_X1 \REGISTERS_reg[4][48]  ( .D(n7215), .CK(CLK), .QN(n20661) );
  DFF_X1 \REGISTERS_reg[4][47]  ( .D(n7214), .CK(CLK), .QN(n20662) );
  DFF_X1 \REGISTERS_reg[4][46]  ( .D(n7213), .CK(CLK), .QN(n20663) );
  DFF_X1 \REGISTERS_reg[4][45]  ( .D(n7212), .CK(CLK), .QN(n20664) );
  DFF_X1 \REGISTERS_reg[4][44]  ( .D(n7211), .CK(CLK), .QN(n20665) );
  DFF_X1 \REGISTERS_reg[4][43]  ( .D(n7210), .CK(CLK), .QN(n20666) );
  DFF_X1 \REGISTERS_reg[4][42]  ( .D(n7209), .CK(CLK), .QN(n20667) );
  DFF_X1 \REGISTERS_reg[4][41]  ( .D(n7208), .CK(CLK), .QN(n20668) );
  DFF_X1 \REGISTERS_reg[4][40]  ( .D(n7207), .CK(CLK), .QN(n20669) );
  DFF_X1 \REGISTERS_reg[4][39]  ( .D(n7206), .CK(CLK), .QN(n20670) );
  DFF_X1 \REGISTERS_reg[4][38]  ( .D(n7205), .CK(CLK), .QN(n20671) );
  DFF_X1 \REGISTERS_reg[4][37]  ( .D(n7204), .CK(CLK), .QN(n20672) );
  DFF_X1 \REGISTERS_reg[4][36]  ( .D(n7203), .CK(CLK), .QN(n20673) );
  DFF_X1 \REGISTERS_reg[4][35]  ( .D(n7202), .CK(CLK), .QN(n20674) );
  DFF_X1 \REGISTERS_reg[4][34]  ( .D(n7201), .CK(CLK), .QN(n20675) );
  DFF_X1 \REGISTERS_reg[4][33]  ( .D(n7200), .CK(CLK), .QN(n20676) );
  DFF_X1 \REGISTERS_reg[4][32]  ( .D(n7199), .CK(CLK), .QN(n20677) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n7198), .CK(CLK), .QN(n20678) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n7197), .CK(CLK), .QN(n20679) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n7196), .CK(CLK), .QN(n20680) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n7195), .CK(CLK), .QN(n20681) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n7194), .CK(CLK), .QN(n20682) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n7193), .CK(CLK), .QN(n20683) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n7192), .CK(CLK), .QN(n20684) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n7191), .CK(CLK), .QN(n20685) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n7190), .CK(CLK), .QN(n20686) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n7189), .CK(CLK), .QN(n20687) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n7188), .CK(CLK), .QN(n20688) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n7187), .CK(CLK), .QN(n20689) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n7186), .CK(CLK), .QN(n20690) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n7185), .CK(CLK), .QN(n20691) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n7184), .CK(CLK), .QN(n20692) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n7183), .CK(CLK), .QN(n20693) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n7182), .CK(CLK), .QN(n20694) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n7181), .CK(CLK), .QN(n20695) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n7180), .CK(CLK), .QN(n20696) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n7179), .CK(CLK), .QN(n20697) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n7178), .CK(CLK), .QN(n20698) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n7177), .CK(CLK), .QN(n20699) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n7176), .CK(CLK), .QN(n20700) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n7175), .CK(CLK), .QN(n20701) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n7174), .CK(CLK), .QN(n20702) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n7173), .CK(CLK), .QN(n20703) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n7172), .CK(CLK), .QN(n20704) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n7171), .CK(CLK), .QN(n20705) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n7170), .CK(CLK), .QN(n20706) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n7169), .CK(CLK), .QN(n20707) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n7168), .CK(CLK), .QN(n20708) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n7167), .CK(CLK), .QN(n20709) );
  DFF_X1 \REGISTERS_reg[19][63]  ( .D(n6270), .CK(CLK), .QN(n20710) );
  DFF_X1 \REGISTERS_reg[19][62]  ( .D(n6269), .CK(CLK), .QN(n20711) );
  DFF_X1 \REGISTERS_reg[19][61]  ( .D(n6268), .CK(CLK), .QN(n20712) );
  DFF_X1 \REGISTERS_reg[19][60]  ( .D(n6267), .CK(CLK), .QN(n20713) );
  DFF_X1 \REGISTERS_reg[19][59]  ( .D(n6266), .CK(CLK), .QN(n20714) );
  DFF_X1 \REGISTERS_reg[19][58]  ( .D(n6265), .CK(CLK), .QN(n20715) );
  DFF_X1 \REGISTERS_reg[19][57]  ( .D(n6264), .CK(CLK), .QN(n20716) );
  DFF_X1 \REGISTERS_reg[19][56]  ( .D(n6263), .CK(CLK), .QN(n20717) );
  DFF_X1 \REGISTERS_reg[19][55]  ( .D(n6262), .CK(CLK), .QN(n20718) );
  DFF_X1 \REGISTERS_reg[19][54]  ( .D(n6261), .CK(CLK), .QN(n20719) );
  DFF_X1 \REGISTERS_reg[19][53]  ( .D(n6260), .CK(CLK), .QN(n20720) );
  DFF_X1 \REGISTERS_reg[19][52]  ( .D(n6259), .CK(CLK), .QN(n20721) );
  DFF_X1 \REGISTERS_reg[19][51]  ( .D(n6258), .CK(CLK), .QN(n20722) );
  DFF_X1 \REGISTERS_reg[19][50]  ( .D(n6257), .CK(CLK), .QN(n20723) );
  DFF_X1 \REGISTERS_reg[19][49]  ( .D(n6256), .CK(CLK), .QN(n20724) );
  DFF_X1 \REGISTERS_reg[19][48]  ( .D(n6255), .CK(CLK), .QN(n20725) );
  DFF_X1 \REGISTERS_reg[19][47]  ( .D(n6254), .CK(CLK), .QN(n20726) );
  DFF_X1 \REGISTERS_reg[19][46]  ( .D(n6253), .CK(CLK), .QN(n20727) );
  DFF_X1 \REGISTERS_reg[19][45]  ( .D(n6252), .CK(CLK), .QN(n20728) );
  DFF_X1 \REGISTERS_reg[19][44]  ( .D(n6251), .CK(CLK), .QN(n20729) );
  DFF_X1 \REGISTERS_reg[19][43]  ( .D(n6250), .CK(CLK), .QN(n20730) );
  DFF_X1 \REGISTERS_reg[19][42]  ( .D(n6249), .CK(CLK), .QN(n20731) );
  DFF_X1 \REGISTERS_reg[19][41]  ( .D(n6248), .CK(CLK), .QN(n20732) );
  DFF_X1 \REGISTERS_reg[19][40]  ( .D(n6247), .CK(CLK), .QN(n20733) );
  DFF_X1 \REGISTERS_reg[19][39]  ( .D(n6246), .CK(CLK), .QN(n20734) );
  DFF_X1 \REGISTERS_reg[19][38]  ( .D(n6245), .CK(CLK), .QN(n20735) );
  DFF_X1 \REGISTERS_reg[19][37]  ( .D(n6244), .CK(CLK), .QN(n20736) );
  DFF_X1 \REGISTERS_reg[19][36]  ( .D(n6243), .CK(CLK), .QN(n20737) );
  DFF_X1 \REGISTERS_reg[19][35]  ( .D(n6242), .CK(CLK), .QN(n20738) );
  DFF_X1 \REGISTERS_reg[19][34]  ( .D(n6241), .CK(CLK), .QN(n20739) );
  DFF_X1 \REGISTERS_reg[19][33]  ( .D(n6240), .CK(CLK), .QN(n20740) );
  DFF_X1 \REGISTERS_reg[19][32]  ( .D(n6239), .CK(CLK), .QN(n20741) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n6238), .CK(CLK), .QN(n20742) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n6237), .CK(CLK), .QN(n20743) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n6236), .CK(CLK), .QN(n20744) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n6235), .CK(CLK), .QN(n20745) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n6234), .CK(CLK), .QN(n20746) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n6233), .CK(CLK), .QN(n20747) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n6232), .CK(CLK), .QN(n20748) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n6231), .CK(CLK), .QN(n20749) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n6230), .CK(CLK), .QN(n20750) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n6229), .CK(CLK), .QN(n20751) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n6228), .CK(CLK), .QN(n20752) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n6227), .CK(CLK), .QN(n20753) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n6226), .CK(CLK), .QN(n20754) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n6225), .CK(CLK), .QN(n20755) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n6224), .CK(CLK), .QN(n20756) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n6223), .CK(CLK), .QN(n20757) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n6222), .CK(CLK), .QN(n20758) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n6221), .CK(CLK), .QN(n20759) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n6220), .CK(CLK), .QN(n20760) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n6219), .CK(CLK), .QN(n20761) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n6218), .CK(CLK), .QN(n20762) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n6217), .CK(CLK), .QN(n20763) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n6216), .CK(CLK), .QN(n20764) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n6215), .CK(CLK), .QN(n20765) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n6214), .CK(CLK), .QN(n20766) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n6213), .CK(CLK), .QN(n20767) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n6212), .CK(CLK), .QN(n20768) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n6211), .CK(CLK), .QN(n20769) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n6210), .CK(CLK), .QN(n20770) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n6209), .CK(CLK), .QN(n20771) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n6208), .CK(CLK), .QN(n20772) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n6207), .CK(CLK), .QN(n20773) );
  DFF_X1 \REGISTERS_reg[17][63]  ( .D(n6398), .CK(CLK), .QN(n21350) );
  DFF_X1 \REGISTERS_reg[17][62]  ( .D(n6397), .CK(CLK), .QN(n21351) );
  DFF_X1 \REGISTERS_reg[17][61]  ( .D(n6396), .CK(CLK), .QN(n21352) );
  DFF_X1 \REGISTERS_reg[17][60]  ( .D(n6395), .CK(CLK), .QN(n21353) );
  DFF_X1 \REGISTERS_reg[17][59]  ( .D(n6394), .CK(CLK), .QN(n21354) );
  DFF_X1 \REGISTERS_reg[17][58]  ( .D(n6393), .CK(CLK), .QN(n21355) );
  DFF_X1 \REGISTERS_reg[17][57]  ( .D(n6392), .CK(CLK), .QN(n21356) );
  DFF_X1 \REGISTERS_reg[17][56]  ( .D(n6391), .CK(CLK), .QN(n21357) );
  DFF_X1 \REGISTERS_reg[17][55]  ( .D(n6390), .CK(CLK), .QN(n21358) );
  DFF_X1 \REGISTERS_reg[17][54]  ( .D(n6389), .CK(CLK), .QN(n21359) );
  DFF_X1 \REGISTERS_reg[17][53]  ( .D(n6388), .CK(CLK), .QN(n21360) );
  DFF_X1 \REGISTERS_reg[17][52]  ( .D(n6387), .CK(CLK), .QN(n21361) );
  DFF_X1 \REGISTERS_reg[17][51]  ( .D(n6386), .CK(CLK), .QN(n21362) );
  DFF_X1 \REGISTERS_reg[17][50]  ( .D(n6385), .CK(CLK), .QN(n21363) );
  DFF_X1 \REGISTERS_reg[17][49]  ( .D(n6384), .CK(CLK), .QN(n21364) );
  DFF_X1 \REGISTERS_reg[17][48]  ( .D(n6383), .CK(CLK), .QN(n21365) );
  DFF_X1 \REGISTERS_reg[17][47]  ( .D(n6382), .CK(CLK), .QN(n21366) );
  DFF_X1 \REGISTERS_reg[17][46]  ( .D(n6381), .CK(CLK), .QN(n21367) );
  DFF_X1 \REGISTERS_reg[17][45]  ( .D(n6380), .CK(CLK), .QN(n21368) );
  DFF_X1 \REGISTERS_reg[17][44]  ( .D(n6379), .CK(CLK), .QN(n21369) );
  DFF_X1 \REGISTERS_reg[17][43]  ( .D(n6378), .CK(CLK), .QN(n21370) );
  DFF_X1 \REGISTERS_reg[17][42]  ( .D(n6377), .CK(CLK), .QN(n21371) );
  DFF_X1 \REGISTERS_reg[17][41]  ( .D(n6376), .CK(CLK), .QN(n21372) );
  DFF_X1 \REGISTERS_reg[17][40]  ( .D(n6375), .CK(CLK), .QN(n21373) );
  DFF_X1 \REGISTERS_reg[17][39]  ( .D(n6374), .CK(CLK), .QN(n21374) );
  DFF_X1 \REGISTERS_reg[17][38]  ( .D(n6373), .CK(CLK), .QN(n21375) );
  DFF_X1 \REGISTERS_reg[17][37]  ( .D(n6372), .CK(CLK), .QN(n21376) );
  DFF_X1 \REGISTERS_reg[17][36]  ( .D(n6371), .CK(CLK), .QN(n21377) );
  DFF_X1 \REGISTERS_reg[17][35]  ( .D(n6370), .CK(CLK), .QN(n21378) );
  DFF_X1 \REGISTERS_reg[17][34]  ( .D(n6369), .CK(CLK), .QN(n21379) );
  DFF_X1 \REGISTERS_reg[17][33]  ( .D(n6368), .CK(CLK), .QN(n21380) );
  DFF_X1 \REGISTERS_reg[17][32]  ( .D(n6367), .CK(CLK), .QN(n21381) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n6366), .CK(CLK), .QN(n21382) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n6365), .CK(CLK), .QN(n21383) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n6364), .CK(CLK), .QN(n21384) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n6363), .CK(CLK), .QN(n21385) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n6362), .CK(CLK), .QN(n21386) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n6361), .CK(CLK), .QN(n21387) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n6360), .CK(CLK), .QN(n21388) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n6359), .CK(CLK), .QN(n21389) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n6358), .CK(CLK), .QN(n21390) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n6357), .CK(CLK), .QN(n21391) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n6356), .CK(CLK), .QN(n21392) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n6355), .CK(CLK), .QN(n21393) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n6354), .CK(CLK), .QN(n21394) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n6353), .CK(CLK), .QN(n21395) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n6352), .CK(CLK), .QN(n21396) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n6351), .CK(CLK), .QN(n21397) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n6350), .CK(CLK), .QN(n21398) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n6349), .CK(CLK), .QN(n21399) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n6348), .CK(CLK), .QN(n21400) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n6347), .CK(CLK), .QN(n21401) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n6346), .CK(CLK), .QN(n21402) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n6345), .CK(CLK), .QN(n21403) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n6344), .CK(CLK), .QN(n21404) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n6343), .CK(CLK), .QN(n21405) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n6342), .CK(CLK), .QN(n21406) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n6341), .CK(CLK), .QN(n21407) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n6340), .CK(CLK), .QN(n21408) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n6339), .CK(CLK), .QN(n21409) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n6338), .CK(CLK), .QN(n21410) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n6337), .CK(CLK), .QN(n21411) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n6336), .CK(CLK), .QN(n21412) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n6335), .CK(CLK), .QN(n21413) );
  DFF_X1 \REGISTERS_reg[31][63]  ( .D(n5502), .CK(CLK), .Q(n17163), .QN(n20774) );
  DFF_X1 \REGISTERS_reg[31][62]  ( .D(n5501), .CK(CLK), .Q(n17184), .QN(n20775) );
  DFF_X1 \REGISTERS_reg[31][61]  ( .D(n5500), .CK(CLK), .Q(n17205), .QN(n20776) );
  DFF_X1 \REGISTERS_reg[31][60]  ( .D(n5499), .CK(CLK), .Q(n17226), .QN(n20777) );
  DFF_X1 \REGISTERS_reg[25][63]  ( .D(n5886), .CK(CLK), .Q(n17161), .QN(n20778) );
  DFF_X1 \REGISTERS_reg[25][62]  ( .D(n5885), .CK(CLK), .Q(n17182), .QN(n20779) );
  DFF_X1 \REGISTERS_reg[25][61]  ( .D(n5884), .CK(CLK), .Q(n17203), .QN(n20780) );
  DFF_X1 \REGISTERS_reg[25][60]  ( .D(n5883), .CK(CLK), .Q(n17224), .QN(n20781) );
  DFF_X1 \REGISTERS_reg[31][59]  ( .D(n5498), .CK(CLK), .Q(n17247), .QN(n20782) );
  DFF_X1 \REGISTERS_reg[31][58]  ( .D(n5497), .CK(CLK), .Q(n17268), .QN(n20783) );
  DFF_X1 \REGISTERS_reg[31][57]  ( .D(n5496), .CK(CLK), .Q(n17289), .QN(n20784) );
  DFF_X1 \REGISTERS_reg[31][56]  ( .D(n5495), .CK(CLK), .Q(n17310), .QN(n20785) );
  DFF_X1 \REGISTERS_reg[31][55]  ( .D(n5494), .CK(CLK), .Q(n17331), .QN(n20786) );
  DFF_X1 \REGISTERS_reg[31][54]  ( .D(n5493), .CK(CLK), .Q(n17352), .QN(n20787) );
  DFF_X1 \REGISTERS_reg[31][53]  ( .D(n5492), .CK(CLK), .Q(n17373), .QN(n20788) );
  DFF_X1 \REGISTERS_reg[31][52]  ( .D(n5491), .CK(CLK), .Q(n17394), .QN(n20789) );
  DFF_X1 \REGISTERS_reg[31][51]  ( .D(n5490), .CK(CLK), .Q(n17415), .QN(n20790) );
  DFF_X1 \REGISTERS_reg[31][50]  ( .D(n5489), .CK(CLK), .Q(n17436), .QN(n20791) );
  DFF_X1 \REGISTERS_reg[31][49]  ( .D(n5488), .CK(CLK), .Q(n17457), .QN(n20792) );
  DFF_X1 \REGISTERS_reg[31][48]  ( .D(n5487), .CK(CLK), .Q(n17478), .QN(n20793) );
  DFF_X1 \REGISTERS_reg[31][47]  ( .D(n5486), .CK(CLK), .Q(n17499), .QN(n20794) );
  DFF_X1 \REGISTERS_reg[31][46]  ( .D(n5485), .CK(CLK), .Q(n17520), .QN(n20795) );
  DFF_X1 \REGISTERS_reg[31][45]  ( .D(n5484), .CK(CLK), .Q(n17541), .QN(n20796) );
  DFF_X1 \REGISTERS_reg[31][44]  ( .D(n5483), .CK(CLK), .Q(n17562), .QN(n20797) );
  DFF_X1 \REGISTERS_reg[31][43]  ( .D(n5482), .CK(CLK), .Q(n17583), .QN(n20798) );
  DFF_X1 \REGISTERS_reg[31][42]  ( .D(n5481), .CK(CLK), .Q(n17604), .QN(n20799) );
  DFF_X1 \REGISTERS_reg[31][41]  ( .D(n5480), .CK(CLK), .Q(n17625), .QN(n20800) );
  DFF_X1 \REGISTERS_reg[31][40]  ( .D(n5479), .CK(CLK), .Q(n17646), .QN(n20801) );
  DFF_X1 \REGISTERS_reg[31][39]  ( .D(n5478), .CK(CLK), .Q(n17667), .QN(n20802) );
  DFF_X1 \REGISTERS_reg[31][38]  ( .D(n5477), .CK(CLK), .Q(n17688), .QN(n20803) );
  DFF_X1 \REGISTERS_reg[31][37]  ( .D(n5476), .CK(CLK), .Q(n17709), .QN(n20804) );
  DFF_X1 \REGISTERS_reg[31][36]  ( .D(n5475), .CK(CLK), .Q(n17730), .QN(n20805) );
  DFF_X1 \REGISTERS_reg[31][35]  ( .D(n5474), .CK(CLK), .Q(n17751), .QN(n20806) );
  DFF_X1 \REGISTERS_reg[31][34]  ( .D(n5473), .CK(CLK), .Q(n17772), .QN(n20807) );
  DFF_X1 \REGISTERS_reg[31][33]  ( .D(n5472), .CK(CLK), .Q(n17793), .QN(n20808) );
  DFF_X1 \REGISTERS_reg[31][32]  ( .D(n5471), .CK(CLK), .Q(n17814), .QN(n20809) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n5470), .CK(CLK), .Q(n17835), .QN(n20810) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n5469), .CK(CLK), .Q(n17856), .QN(n20811) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n5468), .CK(CLK), .Q(n17877), .QN(n20812) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n5467), .CK(CLK), .Q(n17898), .QN(n20813) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n5466), .CK(CLK), .Q(n17919), .QN(n20814) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n5465), .CK(CLK), .Q(n17940), .QN(n20815) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n5464), .CK(CLK), .Q(n17961), .QN(n20816) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n5463), .CK(CLK), .Q(n17982), .QN(n20817) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n5462), .CK(CLK), .Q(n18003), .QN(n20818) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n5461), .CK(CLK), .Q(n18024), .QN(n20819) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n5460), .CK(CLK), .Q(n18045), .QN(n20820) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n5459), .CK(CLK), .Q(n18066), .QN(n20821) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n5458), .CK(CLK), .Q(n18087), .QN(n20822) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n5457), .CK(CLK), .Q(n18108), .QN(n20823) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n5456), .CK(CLK), .Q(n18129), .QN(n20824) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n5455), .CK(CLK), .Q(n18150), .QN(n20825) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n5454), .CK(CLK), .Q(n18171), .QN(n20826) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n5453), .CK(CLK), .Q(n18192), .QN(n20827) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n5452), .CK(CLK), .Q(n18213), .QN(n20828) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n5451), .CK(CLK), .Q(n18234), .QN(n20829) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n5450), .CK(CLK), .Q(n18255), .QN(n20830) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n5449), .CK(CLK), .Q(n18276), .QN(n20831) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n5448), .CK(CLK), .Q(n18297), .QN(n20832)
         );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n5447), .CK(CLK), .Q(n18318), .QN(n20833)
         );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n5446), .CK(CLK), .Q(n18339), .QN(n20834)
         );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n5445), .CK(CLK), .Q(n18360), .QN(n20835)
         );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n5444), .CK(CLK), .Q(n18381), .QN(n20836)
         );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n5443), .CK(CLK), .Q(n18402), .QN(n20837)
         );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n5442), .CK(CLK), .Q(n18423), .QN(n20838)
         );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n5441), .CK(CLK), .Q(n18444), .QN(n20839)
         );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n5440), .CK(CLK), .Q(n18465), .QN(n20840)
         );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n5439), .CK(CLK), .Q(n18486), .QN(n20841)
         );
  DFF_X1 \REGISTERS_reg[25][59]  ( .D(n5882), .CK(CLK), .Q(n17245), .QN(n20842) );
  DFF_X1 \REGISTERS_reg[25][58]  ( .D(n5881), .CK(CLK), .Q(n17266), .QN(n20843) );
  DFF_X1 \REGISTERS_reg[25][57]  ( .D(n5880), .CK(CLK), .Q(n17287), .QN(n20844) );
  DFF_X1 \REGISTERS_reg[25][56]  ( .D(n5879), .CK(CLK), .Q(n17308), .QN(n20845) );
  DFF_X1 \REGISTERS_reg[25][55]  ( .D(n5878), .CK(CLK), .Q(n17329), .QN(n20846) );
  DFF_X1 \REGISTERS_reg[25][54]  ( .D(n5877), .CK(CLK), .Q(n17350), .QN(n20847) );
  DFF_X1 \REGISTERS_reg[25][53]  ( .D(n5876), .CK(CLK), .Q(n17371), .QN(n20848) );
  DFF_X1 \REGISTERS_reg[25][52]  ( .D(n5875), .CK(CLK), .Q(n17392), .QN(n20849) );
  DFF_X1 \REGISTERS_reg[25][51]  ( .D(n5874), .CK(CLK), .Q(n17413), .QN(n20850) );
  DFF_X1 \REGISTERS_reg[25][50]  ( .D(n5873), .CK(CLK), .Q(n17434), .QN(n20851) );
  DFF_X1 \REGISTERS_reg[25][49]  ( .D(n5872), .CK(CLK), .Q(n17455), .QN(n20852) );
  DFF_X1 \REGISTERS_reg[25][48]  ( .D(n5871), .CK(CLK), .Q(n17476), .QN(n20853) );
  DFF_X1 \REGISTERS_reg[25][47]  ( .D(n5870), .CK(CLK), .Q(n17497), .QN(n20854) );
  DFF_X1 \REGISTERS_reg[25][46]  ( .D(n5869), .CK(CLK), .Q(n17518), .QN(n20855) );
  DFF_X1 \REGISTERS_reg[25][45]  ( .D(n5868), .CK(CLK), .Q(n17539), .QN(n20856) );
  DFF_X1 \REGISTERS_reg[25][44]  ( .D(n5867), .CK(CLK), .Q(n17560), .QN(n20857) );
  DFF_X1 \REGISTERS_reg[25][43]  ( .D(n5866), .CK(CLK), .Q(n17581), .QN(n20858) );
  DFF_X1 \REGISTERS_reg[25][42]  ( .D(n5865), .CK(CLK), .Q(n17602), .QN(n20859) );
  DFF_X1 \REGISTERS_reg[25][41]  ( .D(n5864), .CK(CLK), .Q(n17623), .QN(n20860) );
  DFF_X1 \REGISTERS_reg[25][40]  ( .D(n5863), .CK(CLK), .Q(n17644), .QN(n20861) );
  DFF_X1 \REGISTERS_reg[25][39]  ( .D(n5862), .CK(CLK), .Q(n17665), .QN(n20862) );
  DFF_X1 \REGISTERS_reg[25][38]  ( .D(n5861), .CK(CLK), .Q(n17686), .QN(n20863) );
  DFF_X1 \REGISTERS_reg[25][37]  ( .D(n5860), .CK(CLK), .Q(n17707), .QN(n20864) );
  DFF_X1 \REGISTERS_reg[25][36]  ( .D(n5859), .CK(CLK), .Q(n17728), .QN(n20865) );
  DFF_X1 \REGISTERS_reg[25][35]  ( .D(n5858), .CK(CLK), .Q(n17749), .QN(n20866) );
  DFF_X1 \REGISTERS_reg[25][34]  ( .D(n5857), .CK(CLK), .Q(n17770), .QN(n20867) );
  DFF_X1 \REGISTERS_reg[25][33]  ( .D(n5856), .CK(CLK), .Q(n17791), .QN(n20868) );
  DFF_X1 \REGISTERS_reg[25][32]  ( .D(n5855), .CK(CLK), .Q(n17812), .QN(n20869) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n5854), .CK(CLK), .Q(n17833), .QN(n20870) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n5853), .CK(CLK), .Q(n17854), .QN(n20871) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n5852), .CK(CLK), .Q(n17875), .QN(n20872) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n5851), .CK(CLK), .Q(n17896), .QN(n20873) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n5850), .CK(CLK), .Q(n17917), .QN(n20874) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n5849), .CK(CLK), .Q(n17938), .QN(n20875) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n5848), .CK(CLK), .Q(n17959), .QN(n20876) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n5847), .CK(CLK), .Q(n17980), .QN(n20877) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n5846), .CK(CLK), .Q(n18001), .QN(n20878) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n5845), .CK(CLK), .Q(n18022), .QN(n20879) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n5844), .CK(CLK), .Q(n18043), .QN(n20880) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n5843), .CK(CLK), .Q(n18064), .QN(n20881) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n5842), .CK(CLK), .Q(n18085), .QN(n20882) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n5841), .CK(CLK), .Q(n18106), .QN(n20883) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n5840), .CK(CLK), .Q(n18127), .QN(n20884) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n5839), .CK(CLK), .Q(n18148), .QN(n20885) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n5838), .CK(CLK), .Q(n18169), .QN(n20886) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n5837), .CK(CLK), .Q(n18190), .QN(n20887) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n5836), .CK(CLK), .Q(n18211), .QN(n20888) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n5835), .CK(CLK), .Q(n18232), .QN(n20889) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n5834), .CK(CLK), .Q(n18253), .QN(n20890) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n5833), .CK(CLK), .Q(n18274), .QN(n20891) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n5832), .CK(CLK), .Q(n18295), .QN(n20892)
         );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n5831), .CK(CLK), .Q(n18316), .QN(n20893)
         );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n5830), .CK(CLK), .Q(n18337), .QN(n20894)
         );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n5829), .CK(CLK), .Q(n18358), .QN(n20895)
         );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n5828), .CK(CLK), .Q(n18379), .QN(n20896)
         );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n5827), .CK(CLK), .Q(n18400), .QN(n20897)
         );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n5826), .CK(CLK), .Q(n18421), .QN(n20898)
         );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n5825), .CK(CLK), .Q(n18442), .QN(n20899)
         );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n5824), .CK(CLK), .Q(n18463), .QN(n20900)
         );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n5823), .CK(CLK), .Q(n18484), .QN(n20901)
         );
  DFF_X1 \REGISTERS_reg[24][63]  ( .D(n5950), .CK(CLK), .Q(n17156), .QN(n21286) );
  DFF_X1 \REGISTERS_reg[24][62]  ( .D(n5949), .CK(CLK), .Q(n17177), .QN(n21287) );
  DFF_X1 \REGISTERS_reg[24][61]  ( .D(n5948), .CK(CLK), .Q(n17198), .QN(n21288) );
  DFF_X1 \REGISTERS_reg[24][60]  ( .D(n5947), .CK(CLK), .Q(n17219), .QN(n21289) );
  DFF_X1 \REGISTERS_reg[24][59]  ( .D(n5946), .CK(CLK), .Q(n17240), .QN(n21290) );
  DFF_X1 \REGISTERS_reg[24][58]  ( .D(n5945), .CK(CLK), .Q(n17261), .QN(n21291) );
  DFF_X1 \REGISTERS_reg[24][57]  ( .D(n5944), .CK(CLK), .Q(n17282), .QN(n21292) );
  DFF_X1 \REGISTERS_reg[24][56]  ( .D(n5943), .CK(CLK), .Q(n17303), .QN(n21293) );
  DFF_X1 \REGISTERS_reg[24][55]  ( .D(n5942), .CK(CLK), .Q(n17324), .QN(n21294) );
  DFF_X1 \REGISTERS_reg[24][54]  ( .D(n5941), .CK(CLK), .Q(n17345), .QN(n21295) );
  DFF_X1 \REGISTERS_reg[24][53]  ( .D(n5940), .CK(CLK), .Q(n17366), .QN(n21296) );
  DFF_X1 \REGISTERS_reg[24][52]  ( .D(n5939), .CK(CLK), .Q(n17387), .QN(n21297) );
  DFF_X1 \REGISTERS_reg[24][51]  ( .D(n5938), .CK(CLK), .Q(n17408), .QN(n21298) );
  DFF_X1 \REGISTERS_reg[24][50]  ( .D(n5937), .CK(CLK), .Q(n17429), .QN(n21299) );
  DFF_X1 \REGISTERS_reg[24][49]  ( .D(n5936), .CK(CLK), .Q(n17450), .QN(n21300) );
  DFF_X1 \REGISTERS_reg[24][48]  ( .D(n5935), .CK(CLK), .Q(n17471), .QN(n21301) );
  DFF_X1 \REGISTERS_reg[24][47]  ( .D(n5934), .CK(CLK), .Q(n17492), .QN(n21302) );
  DFF_X1 \REGISTERS_reg[24][46]  ( .D(n5933), .CK(CLK), .Q(n17513), .QN(n21303) );
  DFF_X1 \REGISTERS_reg[24][45]  ( .D(n5932), .CK(CLK), .Q(n17534), .QN(n21304) );
  DFF_X1 \REGISTERS_reg[24][44]  ( .D(n5931), .CK(CLK), .Q(n17555), .QN(n21305) );
  DFF_X1 \REGISTERS_reg[24][43]  ( .D(n5930), .CK(CLK), .Q(n17576), .QN(n21306) );
  DFF_X1 \REGISTERS_reg[24][42]  ( .D(n5929), .CK(CLK), .Q(n17597), .QN(n21307) );
  DFF_X1 \REGISTERS_reg[24][41]  ( .D(n5928), .CK(CLK), .Q(n17618), .QN(n21308) );
  DFF_X1 \REGISTERS_reg[24][40]  ( .D(n5927), .CK(CLK), .Q(n17639), .QN(n21309) );
  DFF_X1 \REGISTERS_reg[24][39]  ( .D(n5926), .CK(CLK), .Q(n17660), .QN(n21310) );
  DFF_X1 \REGISTERS_reg[24][38]  ( .D(n5925), .CK(CLK), .Q(n17681), .QN(n21311) );
  DFF_X1 \REGISTERS_reg[24][37]  ( .D(n5924), .CK(CLK), .Q(n17702), .QN(n21312) );
  DFF_X1 \REGISTERS_reg[24][36]  ( .D(n5923), .CK(CLK), .Q(n17723), .QN(n21313) );
  DFF_X1 \REGISTERS_reg[24][35]  ( .D(n5922), .CK(CLK), .Q(n17744), .QN(n21314) );
  DFF_X1 \REGISTERS_reg[24][34]  ( .D(n5921), .CK(CLK), .Q(n17765), .QN(n21315) );
  DFF_X1 \REGISTERS_reg[24][33]  ( .D(n5920), .CK(CLK), .Q(n17786), .QN(n21316) );
  DFF_X1 \REGISTERS_reg[24][32]  ( .D(n5919), .CK(CLK), .Q(n17807), .QN(n21317) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n5918), .CK(CLK), .Q(n17828), .QN(n21318) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n5917), .CK(CLK), .Q(n17849), .QN(n21319) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n5916), .CK(CLK), .Q(n17870), .QN(n21320) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n5915), .CK(CLK), .Q(n17891), .QN(n21321) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n5914), .CK(CLK), .Q(n17912), .QN(n21322) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n5913), .CK(CLK), .Q(n17933), .QN(n21323) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n5912), .CK(CLK), .Q(n17954), .QN(n21324) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n5911), .CK(CLK), .Q(n17975), .QN(n21325) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n5910), .CK(CLK), .Q(n17996), .QN(n21326) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n5909), .CK(CLK), .Q(n18017), .QN(n21327) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n5908), .CK(CLK), .Q(n18038), .QN(n21328) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n5907), .CK(CLK), .Q(n18059), .QN(n21329) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n5906), .CK(CLK), .Q(n18080), .QN(n21330) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n5905), .CK(CLK), .Q(n18101), .QN(n21331) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n5904), .CK(CLK), .Q(n18122), .QN(n21332) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n5903), .CK(CLK), .Q(n18143), .QN(n21333) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n5902), .CK(CLK), .Q(n18164), .QN(n21334) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n5901), .CK(CLK), .Q(n18185), .QN(n21335) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n5900), .CK(CLK), .Q(n18206), .QN(n21336) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n5899), .CK(CLK), .Q(n18227), .QN(n21337) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n5898), .CK(CLK), .Q(n18248), .QN(n21338) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n5897), .CK(CLK), .Q(n18269), .QN(n21339) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n5896), .CK(CLK), .Q(n18290), .QN(n21340)
         );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n5895), .CK(CLK), .Q(n18311), .QN(n21341)
         );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n5894), .CK(CLK), .Q(n18332), .QN(n21342)
         );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n5893), .CK(CLK), .Q(n18353), .QN(n21343)
         );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n5892), .CK(CLK), .Q(n18374), .QN(n21344)
         );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n5891), .CK(CLK), .Q(n18395), .QN(n21345)
         );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n5890), .CK(CLK), .Q(n18416), .QN(n21346)
         );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n5889), .CK(CLK), .Q(n18437), .QN(n21347)
         );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n5888), .CK(CLK), .Q(n18458), .QN(n21348)
         );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n5887), .CK(CLK), .Q(n18479), .QN(n21349)
         );
  DFF_X1 \REGISTERS_reg[8][63]  ( .D(n6974), .CK(CLK), .Q(n24477), .QN(n19686)
         );
  DFF_X1 \REGISTERS_reg[8][62]  ( .D(n6973), .CK(CLK), .Q(n24476), .QN(n19687)
         );
  DFF_X1 \REGISTERS_reg[8][61]  ( .D(n6972), .CK(CLK), .Q(n24475), .QN(n19688)
         );
  DFF_X1 \REGISTERS_reg[8][60]  ( .D(n6971), .CK(CLK), .Q(n24474), .QN(n19689)
         );
  DFF_X1 \REGISTERS_reg[8][59]  ( .D(n6970), .CK(CLK), .Q(n24853), .QN(n19690)
         );
  DFF_X1 \REGISTERS_reg[8][58]  ( .D(n6969), .CK(CLK), .Q(n24852), .QN(n19691)
         );
  DFF_X1 \REGISTERS_reg[8][57]  ( .D(n6968), .CK(CLK), .Q(n24851), .QN(n19692)
         );
  DFF_X1 \REGISTERS_reg[8][56]  ( .D(n6967), .CK(CLK), .Q(n24850), .QN(n19693)
         );
  DFF_X1 \REGISTERS_reg[8][55]  ( .D(n6966), .CK(CLK), .Q(n24849), .QN(n19694)
         );
  DFF_X1 \REGISTERS_reg[8][54]  ( .D(n6965), .CK(CLK), .Q(n24848), .QN(n19695)
         );
  DFF_X1 \REGISTERS_reg[8][53]  ( .D(n6964), .CK(CLK), .Q(n24847), .QN(n19696)
         );
  DFF_X1 \REGISTERS_reg[8][52]  ( .D(n6963), .CK(CLK), .Q(n24846), .QN(n19697)
         );
  DFF_X1 \REGISTERS_reg[8][51]  ( .D(n6962), .CK(CLK), .Q(n24845), .QN(n19698)
         );
  DFF_X1 \REGISTERS_reg[8][50]  ( .D(n6961), .CK(CLK), .Q(n24844), .QN(n19699)
         );
  DFF_X1 \REGISTERS_reg[8][49]  ( .D(n6960), .CK(CLK), .Q(n24843), .QN(n19700)
         );
  DFF_X1 \REGISTERS_reg[8][48]  ( .D(n6959), .CK(CLK), .Q(n24842), .QN(n19701)
         );
  DFF_X1 \REGISTERS_reg[8][47]  ( .D(n6958), .CK(CLK), .Q(n24841), .QN(n19702)
         );
  DFF_X1 \REGISTERS_reg[8][46]  ( .D(n6957), .CK(CLK), .Q(n24840), .QN(n19703)
         );
  DFF_X1 \REGISTERS_reg[8][45]  ( .D(n6956), .CK(CLK), .Q(n24839), .QN(n19704)
         );
  DFF_X1 \REGISTERS_reg[8][44]  ( .D(n6955), .CK(CLK), .Q(n24838), .QN(n19705)
         );
  DFF_X1 \REGISTERS_reg[8][43]  ( .D(n6954), .CK(CLK), .Q(n24837), .QN(n19706)
         );
  DFF_X1 \REGISTERS_reg[8][42]  ( .D(n6953), .CK(CLK), .Q(n24836), .QN(n19707)
         );
  DFF_X1 \REGISTERS_reg[8][41]  ( .D(n6952), .CK(CLK), .Q(n24835), .QN(n19708)
         );
  DFF_X1 \REGISTERS_reg[8][40]  ( .D(n6951), .CK(CLK), .Q(n24834), .QN(n19709)
         );
  DFF_X1 \REGISTERS_reg[8][39]  ( .D(n6950), .CK(CLK), .Q(n24833), .QN(n19710)
         );
  DFF_X1 \REGISTERS_reg[8][38]  ( .D(n6949), .CK(CLK), .Q(n24832), .QN(n19711)
         );
  DFF_X1 \REGISTERS_reg[8][37]  ( .D(n6948), .CK(CLK), .Q(n24831), .QN(n19712)
         );
  DFF_X1 \REGISTERS_reg[8][36]  ( .D(n6947), .CK(CLK), .Q(n24830), .QN(n19713)
         );
  DFF_X1 \REGISTERS_reg[8][35]  ( .D(n6946), .CK(CLK), .Q(n24829), .QN(n19714)
         );
  DFF_X1 \REGISTERS_reg[8][34]  ( .D(n6945), .CK(CLK), .Q(n24828), .QN(n19715)
         );
  DFF_X1 \REGISTERS_reg[8][33]  ( .D(n6944), .CK(CLK), .Q(n24827), .QN(n19716)
         );
  DFF_X1 \REGISTERS_reg[8][32]  ( .D(n6943), .CK(CLK), .Q(n24826), .QN(n19717)
         );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n6942), .CK(CLK), .Q(n24825), .QN(n19718)
         );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n6941), .CK(CLK), .Q(n24824), .QN(n19719)
         );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n6940), .CK(CLK), .Q(n24823), .QN(n19720)
         );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n6939), .CK(CLK), .Q(n24822), .QN(n19721)
         );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n6938), .CK(CLK), .Q(n24821), .QN(n19722)
         );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n6937), .CK(CLK), .Q(n24820), .QN(n19723)
         );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n6936), .CK(CLK), .Q(n24819), .QN(n19724)
         );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n6935), .CK(CLK), .Q(n24818), .QN(n19725)
         );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n6934), .CK(CLK), .Q(n24817), .QN(n19726)
         );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n6933), .CK(CLK), .Q(n24816), .QN(n19727)
         );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n6932), .CK(CLK), .Q(n24815), .QN(n19728)
         );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n6931), .CK(CLK), .Q(n24814), .QN(n19729)
         );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n6930), .CK(CLK), .Q(n24813), .QN(n19730)
         );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n6929), .CK(CLK), .Q(n24812), .QN(n19731)
         );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n6928), .CK(CLK), .Q(n24811), .QN(n19732)
         );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n6927), .CK(CLK), .Q(n24810), .QN(n19733)
         );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n6926), .CK(CLK), .Q(n24809), .QN(n19734)
         );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n6925), .CK(CLK), .Q(n24808), .QN(n19735)
         );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n6924), .CK(CLK), .Q(n24807), .QN(n19736)
         );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n6923), .CK(CLK), .Q(n24806), .QN(n19737)
         );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n6922), .CK(CLK), .Q(n24805), .QN(n19738)
         );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n6921), .CK(CLK), .Q(n24804), .QN(n19739)
         );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n6920), .CK(CLK), .Q(n24803), .QN(n19740)
         );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n6919), .CK(CLK), .Q(n24802), .QN(n19741)
         );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n6918), .CK(CLK), .Q(n24801), .QN(n19742)
         );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n6917), .CK(CLK), .Q(n24800), .QN(n19743)
         );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n6916), .CK(CLK), .Q(n24799), .QN(n19744)
         );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n6915), .CK(CLK), .Q(n24798), .QN(n19745)
         );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n6914), .CK(CLK), .Q(n24797), .QN(n19746)
         );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n6913), .CK(CLK), .Q(n24796), .QN(n19747)
         );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n6912), .CK(CLK), .Q(n24795), .QN(n19748)
         );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n6911), .CK(CLK), .Q(n24794), .QN(n19749)
         );
  DFF_X1 \REGISTERS_reg[23][63]  ( .D(n6014), .CK(CLK), .Q(n17157), .QN(n21030) );
  DFF_X1 \REGISTERS_reg[23][62]  ( .D(n6013), .CK(CLK), .Q(n17178), .QN(n21031) );
  DFF_X1 \REGISTERS_reg[23][61]  ( .D(n6012), .CK(CLK), .Q(n17199), .QN(n21032) );
  DFF_X1 \REGISTERS_reg[23][60]  ( .D(n6011), .CK(CLK), .Q(n17220), .QN(n21033) );
  DFF_X1 \REGISTERS_reg[23][59]  ( .D(n6010), .CK(CLK), .Q(n17241), .QN(n21034) );
  DFF_X1 \REGISTERS_reg[23][58]  ( .D(n6009), .CK(CLK), .Q(n17262), .QN(n21035) );
  DFF_X1 \REGISTERS_reg[23][57]  ( .D(n6008), .CK(CLK), .Q(n17283), .QN(n21036) );
  DFF_X1 \REGISTERS_reg[23][56]  ( .D(n6007), .CK(CLK), .Q(n17304), .QN(n21037) );
  DFF_X1 \REGISTERS_reg[23][55]  ( .D(n6006), .CK(CLK), .Q(n17325), .QN(n21038) );
  DFF_X1 \REGISTERS_reg[23][54]  ( .D(n6005), .CK(CLK), .Q(n17346), .QN(n21039) );
  DFF_X1 \REGISTERS_reg[23][53]  ( .D(n6004), .CK(CLK), .Q(n17367), .QN(n21040) );
  DFF_X1 \REGISTERS_reg[23][52]  ( .D(n6003), .CK(CLK), .Q(n17388), .QN(n21041) );
  DFF_X1 \REGISTERS_reg[23][51]  ( .D(n6002), .CK(CLK), .Q(n17409), .QN(n21042) );
  DFF_X1 \REGISTERS_reg[23][50]  ( .D(n6001), .CK(CLK), .Q(n17430), .QN(n21043) );
  DFF_X1 \REGISTERS_reg[23][49]  ( .D(n6000), .CK(CLK), .Q(n17451), .QN(n21044) );
  DFF_X1 \REGISTERS_reg[23][48]  ( .D(n5999), .CK(CLK), .Q(n17472), .QN(n21045) );
  DFF_X1 \REGISTERS_reg[23][47]  ( .D(n5998), .CK(CLK), .Q(n17493), .QN(n21046) );
  DFF_X1 \REGISTERS_reg[23][46]  ( .D(n5997), .CK(CLK), .Q(n17514), .QN(n21047) );
  DFF_X1 \REGISTERS_reg[23][45]  ( .D(n5996), .CK(CLK), .Q(n17535), .QN(n21048) );
  DFF_X1 \REGISTERS_reg[23][44]  ( .D(n5995), .CK(CLK), .Q(n17556), .QN(n21049) );
  DFF_X1 \REGISTERS_reg[23][43]  ( .D(n5994), .CK(CLK), .Q(n17577), .QN(n21050) );
  DFF_X1 \REGISTERS_reg[23][42]  ( .D(n5993), .CK(CLK), .Q(n17598), .QN(n21051) );
  DFF_X1 \REGISTERS_reg[23][41]  ( .D(n5992), .CK(CLK), .Q(n17619), .QN(n21052) );
  DFF_X1 \REGISTERS_reg[23][40]  ( .D(n5991), .CK(CLK), .Q(n17640), .QN(n21053) );
  DFF_X1 \REGISTERS_reg[23][39]  ( .D(n5990), .CK(CLK), .Q(n17661), .QN(n21054) );
  DFF_X1 \REGISTERS_reg[23][38]  ( .D(n5989), .CK(CLK), .Q(n17682), .QN(n21055) );
  DFF_X1 \REGISTERS_reg[23][37]  ( .D(n5988), .CK(CLK), .Q(n17703), .QN(n21056) );
  DFF_X1 \REGISTERS_reg[23][36]  ( .D(n5987), .CK(CLK), .Q(n17724), .QN(n21057) );
  DFF_X1 \REGISTERS_reg[23][35]  ( .D(n5986), .CK(CLK), .Q(n17745), .QN(n21058) );
  DFF_X1 \REGISTERS_reg[23][34]  ( .D(n5985), .CK(CLK), .Q(n17766), .QN(n21059) );
  DFF_X1 \REGISTERS_reg[23][33]  ( .D(n5984), .CK(CLK), .Q(n17787), .QN(n21060) );
  DFF_X1 \REGISTERS_reg[23][32]  ( .D(n5983), .CK(CLK), .Q(n17808), .QN(n21061) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n5982), .CK(CLK), .Q(n17829), .QN(n21062) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n5981), .CK(CLK), .Q(n17850), .QN(n21063) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n5980), .CK(CLK), .Q(n17871), .QN(n21064) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n5979), .CK(CLK), .Q(n17892), .QN(n21065) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n5978), .CK(CLK), .Q(n17913), .QN(n21066) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n5977), .CK(CLK), .Q(n17934), .QN(n21067) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n5976), .CK(CLK), .Q(n17955), .QN(n21068) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n5975), .CK(CLK), .Q(n17976), .QN(n21069) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n5974), .CK(CLK), .Q(n17997), .QN(n21070) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n5973), .CK(CLK), .Q(n18018), .QN(n21071) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n5972), .CK(CLK), .Q(n18039), .QN(n21072) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n5971), .CK(CLK), .Q(n18060), .QN(n21073) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n5970), .CK(CLK), .Q(n18081), .QN(n21074) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n5969), .CK(CLK), .Q(n18102), .QN(n21075) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n5968), .CK(CLK), .Q(n18123), .QN(n21076) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n5967), .CK(CLK), .Q(n18144), .QN(n21077) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n5966), .CK(CLK), .Q(n18165), .QN(n21078) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n5965), .CK(CLK), .Q(n18186), .QN(n21079) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n5964), .CK(CLK), .Q(n18207), .QN(n21080) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n5963), .CK(CLK), .Q(n18228), .QN(n21081) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n5962), .CK(CLK), .Q(n18249), .QN(n21082) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n5961), .CK(CLK), .Q(n18270), .QN(n21083) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n5960), .CK(CLK), .Q(n18291), .QN(n21084)
         );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n5959), .CK(CLK), .Q(n18312), .QN(n21085)
         );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n5958), .CK(CLK), .Q(n18333), .QN(n21086)
         );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n5957), .CK(CLK), .Q(n18354), .QN(n21087)
         );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n5956), .CK(CLK), .Q(n18375), .QN(n21088)
         );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n5955), .CK(CLK), .Q(n18396), .QN(n21089)
         );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n5954), .CK(CLK), .Q(n18417), .QN(n21090)
         );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n5953), .CK(CLK), .Q(n18438), .QN(n21091)
         );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n5952), .CK(CLK), .Q(n18459), .QN(n21092)
         );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n5951), .CK(CLK), .Q(n18480), .QN(n21093)
         );
  DFF_X1 \REGISTERS_reg[16][63]  ( .D(n6462), .CK(CLK), .Q(n17148), .QN(n20902) );
  DFF_X1 \REGISTERS_reg[16][62]  ( .D(n6461), .CK(CLK), .Q(n17169), .QN(n20903) );
  DFF_X1 \REGISTERS_reg[16][61]  ( .D(n6460), .CK(CLK), .Q(n17190), .QN(n20904) );
  DFF_X1 \REGISTERS_reg[16][60]  ( .D(n6459), .CK(CLK), .Q(n17211), .QN(n20905) );
  DFF_X1 \REGISTERS_reg[16][59]  ( .D(n6458), .CK(CLK), .Q(n17232), .QN(n20906) );
  DFF_X1 \REGISTERS_reg[16][58]  ( .D(n6457), .CK(CLK), .Q(n17253), .QN(n20907) );
  DFF_X1 \REGISTERS_reg[16][57]  ( .D(n6456), .CK(CLK), .Q(n17274), .QN(n20908) );
  DFF_X1 \REGISTERS_reg[16][56]  ( .D(n6455), .CK(CLK), .Q(n17295), .QN(n20909) );
  DFF_X1 \REGISTERS_reg[16][55]  ( .D(n6454), .CK(CLK), .Q(n17316), .QN(n20910) );
  DFF_X1 \REGISTERS_reg[16][54]  ( .D(n6453), .CK(CLK), .Q(n17337), .QN(n20911) );
  DFF_X1 \REGISTERS_reg[16][53]  ( .D(n6452), .CK(CLK), .Q(n17358), .QN(n20912) );
  DFF_X1 \REGISTERS_reg[16][52]  ( .D(n6451), .CK(CLK), .Q(n17379), .QN(n20913) );
  DFF_X1 \REGISTERS_reg[16][51]  ( .D(n6450), .CK(CLK), .Q(n17400), .QN(n20914) );
  DFF_X1 \REGISTERS_reg[16][50]  ( .D(n6449), .CK(CLK), .Q(n17421), .QN(n20915) );
  DFF_X1 \REGISTERS_reg[16][49]  ( .D(n6448), .CK(CLK), .Q(n17442), .QN(n20916) );
  DFF_X1 \REGISTERS_reg[16][48]  ( .D(n6447), .CK(CLK), .Q(n17463), .QN(n20917) );
  DFF_X1 \REGISTERS_reg[16][47]  ( .D(n6446), .CK(CLK), .Q(n17484), .QN(n20918) );
  DFF_X1 \REGISTERS_reg[16][46]  ( .D(n6445), .CK(CLK), .Q(n17505), .QN(n20919) );
  DFF_X1 \REGISTERS_reg[16][45]  ( .D(n6444), .CK(CLK), .Q(n17526), .QN(n20920) );
  DFF_X1 \REGISTERS_reg[16][44]  ( .D(n6443), .CK(CLK), .Q(n17547), .QN(n20921) );
  DFF_X1 \REGISTERS_reg[16][43]  ( .D(n6442), .CK(CLK), .Q(n17568), .QN(n20922) );
  DFF_X1 \REGISTERS_reg[16][42]  ( .D(n6441), .CK(CLK), .Q(n17589), .QN(n20923) );
  DFF_X1 \REGISTERS_reg[16][41]  ( .D(n6440), .CK(CLK), .Q(n17610), .QN(n20924) );
  DFF_X1 \REGISTERS_reg[16][40]  ( .D(n6439), .CK(CLK), .Q(n17631), .QN(n20925) );
  DFF_X1 \REGISTERS_reg[16][39]  ( .D(n6438), .CK(CLK), .Q(n17652), .QN(n20926) );
  DFF_X1 \REGISTERS_reg[16][38]  ( .D(n6437), .CK(CLK), .Q(n17673), .QN(n20927) );
  DFF_X1 \REGISTERS_reg[16][37]  ( .D(n6436), .CK(CLK), .Q(n17694), .QN(n20928) );
  DFF_X1 \REGISTERS_reg[16][36]  ( .D(n6435), .CK(CLK), .Q(n17715), .QN(n20929) );
  DFF_X1 \REGISTERS_reg[16][35]  ( .D(n6434), .CK(CLK), .Q(n17736), .QN(n20930) );
  DFF_X1 \REGISTERS_reg[16][34]  ( .D(n6433), .CK(CLK), .Q(n17757), .QN(n20931) );
  DFF_X1 \REGISTERS_reg[16][33]  ( .D(n6432), .CK(CLK), .Q(n17778), .QN(n20932) );
  DFF_X1 \REGISTERS_reg[16][32]  ( .D(n6431), .CK(CLK), .Q(n17799), .QN(n20933) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n6430), .CK(CLK), .Q(n17820), .QN(n20934) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n6429), .CK(CLK), .Q(n17841), .QN(n20935) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n6428), .CK(CLK), .Q(n17862), .QN(n20936) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n6427), .CK(CLK), .Q(n17883), .QN(n20937) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n6426), .CK(CLK), .Q(n17904), .QN(n20938) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n6425), .CK(CLK), .Q(n17925), .QN(n20939) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n6424), .CK(CLK), .Q(n17946), .QN(n20940) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n6423), .CK(CLK), .Q(n17967), .QN(n20941) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n6422), .CK(CLK), .Q(n17988), .QN(n20942) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n6421), .CK(CLK), .Q(n18009), .QN(n20943) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n6420), .CK(CLK), .Q(n18030), .QN(n20944) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n6419), .CK(CLK), .Q(n18051), .QN(n20945) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n6418), .CK(CLK), .Q(n18072), .QN(n20946) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n6417), .CK(CLK), .Q(n18093), .QN(n20947) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n6416), .CK(CLK), .Q(n18114), .QN(n20948) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n6415), .CK(CLK), .Q(n18135), .QN(n20949) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n6414), .CK(CLK), .Q(n18156), .QN(n20950) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n6413), .CK(CLK), .Q(n18177), .QN(n20951) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n6412), .CK(CLK), .Q(n18198), .QN(n20952) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n6411), .CK(CLK), .Q(n18219), .QN(n20953) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n6410), .CK(CLK), .Q(n18240), .QN(n20954) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n6409), .CK(CLK), .Q(n18261), .QN(n20955) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n6408), .CK(CLK), .Q(n18282), .QN(n20956)
         );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n6407), .CK(CLK), .Q(n18303), .QN(n20957)
         );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n6406), .CK(CLK), .Q(n18324), .QN(n20958)
         );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n6405), .CK(CLK), .Q(n18345), .QN(n20959)
         );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n6404), .CK(CLK), .Q(n18366), .QN(n20960)
         );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n6403), .CK(CLK), .Q(n18387), .QN(n20961)
         );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n6402), .CK(CLK), .Q(n18408), .QN(n20962)
         );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n6401), .CK(CLK), .Q(n18429), .QN(n20963)
         );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n6400), .CK(CLK), .Q(n18450), .QN(n20964)
         );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n6399), .CK(CLK), .Q(n18471), .QN(n20965)
         );
  DFF_X1 \REGISTERS_reg[14][63]  ( .D(n6590), .CK(CLK), .Q(n17149), .QN(n21414) );
  DFF_X1 \REGISTERS_reg[14][62]  ( .D(n6589), .CK(CLK), .Q(n17170), .QN(n21415) );
  DFF_X1 \REGISTERS_reg[14][61]  ( .D(n6588), .CK(CLK), .Q(n17191), .QN(n21416) );
  DFF_X1 \REGISTERS_reg[14][60]  ( .D(n6587), .CK(CLK), .Q(n17212), .QN(n21417) );
  DFF_X1 \REGISTERS_reg[14][59]  ( .D(n6586), .CK(CLK), .Q(n17233), .QN(n21418) );
  DFF_X1 \REGISTERS_reg[14][58]  ( .D(n6585), .CK(CLK), .Q(n17254), .QN(n21419) );
  DFF_X1 \REGISTERS_reg[14][57]  ( .D(n6584), .CK(CLK), .Q(n17275), .QN(n21420) );
  DFF_X1 \REGISTERS_reg[14][56]  ( .D(n6583), .CK(CLK), .Q(n17296), .QN(n21421) );
  DFF_X1 \REGISTERS_reg[14][55]  ( .D(n6582), .CK(CLK), .Q(n17317), .QN(n21422) );
  DFF_X1 \REGISTERS_reg[14][54]  ( .D(n6581), .CK(CLK), .Q(n17338), .QN(n21423) );
  DFF_X1 \REGISTERS_reg[14][53]  ( .D(n6580), .CK(CLK), .Q(n17359), .QN(n21424) );
  DFF_X1 \REGISTERS_reg[14][52]  ( .D(n6579), .CK(CLK), .Q(n17380), .QN(n21425) );
  DFF_X1 \REGISTERS_reg[14][51]  ( .D(n6578), .CK(CLK), .Q(n17401), .QN(n21426) );
  DFF_X1 \REGISTERS_reg[14][50]  ( .D(n6577), .CK(CLK), .Q(n17422), .QN(n21427) );
  DFF_X1 \REGISTERS_reg[14][49]  ( .D(n6576), .CK(CLK), .Q(n17443), .QN(n21428) );
  DFF_X1 \REGISTERS_reg[14][48]  ( .D(n6575), .CK(CLK), .Q(n17464), .QN(n21429) );
  DFF_X1 \REGISTERS_reg[14][47]  ( .D(n6574), .CK(CLK), .Q(n17485), .QN(n21430) );
  DFF_X1 \REGISTERS_reg[14][46]  ( .D(n6573), .CK(CLK), .Q(n17506), .QN(n21431) );
  DFF_X1 \REGISTERS_reg[14][45]  ( .D(n6572), .CK(CLK), .Q(n17527), .QN(n21432) );
  DFF_X1 \REGISTERS_reg[14][44]  ( .D(n6571), .CK(CLK), .Q(n17548), .QN(n21433) );
  DFF_X1 \REGISTERS_reg[14][43]  ( .D(n6570), .CK(CLK), .Q(n17569), .QN(n21434) );
  DFF_X1 \REGISTERS_reg[14][42]  ( .D(n6569), .CK(CLK), .Q(n17590), .QN(n21435) );
  DFF_X1 \REGISTERS_reg[14][41]  ( .D(n6568), .CK(CLK), .Q(n17611), .QN(n21436) );
  DFF_X1 \REGISTERS_reg[14][40]  ( .D(n6567), .CK(CLK), .Q(n17632), .QN(n21437) );
  DFF_X1 \REGISTERS_reg[14][39]  ( .D(n6566), .CK(CLK), .Q(n17653), .QN(n21438) );
  DFF_X1 \REGISTERS_reg[14][38]  ( .D(n6565), .CK(CLK), .Q(n17674), .QN(n21439) );
  DFF_X1 \REGISTERS_reg[14][37]  ( .D(n6564), .CK(CLK), .Q(n17695), .QN(n21440) );
  DFF_X1 \REGISTERS_reg[14][36]  ( .D(n6563), .CK(CLK), .Q(n17716), .QN(n21441) );
  DFF_X1 \REGISTERS_reg[14][35]  ( .D(n6562), .CK(CLK), .Q(n17737), .QN(n21442) );
  DFF_X1 \REGISTERS_reg[14][34]  ( .D(n6561), .CK(CLK), .Q(n17758), .QN(n21443) );
  DFF_X1 \REGISTERS_reg[14][33]  ( .D(n6560), .CK(CLK), .Q(n17779), .QN(n21444) );
  DFF_X1 \REGISTERS_reg[14][32]  ( .D(n6559), .CK(CLK), .Q(n17800), .QN(n21445) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n6558), .CK(CLK), .Q(n17821), .QN(n21446) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n6557), .CK(CLK), .Q(n17842), .QN(n21447) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n6556), .CK(CLK), .Q(n17863), .QN(n21448) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n6555), .CK(CLK), .Q(n17884), .QN(n21449) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n6554), .CK(CLK), .Q(n17905), .QN(n21450) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n6553), .CK(CLK), .Q(n17926), .QN(n21451) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n6552), .CK(CLK), .Q(n17947), .QN(n21452) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n6551), .CK(CLK), .Q(n17968), .QN(n21453) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n6550), .CK(CLK), .Q(n17989), .QN(n21454) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n6549), .CK(CLK), .Q(n18010), .QN(n21455) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n6548), .CK(CLK), .Q(n18031), .QN(n21456) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n6547), .CK(CLK), .Q(n18052), .QN(n21457) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n6546), .CK(CLK), .Q(n18073), .QN(n21458) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n6545), .CK(CLK), .Q(n18094), .QN(n21459) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n6544), .CK(CLK), .Q(n18115), .QN(n21460) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n6543), .CK(CLK), .Q(n18136), .QN(n21461) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n6542), .CK(CLK), .Q(n18157), .QN(n21462) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n6541), .CK(CLK), .Q(n18178), .QN(n21463) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n6540), .CK(CLK), .Q(n18199), .QN(n21464) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n6539), .CK(CLK), .Q(n18220), .QN(n21465) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n6538), .CK(CLK), .Q(n18241), .QN(n21466) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n6537), .CK(CLK), .Q(n18262), .QN(n21467) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n6536), .CK(CLK), .Q(n18283), .QN(n21468)
         );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n6535), .CK(CLK), .Q(n18304), .QN(n21469)
         );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n6534), .CK(CLK), .Q(n18325), .QN(n21470)
         );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n6533), .CK(CLK), .Q(n18346), .QN(n21471)
         );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n6532), .CK(CLK), .Q(n18367), .QN(n21472)
         );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n6531), .CK(CLK), .Q(n18388), .QN(n21473)
         );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n6530), .CK(CLK), .Q(n18409), .QN(n21474)
         );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n6529), .CK(CLK), .Q(n18430), .QN(n21475)
         );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n6528), .CK(CLK), .Q(n18451), .QN(n21476)
         );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n6527), .CK(CLK), .Q(n18472), .QN(n21477)
         );
  DFF_X1 \REGISTERS_reg[30][63]  ( .D(n5566), .CK(CLK), .Q(n24441), .QN(n20262) );
  DFF_X1 \REGISTERS_reg[30][62]  ( .D(n5565), .CK(CLK), .Q(n24439), .QN(n20263) );
  DFF_X1 \REGISTERS_reg[30][61]  ( .D(n5564), .CK(CLK), .Q(n24437), .QN(n20264) );
  DFF_X1 \REGISTERS_reg[30][60]  ( .D(n5563), .CK(CLK), .Q(n24435), .QN(n20265) );
  DFF_X1 \REGISTERS_reg[28][63]  ( .D(n5694), .CK(CLK), .Q(n24085), .QN(n20266) );
  DFF_X1 \REGISTERS_reg[28][62]  ( .D(n5693), .CK(CLK), .Q(n24083), .QN(n20267) );
  DFF_X1 \REGISTERS_reg[28][61]  ( .D(n5692), .CK(CLK), .Q(n24081), .QN(n20268) );
  DFF_X1 \REGISTERS_reg[28][60]  ( .D(n5691), .CK(CLK), .Q(n24079), .QN(n20269) );
  DFF_X1 \REGISTERS_reg[30][59]  ( .D(n5562), .CK(CLK), .Q(n24433), .QN(n20462) );
  DFF_X1 \REGISTERS_reg[30][58]  ( .D(n5561), .CK(CLK), .Q(n24431), .QN(n20463) );
  DFF_X1 \REGISTERS_reg[30][57]  ( .D(n5560), .CK(CLK), .Q(n24429), .QN(n20464) );
  DFF_X1 \REGISTERS_reg[30][56]  ( .D(n5559), .CK(CLK), .Q(n24427), .QN(n20465) );
  DFF_X1 \REGISTERS_reg[30][55]  ( .D(n5558), .CK(CLK), .Q(n24425), .QN(n20466) );
  DFF_X1 \REGISTERS_reg[30][54]  ( .D(n5557), .CK(CLK), .Q(n24423), .QN(n20467) );
  DFF_X1 \REGISTERS_reg[30][53]  ( .D(n5556), .CK(CLK), .Q(n24421), .QN(n20468) );
  DFF_X1 \REGISTERS_reg[30][52]  ( .D(n5555), .CK(CLK), .Q(n24419), .QN(n20469) );
  DFF_X1 \REGISTERS_reg[30][51]  ( .D(n5554), .CK(CLK), .Q(n24417), .QN(n20470) );
  DFF_X1 \REGISTERS_reg[30][50]  ( .D(n5553), .CK(CLK), .Q(n24415), .QN(n20471) );
  DFF_X1 \REGISTERS_reg[30][49]  ( .D(n5552), .CK(CLK), .Q(n24413), .QN(n20472) );
  DFF_X1 \REGISTERS_reg[30][48]  ( .D(n5551), .CK(CLK), .Q(n24411), .QN(n20473) );
  DFF_X1 \REGISTERS_reg[30][47]  ( .D(n5550), .CK(CLK), .Q(n24409), .QN(n20474) );
  DFF_X1 \REGISTERS_reg[30][46]  ( .D(n5549), .CK(CLK), .Q(n24407), .QN(n20475) );
  DFF_X1 \REGISTERS_reg[30][45]  ( .D(n5548), .CK(CLK), .Q(n24405), .QN(n20476) );
  DFF_X1 \REGISTERS_reg[30][44]  ( .D(n5547), .CK(CLK), .Q(n24403), .QN(n20477) );
  DFF_X1 \REGISTERS_reg[30][43]  ( .D(n5546), .CK(CLK), .Q(n24401), .QN(n20478) );
  DFF_X1 \REGISTERS_reg[30][42]  ( .D(n5545), .CK(CLK), .Q(n24399), .QN(n20479) );
  DFF_X1 \REGISTERS_reg[30][41]  ( .D(n5544), .CK(CLK), .Q(n24397), .QN(n20480) );
  DFF_X1 \REGISTERS_reg[30][40]  ( .D(n5543), .CK(CLK), .Q(n24395), .QN(n20481) );
  DFF_X1 \REGISTERS_reg[30][39]  ( .D(n5542), .CK(CLK), .Q(n24393), .QN(n20482) );
  DFF_X1 \REGISTERS_reg[30][38]  ( .D(n5541), .CK(CLK), .Q(n24391), .QN(n20483) );
  DFF_X1 \REGISTERS_reg[30][37]  ( .D(n5540), .CK(CLK), .Q(n24389), .QN(n20484) );
  DFF_X1 \REGISTERS_reg[30][36]  ( .D(n5539), .CK(CLK), .Q(n24387), .QN(n20485) );
  DFF_X1 \REGISTERS_reg[30][35]  ( .D(n5538), .CK(CLK), .Q(n24385), .QN(n20486) );
  DFF_X1 \REGISTERS_reg[30][34]  ( .D(n5537), .CK(CLK), .Q(n24383), .QN(n20487) );
  DFF_X1 \REGISTERS_reg[30][33]  ( .D(n5536), .CK(CLK), .Q(n24381), .QN(n20488) );
  DFF_X1 \REGISTERS_reg[30][32]  ( .D(n5535), .CK(CLK), .Q(n24379), .QN(n20489) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n5534), .CK(CLK), .Q(n24377), .QN(n20490) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n5533), .CK(CLK), .Q(n24375), .QN(n20491) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n5532), .CK(CLK), .Q(n24373), .QN(n20492) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n5531), .CK(CLK), .Q(n24371), .QN(n20493) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n5530), .CK(CLK), .Q(n24369), .QN(n20494) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n5529), .CK(CLK), .Q(n24367), .QN(n20495) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n5528), .CK(CLK), .Q(n24365), .QN(n20496) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n5527), .CK(CLK), .Q(n24363), .QN(n20497) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n5526), .CK(CLK), .Q(n24361), .QN(n20498) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n5525), .CK(CLK), .Q(n24359), .QN(n20499) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n5524), .CK(CLK), .Q(n24357), .QN(n20500) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n5523), .CK(CLK), .Q(n24355), .QN(n20501) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n5522), .CK(CLK), .Q(n24353), .QN(n20502) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n5521), .CK(CLK), .Q(n24351), .QN(n20503) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n5520), .CK(CLK), .Q(n24349), .QN(n20504) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n5519), .CK(CLK), .Q(n24347), .QN(n20505) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n5518), .CK(CLK), .Q(n24345), .QN(n20506) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n5517), .CK(CLK), .Q(n24343), .QN(n20507) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n5516), .CK(CLK), .Q(n24341), .QN(n20508) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n5515), .CK(CLK), .Q(n24339), .QN(n20509) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n5514), .CK(CLK), .Q(n24465), .QN(n20510) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n5513), .CK(CLK), .Q(n24463), .QN(n20511) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n5512), .CK(CLK), .Q(n24461), .QN(n20512)
         );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n5511), .CK(CLK), .Q(n24459), .QN(n20513)
         );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n5510), .CK(CLK), .Q(n24457), .QN(n20514)
         );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n5509), .CK(CLK), .Q(n24455), .QN(n20515)
         );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n5508), .CK(CLK), .Q(n24453), .QN(n20516)
         );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n5507), .CK(CLK), .Q(n24451), .QN(n20517)
         );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n5506), .CK(CLK), .Q(n24449), .QN(n20518)
         );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n5505), .CK(CLK), .Q(n24447), .QN(n20519)
         );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n5504), .CK(CLK), .Q(n24445), .QN(n20520)
         );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n5503), .CK(CLK), .Q(n24443), .QN(n20521)
         );
  DFF_X1 \REGISTERS_reg[28][59]  ( .D(n5690), .CK(CLK), .Q(n24205), .QN(n20522) );
  DFF_X1 \REGISTERS_reg[28][58]  ( .D(n5689), .CK(CLK), .Q(n24203), .QN(n20523) );
  DFF_X1 \REGISTERS_reg[28][57]  ( .D(n5688), .CK(CLK), .Q(n24201), .QN(n20524) );
  DFF_X1 \REGISTERS_reg[28][56]  ( .D(n5687), .CK(CLK), .Q(n24199), .QN(n20525) );
  DFF_X1 \REGISTERS_reg[28][55]  ( .D(n5686), .CK(CLK), .Q(n24197), .QN(n20526) );
  DFF_X1 \REGISTERS_reg[28][54]  ( .D(n5685), .CK(CLK), .Q(n24195), .QN(n20527) );
  DFF_X1 \REGISTERS_reg[28][53]  ( .D(n5684), .CK(CLK), .Q(n24193), .QN(n20528) );
  DFF_X1 \REGISTERS_reg[28][52]  ( .D(n5683), .CK(CLK), .Q(n24191), .QN(n20529) );
  DFF_X1 \REGISTERS_reg[28][51]  ( .D(n5682), .CK(CLK), .Q(n24189), .QN(n20530) );
  DFF_X1 \REGISTERS_reg[28][50]  ( .D(n5681), .CK(CLK), .Q(n24187), .QN(n20531) );
  DFF_X1 \REGISTERS_reg[28][49]  ( .D(n5680), .CK(CLK), .Q(n24185), .QN(n20532) );
  DFF_X1 \REGISTERS_reg[28][48]  ( .D(n5679), .CK(CLK), .Q(n24183), .QN(n20533) );
  DFF_X1 \REGISTERS_reg[28][47]  ( .D(n5678), .CK(CLK), .Q(n24181), .QN(n20534) );
  DFF_X1 \REGISTERS_reg[28][46]  ( .D(n5677), .CK(CLK), .Q(n24179), .QN(n20535) );
  DFF_X1 \REGISTERS_reg[28][45]  ( .D(n5676), .CK(CLK), .Q(n24177), .QN(n20536) );
  DFF_X1 \REGISTERS_reg[28][44]  ( .D(n5675), .CK(CLK), .Q(n24175), .QN(n20537) );
  DFF_X1 \REGISTERS_reg[28][43]  ( .D(n5674), .CK(CLK), .Q(n24173), .QN(n20538) );
  DFF_X1 \REGISTERS_reg[28][42]  ( .D(n5673), .CK(CLK), .Q(n24171), .QN(n20539) );
  DFF_X1 \REGISTERS_reg[28][41]  ( .D(n5672), .CK(CLK), .Q(n24169), .QN(n20540) );
  DFF_X1 \REGISTERS_reg[28][40]  ( .D(n5671), .CK(CLK), .Q(n24167), .QN(n20541) );
  DFF_X1 \REGISTERS_reg[28][39]  ( .D(n5670), .CK(CLK), .Q(n24165), .QN(n20542) );
  DFF_X1 \REGISTERS_reg[28][38]  ( .D(n5669), .CK(CLK), .Q(n24163), .QN(n20543) );
  DFF_X1 \REGISTERS_reg[28][37]  ( .D(n5668), .CK(CLK), .Q(n24161), .QN(n20544) );
  DFF_X1 \REGISTERS_reg[28][36]  ( .D(n5667), .CK(CLK), .Q(n24159), .QN(n20545) );
  DFF_X1 \REGISTERS_reg[28][35]  ( .D(n5666), .CK(CLK), .Q(n24157), .QN(n20546) );
  DFF_X1 \REGISTERS_reg[28][34]  ( .D(n5665), .CK(CLK), .Q(n24155), .QN(n20547) );
  DFF_X1 \REGISTERS_reg[28][33]  ( .D(n5664), .CK(CLK), .Q(n24153), .QN(n20548) );
  DFF_X1 \REGISTERS_reg[28][32]  ( .D(n5663), .CK(CLK), .Q(n24151), .QN(n20549) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n5662), .CK(CLK), .Q(n24149), .QN(n20550) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n5661), .CK(CLK), .Q(n24147), .QN(n20551) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n5660), .CK(CLK), .Q(n24145), .QN(n20552) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n5659), .CK(CLK), .Q(n24143), .QN(n20553) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n5658), .CK(CLK), .Q(n24141), .QN(n20554) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n5657), .CK(CLK), .Q(n24139), .QN(n20555) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n5656), .CK(CLK), .Q(n24137), .QN(n20556) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n5655), .CK(CLK), .Q(n24135), .QN(n20557) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n5654), .CK(CLK), .Q(n24133), .QN(n20558) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n5653), .CK(CLK), .Q(n24131), .QN(n20559) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n5652), .CK(CLK), .Q(n24129), .QN(n20560) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n5651), .CK(CLK), .Q(n24127), .QN(n20561) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n5650), .CK(CLK), .Q(n24125), .QN(n20562) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n5649), .CK(CLK), .Q(n24123), .QN(n20563) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n5648), .CK(CLK), .Q(n24121), .QN(n20564) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n5647), .CK(CLK), .Q(n24119), .QN(n20565) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n5646), .CK(CLK), .Q(n24117), .QN(n20566) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n5645), .CK(CLK), .Q(n24115), .QN(n20567) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n5644), .CK(CLK), .Q(n24113), .QN(n20568) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n5643), .CK(CLK), .Q(n24111), .QN(n20569) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n5642), .CK(CLK), .Q(n24109), .QN(n20570) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n5641), .CK(CLK), .Q(n24107), .QN(n20571) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n5640), .CK(CLK), .Q(n24105), .QN(n20572)
         );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n5639), .CK(CLK), .Q(n24103), .QN(n20573)
         );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n5638), .CK(CLK), .Q(n24101), .QN(n20574)
         );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n5637), .CK(CLK), .Q(n24099), .QN(n20575)
         );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n5636), .CK(CLK), .Q(n24097), .QN(n20576)
         );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n5635), .CK(CLK), .Q(n24095), .QN(n20577)
         );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n5634), .CK(CLK), .Q(n24093), .QN(n20578)
         );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n5633), .CK(CLK), .Q(n24091), .QN(n20579)
         );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n5632), .CK(CLK), .Q(n24089), .QN(n20580)
         );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n5631), .CK(CLK), .Q(n24087), .QN(n20581)
         );
  DFF_X1 \REGISTERS_reg[10][63]  ( .D(n6846), .CK(CLK), .Q(n23957), .QN(n20582) );
  DFF_X1 \REGISTERS_reg[10][62]  ( .D(n6845), .CK(CLK), .Q(n23956), .QN(n20583) );
  DFF_X1 \REGISTERS_reg[10][61]  ( .D(n6844), .CK(CLK), .Q(n23955), .QN(n20584) );
  DFF_X1 \REGISTERS_reg[10][60]  ( .D(n6843), .CK(CLK), .Q(n23954), .QN(n20585) );
  DFF_X1 \REGISTERS_reg[10][59]  ( .D(n6842), .CK(CLK), .Q(n24077), .QN(n20586) );
  DFF_X1 \REGISTERS_reg[10][58]  ( .D(n6841), .CK(CLK), .Q(n24076), .QN(n20587) );
  DFF_X1 \REGISTERS_reg[10][57]  ( .D(n6840), .CK(CLK), .Q(n24075), .QN(n20588) );
  DFF_X1 \REGISTERS_reg[10][56]  ( .D(n6839), .CK(CLK), .Q(n24074), .QN(n20589) );
  DFF_X1 \REGISTERS_reg[10][55]  ( .D(n6838), .CK(CLK), .Q(n24073), .QN(n20590) );
  DFF_X1 \REGISTERS_reg[10][54]  ( .D(n6837), .CK(CLK), .Q(n24072), .QN(n20591) );
  DFF_X1 \REGISTERS_reg[10][53]  ( .D(n6836), .CK(CLK), .Q(n24071), .QN(n20592) );
  DFF_X1 \REGISTERS_reg[10][52]  ( .D(n6835), .CK(CLK), .Q(n24070), .QN(n20593) );
  DFF_X1 \REGISTERS_reg[10][51]  ( .D(n6834), .CK(CLK), .Q(n24069), .QN(n20594) );
  DFF_X1 \REGISTERS_reg[10][50]  ( .D(n6833), .CK(CLK), .Q(n24068), .QN(n20595) );
  DFF_X1 \REGISTERS_reg[10][49]  ( .D(n6832), .CK(CLK), .Q(n24067), .QN(n20596) );
  DFF_X1 \REGISTERS_reg[10][48]  ( .D(n6831), .CK(CLK), .Q(n24066), .QN(n20597) );
  DFF_X1 \REGISTERS_reg[10][47]  ( .D(n6830), .CK(CLK), .Q(n24065), .QN(n20598) );
  DFF_X1 \REGISTERS_reg[10][46]  ( .D(n6829), .CK(CLK), .Q(n24064), .QN(n20599) );
  DFF_X1 \REGISTERS_reg[10][45]  ( .D(n6828), .CK(CLK), .Q(n24063), .QN(n20600) );
  DFF_X1 \REGISTERS_reg[10][44]  ( .D(n6827), .CK(CLK), .Q(n24062), .QN(n20601) );
  DFF_X1 \REGISTERS_reg[10][43]  ( .D(n6826), .CK(CLK), .Q(n24061), .QN(n20602) );
  DFF_X1 \REGISTERS_reg[10][42]  ( .D(n6825), .CK(CLK), .Q(n24060), .QN(n20603) );
  DFF_X1 \REGISTERS_reg[10][41]  ( .D(n6824), .CK(CLK), .Q(n24059), .QN(n20604) );
  DFF_X1 \REGISTERS_reg[10][40]  ( .D(n6823), .CK(CLK), .Q(n24058), .QN(n20605) );
  DFF_X1 \REGISTERS_reg[10][39]  ( .D(n6822), .CK(CLK), .Q(n24057), .QN(n20606) );
  DFF_X1 \REGISTERS_reg[10][38]  ( .D(n6821), .CK(CLK), .Q(n24056), .QN(n20607) );
  DFF_X1 \REGISTERS_reg[10][37]  ( .D(n6820), .CK(CLK), .Q(n24055), .QN(n20608) );
  DFF_X1 \REGISTERS_reg[10][36]  ( .D(n6819), .CK(CLK), .Q(n24054), .QN(n20609) );
  DFF_X1 \REGISTERS_reg[10][35]  ( .D(n6818), .CK(CLK), .Q(n24053), .QN(n20610) );
  DFF_X1 \REGISTERS_reg[10][34]  ( .D(n6817), .CK(CLK), .Q(n24052), .QN(n20611) );
  DFF_X1 \REGISTERS_reg[10][33]  ( .D(n6816), .CK(CLK), .Q(n24051), .QN(n20612) );
  DFF_X1 \REGISTERS_reg[10][32]  ( .D(n6815), .CK(CLK), .Q(n24050), .QN(n20613) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n6814), .CK(CLK), .Q(n24049), .QN(n20614) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n6813), .CK(CLK), .Q(n24048), .QN(n20615) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n6812), .CK(CLK), .Q(n24047), .QN(n20616) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n6811), .CK(CLK), .Q(n24046), .QN(n20617) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n6810), .CK(CLK), .Q(n24045), .QN(n20618) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n6809), .CK(CLK), .Q(n24044), .QN(n20619) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n6808), .CK(CLK), .Q(n24043), .QN(n20620) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n6807), .CK(CLK), .Q(n24042), .QN(n20621) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n6806), .CK(CLK), .Q(n24041), .QN(n20622) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n6805), .CK(CLK), .Q(n24040), .QN(n20623) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n6804), .CK(CLK), .Q(n24039), .QN(n20624) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n6803), .CK(CLK), .Q(n24038), .QN(n20625) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n6802), .CK(CLK), .Q(n24037), .QN(n20626) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n6801), .CK(CLK), .Q(n24036), .QN(n20627) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n6800), .CK(CLK), .Q(n24035), .QN(n20628) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n6799), .CK(CLK), .Q(n24034), .QN(n20629) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n6798), .CK(CLK), .Q(n24033), .QN(n20630) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n6797), .CK(CLK), .Q(n24032), .QN(n20631) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n6796), .CK(CLK), .Q(n24031), .QN(n20632) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n6795), .CK(CLK), .Q(n24030), .QN(n20633) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n6794), .CK(CLK), .Q(n24029), .QN(n20634) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n6793), .CK(CLK), .Q(n24028), .QN(n20635) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n6792), .CK(CLK), .Q(n24027), .QN(n20636)
         );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n6791), .CK(CLK), .Q(n24026), .QN(n20637)
         );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n6790), .CK(CLK), .Q(n24025), .QN(n20638)
         );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n6789), .CK(CLK), .Q(n24024), .QN(n20639)
         );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n6788), .CK(CLK), .Q(n24023), .QN(n20640)
         );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n6787), .CK(CLK), .Q(n24022), .QN(n20641)
         );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n6786), .CK(CLK), .Q(n24021), .QN(n20642)
         );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n6785), .CK(CLK), .Q(n24020), .QN(n20643)
         );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n6784), .CK(CLK), .Q(n24019), .QN(n20644)
         );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n6783), .CK(CLK), .Q(n24018), .QN(n20645)
         );
  DFF_X1 \REGISTERS_reg[6][63]  ( .D(n7102), .CK(CLK), .Q(n24481), .QN(n19622)
         );
  DFF_X1 \REGISTERS_reg[6][62]  ( .D(n7101), .CK(CLK), .Q(n24480), .QN(n19623)
         );
  DFF_X1 \REGISTERS_reg[6][61]  ( .D(n7100), .CK(CLK), .Q(n24479), .QN(n19624)
         );
  DFF_X1 \REGISTERS_reg[6][60]  ( .D(n7099), .CK(CLK), .Q(n24478), .QN(n19625)
         );
  DFF_X1 \REGISTERS_reg[6][59]  ( .D(n7098), .CK(CLK), .Q(n24913), .QN(n19626)
         );
  DFF_X1 \REGISTERS_reg[6][58]  ( .D(n7097), .CK(CLK), .Q(n24912), .QN(n19627)
         );
  DFF_X1 \REGISTERS_reg[6][57]  ( .D(n7096), .CK(CLK), .Q(n24911), .QN(n19628)
         );
  DFF_X1 \REGISTERS_reg[6][56]  ( .D(n7095), .CK(CLK), .Q(n24910), .QN(n19629)
         );
  DFF_X1 \REGISTERS_reg[6][55]  ( .D(n7094), .CK(CLK), .Q(n24909), .QN(n19630)
         );
  DFF_X1 \REGISTERS_reg[6][54]  ( .D(n7093), .CK(CLK), .Q(n24908), .QN(n19631)
         );
  DFF_X1 \REGISTERS_reg[6][53]  ( .D(n7092), .CK(CLK), .Q(n24907), .QN(n19632)
         );
  DFF_X1 \REGISTERS_reg[6][52]  ( .D(n7091), .CK(CLK), .Q(n24906), .QN(n19633)
         );
  DFF_X1 \REGISTERS_reg[6][51]  ( .D(n7090), .CK(CLK), .Q(n24905), .QN(n19634)
         );
  DFF_X1 \REGISTERS_reg[6][50]  ( .D(n7089), .CK(CLK), .Q(n24904), .QN(n19635)
         );
  DFF_X1 \REGISTERS_reg[6][49]  ( .D(n7088), .CK(CLK), .Q(n24903), .QN(n19636)
         );
  DFF_X1 \REGISTERS_reg[6][48]  ( .D(n7087), .CK(CLK), .Q(n24902), .QN(n19637)
         );
  DFF_X1 \REGISTERS_reg[6][47]  ( .D(n7086), .CK(CLK), .Q(n24901), .QN(n19638)
         );
  DFF_X1 \REGISTERS_reg[6][46]  ( .D(n7085), .CK(CLK), .Q(n24900), .QN(n19639)
         );
  DFF_X1 \REGISTERS_reg[6][45]  ( .D(n7084), .CK(CLK), .Q(n24899), .QN(n19640)
         );
  DFF_X1 \REGISTERS_reg[6][44]  ( .D(n7083), .CK(CLK), .Q(n24898), .QN(n19641)
         );
  DFF_X1 \REGISTERS_reg[6][43]  ( .D(n7082), .CK(CLK), .Q(n24897), .QN(n19642)
         );
  DFF_X1 \REGISTERS_reg[6][42]  ( .D(n7081), .CK(CLK), .Q(n24896), .QN(n19643)
         );
  DFF_X1 \REGISTERS_reg[6][41]  ( .D(n7080), .CK(CLK), .Q(n24895), .QN(n19644)
         );
  DFF_X1 \REGISTERS_reg[6][40]  ( .D(n7079), .CK(CLK), .Q(n24894), .QN(n19645)
         );
  DFF_X1 \REGISTERS_reg[6][39]  ( .D(n7078), .CK(CLK), .Q(n24893), .QN(n19646)
         );
  DFF_X1 \REGISTERS_reg[6][38]  ( .D(n7077), .CK(CLK), .Q(n24892), .QN(n19647)
         );
  DFF_X1 \REGISTERS_reg[6][37]  ( .D(n7076), .CK(CLK), .Q(n24891), .QN(n19648)
         );
  DFF_X1 \REGISTERS_reg[6][36]  ( .D(n7075), .CK(CLK), .Q(n24890), .QN(n19649)
         );
  DFF_X1 \REGISTERS_reg[6][35]  ( .D(n7074), .CK(CLK), .Q(n24889), .QN(n19650)
         );
  DFF_X1 \REGISTERS_reg[6][34]  ( .D(n7073), .CK(CLK), .Q(n24888), .QN(n19651)
         );
  DFF_X1 \REGISTERS_reg[6][33]  ( .D(n7072), .CK(CLK), .Q(n24887), .QN(n19652)
         );
  DFF_X1 \REGISTERS_reg[6][32]  ( .D(n7071), .CK(CLK), .Q(n24886), .QN(n19653)
         );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n7070), .CK(CLK), .Q(n24885), .QN(n19654)
         );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n7069), .CK(CLK), .Q(n24884), .QN(n19655)
         );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n7068), .CK(CLK), .Q(n24883), .QN(n19656)
         );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n7067), .CK(CLK), .Q(n24882), .QN(n19657)
         );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n7066), .CK(CLK), .Q(n24881), .QN(n19658)
         );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n7065), .CK(CLK), .Q(n24880), .QN(n19659)
         );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n7064), .CK(CLK), .Q(n24879), .QN(n19660)
         );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n7063), .CK(CLK), .Q(n24878), .QN(n19661)
         );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n7062), .CK(CLK), .Q(n24877), .QN(n19662)
         );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n7061), .CK(CLK), .Q(n24876), .QN(n19663)
         );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n7060), .CK(CLK), .Q(n24875), .QN(n19664)
         );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n7059), .CK(CLK), .Q(n24874), .QN(n19665)
         );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n7058), .CK(CLK), .Q(n24873), .QN(n19666)
         );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n7057), .CK(CLK), .Q(n24872), .QN(n19667)
         );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n7056), .CK(CLK), .Q(n24871), .QN(n19668)
         );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n7055), .CK(CLK), .Q(n24870), .QN(n19669)
         );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n7054), .CK(CLK), .Q(n24869), .QN(n19670)
         );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n7053), .CK(CLK), .Q(n24868), .QN(n19671)
         );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n7052), .CK(CLK), .Q(n24867), .QN(n19672)
         );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n7051), .CK(CLK), .Q(n24866), .QN(n19673)
         );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n7050), .CK(CLK), .Q(n24865), .QN(n19674)
         );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n7049), .CK(CLK), .Q(n24864), .QN(n19675)
         );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n7048), .CK(CLK), .Q(n24863), .QN(n19676)
         );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n7047), .CK(CLK), .Q(n24862), .QN(n19677)
         );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n7046), .CK(CLK), .Q(n24861), .QN(n19678)
         );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n7045), .CK(CLK), .Q(n24860), .QN(n19679)
         );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n7044), .CK(CLK), .Q(n24859), .QN(n19680)
         );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n7043), .CK(CLK), .Q(n24858), .QN(n19681)
         );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n7042), .CK(CLK), .Q(n24857), .QN(n19682)
         );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n7041), .CK(CLK), .Q(n24856), .QN(n19683)
         );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n7040), .CK(CLK), .Q(n24855), .QN(n19684)
         );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n7039), .CK(CLK), .Q(n24854), .QN(n19685)
         );
  DFF_X1 \REGISTERS_reg[3][63]  ( .D(n7294), .CK(CLK), .Q(n24311), .QN(n20198)
         );
  DFF_X1 \REGISTERS_reg[3][62]  ( .D(n7293), .CK(CLK), .Q(n24308), .QN(n20199)
         );
  DFF_X1 \REGISTERS_reg[3][61]  ( .D(n7292), .CK(CLK), .Q(n24305), .QN(n20200)
         );
  DFF_X1 \REGISTERS_reg[3][60]  ( .D(n7291), .CK(CLK), .Q(n24302), .QN(n20201)
         );
  DFF_X1 \REGISTERS_reg[3][59]  ( .D(n7290), .CK(CLK), .Q(n24300), .QN(n20202)
         );
  DFF_X1 \REGISTERS_reg[3][58]  ( .D(n7289), .CK(CLK), .Q(n24298), .QN(n20203)
         );
  DFF_X1 \REGISTERS_reg[3][57]  ( .D(n7288), .CK(CLK), .Q(n24296), .QN(n20204)
         );
  DFF_X1 \REGISTERS_reg[3][56]  ( .D(n7287), .CK(CLK), .Q(n24294), .QN(n20205)
         );
  DFF_X1 \REGISTERS_reg[3][55]  ( .D(n7286), .CK(CLK), .Q(n24292), .QN(n20206)
         );
  DFF_X1 \REGISTERS_reg[3][54]  ( .D(n7285), .CK(CLK), .Q(n24290), .QN(n20207)
         );
  DFF_X1 \REGISTERS_reg[3][53]  ( .D(n7284), .CK(CLK), .Q(n24288), .QN(n20208)
         );
  DFF_X1 \REGISTERS_reg[3][52]  ( .D(n7283), .CK(CLK), .Q(n24286), .QN(n20209)
         );
  DFF_X1 \REGISTERS_reg[3][51]  ( .D(n7282), .CK(CLK), .Q(n24284), .QN(n20210)
         );
  DFF_X1 \REGISTERS_reg[3][50]  ( .D(n7281), .CK(CLK), .Q(n24282), .QN(n20211)
         );
  DFF_X1 \REGISTERS_reg[3][49]  ( .D(n7280), .CK(CLK), .Q(n24280), .QN(n20212)
         );
  DFF_X1 \REGISTERS_reg[3][48]  ( .D(n7279), .CK(CLK), .Q(n24278), .QN(n20213)
         );
  DFF_X1 \REGISTERS_reg[3][47]  ( .D(n7278), .CK(CLK), .Q(n24276), .QN(n20214)
         );
  DFF_X1 \REGISTERS_reg[3][46]  ( .D(n7277), .CK(CLK), .Q(n24274), .QN(n20215)
         );
  DFF_X1 \REGISTERS_reg[3][45]  ( .D(n7276), .CK(CLK), .Q(n24272), .QN(n20216)
         );
  DFF_X1 \REGISTERS_reg[3][44]  ( .D(n7275), .CK(CLK), .Q(n24270), .QN(n20217)
         );
  DFF_X1 \REGISTERS_reg[3][43]  ( .D(n7274), .CK(CLK), .Q(n24268), .QN(n20218)
         );
  DFF_X1 \REGISTERS_reg[3][42]  ( .D(n7273), .CK(CLK), .Q(n24266), .QN(n20219)
         );
  DFF_X1 \REGISTERS_reg[3][41]  ( .D(n7272), .CK(CLK), .Q(n24264), .QN(n20220)
         );
  DFF_X1 \REGISTERS_reg[3][40]  ( .D(n7271), .CK(CLK), .Q(n24262), .QN(n20221)
         );
  DFF_X1 \REGISTERS_reg[3][39]  ( .D(n7270), .CK(CLK), .Q(n24260), .QN(n20222)
         );
  DFF_X1 \REGISTERS_reg[3][38]  ( .D(n7269), .CK(CLK), .Q(n24258), .QN(n20223)
         );
  DFF_X1 \REGISTERS_reg[3][37]  ( .D(n7268), .CK(CLK), .Q(n24256), .QN(n20224)
         );
  DFF_X1 \REGISTERS_reg[3][36]  ( .D(n7267), .CK(CLK), .Q(n24254), .QN(n20225)
         );
  DFF_X1 \REGISTERS_reg[3][35]  ( .D(n7266), .CK(CLK), .Q(n24252), .QN(n20226)
         );
  DFF_X1 \REGISTERS_reg[3][34]  ( .D(n7265), .CK(CLK), .Q(n24250), .QN(n20227)
         );
  DFF_X1 \REGISTERS_reg[3][33]  ( .D(n7264), .CK(CLK), .Q(n24248), .QN(n20228)
         );
  DFF_X1 \REGISTERS_reg[3][32]  ( .D(n7263), .CK(CLK), .Q(n24246), .QN(n20229)
         );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n7262), .CK(CLK), .Q(n24244), .QN(n20230)
         );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n7261), .CK(CLK), .Q(n24242), .QN(n20231)
         );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n7260), .CK(CLK), .Q(n24240), .QN(n20232)
         );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n7259), .CK(CLK), .Q(n24238), .QN(n20233)
         );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n7258), .CK(CLK), .Q(n24236), .QN(n20234)
         );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n7257), .CK(CLK), .Q(n24234), .QN(n20235)
         );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n7256), .CK(CLK), .Q(n24232), .QN(n20236)
         );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n7255), .CK(CLK), .Q(n24230), .QN(n20237)
         );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n7254), .CK(CLK), .Q(n24228), .QN(n20238)
         );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n7253), .CK(CLK), .Q(n24226), .QN(n20239)
         );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n7252), .CK(CLK), .Q(n24224), .QN(n20240)
         );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n7251), .CK(CLK), .Q(n24222), .QN(n20241)
         );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n7250), .CK(CLK), .Q(n24220), .QN(n20242)
         );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n7249), .CK(CLK), .Q(n24218), .QN(n20243)
         );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n7248), .CK(CLK), .Q(n24216), .QN(n20244)
         );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n7247), .CK(CLK), .Q(n24214), .QN(n20245)
         );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n7246), .CK(CLK), .Q(n24212), .QN(n20246)
         );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n7245), .CK(CLK), .Q(n24210), .QN(n20247)
         );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n7244), .CK(CLK), .Q(n24208), .QN(n20248)
         );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n7243), .CK(CLK), .Q(n24206), .QN(n20249)
         );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n7242), .CK(CLK), .Q(n24336), .QN(n20250)
         );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n7241), .CK(CLK), .Q(n24334), .QN(n20251)
         );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n7240), .CK(CLK), .Q(n24332), .QN(n20252)
         );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n7239), .CK(CLK), .Q(n24330), .QN(n20253)
         );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n7238), .CK(CLK), .Q(n24328), .QN(n20254)
         );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n7237), .CK(CLK), .Q(n24326), .QN(n20255)
         );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n7236), .CK(CLK), .Q(n24324), .QN(n20256)
         );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n7235), .CK(CLK), .Q(n24322), .QN(n20257)
         );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n7234), .CK(CLK), .Q(n24320), .QN(n20258)
         );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n7233), .CK(CLK), .Q(n24318), .QN(n20259)
         );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n7232), .CK(CLK), .Q(n24316), .QN(n20260)
         );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n7231), .CK(CLK), .Q(n24314), .QN(n20261)
         );
  DFF_X1 \REGISTERS_reg[22][63]  ( .D(n6078), .CK(CLK), .Q(n24613), .QN(n19877) );
  DFF_X1 \REGISTERS_reg[22][62]  ( .D(n6077), .CK(CLK), .Q(n24611), .QN(n19878) );
  DFF_X1 \REGISTERS_reg[22][61]  ( .D(n6076), .CK(CLK), .Q(n24609), .QN(n19879) );
  DFF_X1 \REGISTERS_reg[22][60]  ( .D(n6075), .CK(CLK), .Q(n24607), .QN(n19880) );
  DFF_X1 \REGISTERS_reg[22][59]  ( .D(n6074), .CK(CLK), .Q(n24673), .QN(n19881) );
  DFF_X1 \REGISTERS_reg[22][58]  ( .D(n6073), .CK(CLK), .Q(n24672), .QN(n19882) );
  DFF_X1 \REGISTERS_reg[22][57]  ( .D(n6072), .CK(CLK), .Q(n24671), .QN(n19883) );
  DFF_X1 \REGISTERS_reg[22][56]  ( .D(n6071), .CK(CLK), .Q(n24670), .QN(n19884) );
  DFF_X1 \REGISTERS_reg[22][55]  ( .D(n6070), .CK(CLK), .Q(n24669), .QN(n19885) );
  DFF_X1 \REGISTERS_reg[22][54]  ( .D(n6069), .CK(CLK), .Q(n24668), .QN(n19886) );
  DFF_X1 \REGISTERS_reg[22][53]  ( .D(n6068), .CK(CLK), .Q(n24667), .QN(n19887) );
  DFF_X1 \REGISTERS_reg[22][52]  ( .D(n6067), .CK(CLK), .Q(n24666), .QN(n19888) );
  DFF_X1 \REGISTERS_reg[22][51]  ( .D(n6066), .CK(CLK), .Q(n24665), .QN(n19889) );
  DFF_X1 \REGISTERS_reg[22][50]  ( .D(n6065), .CK(CLK), .Q(n24664), .QN(n19890) );
  DFF_X1 \REGISTERS_reg[22][49]  ( .D(n6064), .CK(CLK), .Q(n24663), .QN(n19891) );
  DFF_X1 \REGISTERS_reg[22][48]  ( .D(n6063), .CK(CLK), .Q(n24662), .QN(n19892) );
  DFF_X1 \REGISTERS_reg[22][47]  ( .D(n6062), .CK(CLK), .Q(n24661), .QN(n19893) );
  DFF_X1 \REGISTERS_reg[22][46]  ( .D(n6061), .CK(CLK), .Q(n24660), .QN(n19894) );
  DFF_X1 \REGISTERS_reg[22][45]  ( .D(n6060), .CK(CLK), .Q(n24659), .QN(n19895) );
  DFF_X1 \REGISTERS_reg[22][44]  ( .D(n6059), .CK(CLK), .Q(n24658), .QN(n19896) );
  DFF_X1 \REGISTERS_reg[22][43]  ( .D(n6058), .CK(CLK), .Q(n24657), .QN(n19897) );
  DFF_X1 \REGISTERS_reg[22][42]  ( .D(n6057), .CK(CLK), .Q(n24656), .QN(n19898) );
  DFF_X1 \REGISTERS_reg[22][41]  ( .D(n6056), .CK(CLK), .Q(n24655), .QN(n19899) );
  DFF_X1 \REGISTERS_reg[22][40]  ( .D(n6055), .CK(CLK), .Q(n24654), .QN(n19900) );
  DFF_X1 \REGISTERS_reg[22][39]  ( .D(n6054), .CK(CLK), .Q(n24653), .QN(n19901) );
  DFF_X1 \REGISTERS_reg[22][38]  ( .D(n6053), .CK(CLK), .Q(n24652), .QN(n19902) );
  DFF_X1 \REGISTERS_reg[22][37]  ( .D(n6052), .CK(CLK), .Q(n24651), .QN(n19903) );
  DFF_X1 \REGISTERS_reg[22][36]  ( .D(n6051), .CK(CLK), .Q(n24650), .QN(n19904) );
  DFF_X1 \REGISTERS_reg[22][35]  ( .D(n6050), .CK(CLK), .Q(n24649), .QN(n19905) );
  DFF_X1 \REGISTERS_reg[22][34]  ( .D(n6049), .CK(CLK), .Q(n24648), .QN(n19906) );
  DFF_X1 \REGISTERS_reg[22][33]  ( .D(n6048), .CK(CLK), .Q(n24647), .QN(n19907) );
  DFF_X1 \REGISTERS_reg[22][32]  ( .D(n6047), .CK(CLK), .Q(n24646), .QN(n19908) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n6046), .CK(CLK), .Q(n24645), .QN(n19909) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n6045), .CK(CLK), .Q(n24644), .QN(n19910) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n6044), .CK(CLK), .Q(n24643), .QN(n19911) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n6043), .CK(CLK), .Q(n24642), .QN(n19912) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n6042), .CK(CLK), .Q(n24641), .QN(n19913) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n6041), .CK(CLK), .Q(n24640), .QN(n19914) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n6040), .CK(CLK), .Q(n24639), .QN(n19915) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n6039), .CK(CLK), .Q(n24638), .QN(n19916) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n6038), .CK(CLK), .Q(n24637), .QN(n19917) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n6037), .CK(CLK), .Q(n24636), .QN(n19918) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n6036), .CK(CLK), .Q(n24635), .QN(n19919) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n6035), .CK(CLK), .Q(n24634), .QN(n19920) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n6034), .CK(CLK), .Q(n24633), .QN(n19921) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n6033), .CK(CLK), .Q(n24632), .QN(n19922) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n6032), .CK(CLK), .Q(n24631), .QN(n19923) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n6031), .CK(CLK), .Q(n24630), .QN(n19924) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n6030), .CK(CLK), .Q(n24629), .QN(n19925) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n6029), .CK(CLK), .Q(n24628), .QN(n19926) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n6028), .CK(CLK), .Q(n24627), .QN(n19927) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n6027), .CK(CLK), .Q(n24626), .QN(n19928) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n6026), .CK(CLK), .Q(n24625), .QN(n19929) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n6025), .CK(CLK), .Q(n24624), .QN(n19930) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n6024), .CK(CLK), .Q(n24623), .QN(n19931)
         );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n6023), .CK(CLK), .Q(n24622), .QN(n19932)
         );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n6022), .CK(CLK), .Q(n24621), .QN(n19933)
         );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n6021), .CK(CLK), .Q(n24620), .QN(n19934)
         );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n6020), .CK(CLK), .Q(n24619), .QN(n19935)
         );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n6019), .CK(CLK), .Q(n24618), .QN(n19936)
         );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n6018), .CK(CLK), .Q(n24617), .QN(n19937)
         );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n6017), .CK(CLK), .Q(n24616), .QN(n19938)
         );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n6016), .CK(CLK), .Q(n24615), .QN(n19939)
         );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n6015), .CK(CLK), .Q(n24614), .QN(n19940)
         );
  DFF_X1 \OUT2_reg[63]  ( .D(n5374), .CK(CLK), .Q(OUT2[63]) );
  NOR3_X1 U18481 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(n25046), .ZN(n23931)
         );
  NOR3_X1 U18482 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(n25244), .ZN(n22734)
         );
  NOR3_X1 U18483 ( .A1(n25046), .A2(ADD_RD2[2]), .A3(n19492), .ZN(n23934) );
  NOR3_X1 U18484 ( .A1(n25244), .A2(ADD_RD1[2]), .A3(n19487), .ZN(n22737) );
  BUF_X1 U18485 ( .A(n25570), .Z(n25572) );
  BUF_X1 U18486 ( .A(n25570), .Z(n25573) );
  BUF_X1 U18487 ( .A(n25570), .Z(n25574) );
  BUF_X1 U18488 ( .A(n25571), .Z(n25575) );
  BUF_X1 U18489 ( .A(n25571), .Z(n25576) );
  BUF_X1 U18490 ( .A(n21479), .Z(n25770) );
  BUF_X1 U18491 ( .A(n21479), .Z(n25771) );
  BUF_X1 U18492 ( .A(n21479), .Z(n25772) );
  BUF_X1 U18493 ( .A(n21479), .Z(n25773) );
  BUF_X1 U18494 ( .A(n22798), .Z(n24998) );
  BUF_X1 U18495 ( .A(n22798), .Z(n24999) );
  BUF_X1 U18496 ( .A(n22798), .Z(n25000) );
  BUF_X1 U18497 ( .A(n22798), .Z(n25001) );
  BUF_X1 U18498 ( .A(n22798), .Z(n25002) );
  BUF_X1 U18499 ( .A(n21601), .Z(n25196) );
  BUF_X1 U18500 ( .A(n21601), .Z(n25197) );
  BUF_X1 U18501 ( .A(n21601), .Z(n25198) );
  BUF_X1 U18502 ( .A(n21601), .Z(n25199) );
  BUF_X1 U18503 ( .A(n21601), .Z(n25200) );
  BUF_X1 U18504 ( .A(n25595), .Z(n25597) );
  BUF_X1 U18505 ( .A(n25557), .Z(n25559) );
  BUF_X1 U18506 ( .A(n25467), .Z(n25469) );
  BUF_X1 U18507 ( .A(n25634), .Z(n25636) );
  BUF_X1 U18508 ( .A(n25441), .Z(n25443) );
  BUF_X1 U18509 ( .A(n25402), .Z(n25404) );
  BUF_X1 U18510 ( .A(n25480), .Z(n25482) );
  BUF_X1 U18511 ( .A(n25762), .Z(n25764) );
  BUF_X1 U18512 ( .A(n25454), .Z(n25456) );
  BUF_X1 U18513 ( .A(n25376), .Z(n25378) );
  BUF_X1 U18514 ( .A(n25531), .Z(n25533) );
  BUF_X1 U18515 ( .A(n25724), .Z(n25726) );
  BUF_X1 U18516 ( .A(n25647), .Z(n25649) );
  BUF_X1 U18517 ( .A(n25415), .Z(n25417) );
  BUF_X1 U18518 ( .A(n25389), .Z(n25391) );
  BUF_X1 U18519 ( .A(n25621), .Z(n25623) );
  BUF_X1 U18520 ( .A(n25544), .Z(n25546) );
  BUF_X1 U18521 ( .A(n25518), .Z(n25520) );
  BUF_X1 U18522 ( .A(n25737), .Z(n25739) );
  BUF_X1 U18523 ( .A(n25428), .Z(n25430) );
  BUF_X1 U18524 ( .A(n25493), .Z(n25495) );
  BUF_X1 U18525 ( .A(n25608), .Z(n25610) );
  BUF_X1 U18526 ( .A(n25660), .Z(n25662) );
  BUF_X1 U18527 ( .A(n25673), .Z(n25675) );
  BUF_X1 U18528 ( .A(n25698), .Z(n25700) );
  BUF_X1 U18529 ( .A(n25711), .Z(n25713) );
  BUF_X1 U18530 ( .A(n25595), .Z(n25598) );
  BUF_X1 U18531 ( .A(n25595), .Z(n25599) );
  BUF_X1 U18532 ( .A(n25596), .Z(n25600) );
  BUF_X1 U18533 ( .A(n25596), .Z(n25601) );
  BUF_X1 U18534 ( .A(n25557), .Z(n25560) );
  BUF_X1 U18535 ( .A(n25557), .Z(n25561) );
  BUF_X1 U18536 ( .A(n25558), .Z(n25562) );
  BUF_X1 U18537 ( .A(n25558), .Z(n25563) );
  BUF_X1 U18538 ( .A(n25467), .Z(n25470) );
  BUF_X1 U18539 ( .A(n25467), .Z(n25471) );
  BUF_X1 U18540 ( .A(n25468), .Z(n25472) );
  BUF_X1 U18541 ( .A(n25468), .Z(n25473) );
  BUF_X1 U18542 ( .A(n25634), .Z(n25637) );
  BUF_X1 U18543 ( .A(n25634), .Z(n25638) );
  BUF_X1 U18544 ( .A(n25635), .Z(n25639) );
  BUF_X1 U18545 ( .A(n25635), .Z(n25640) );
  BUF_X1 U18546 ( .A(n25441), .Z(n25444) );
  BUF_X1 U18547 ( .A(n25441), .Z(n25445) );
  BUF_X1 U18548 ( .A(n25442), .Z(n25446) );
  BUF_X1 U18549 ( .A(n25402), .Z(n25405) );
  BUF_X1 U18550 ( .A(n25402), .Z(n25406) );
  BUF_X1 U18551 ( .A(n25403), .Z(n25407) );
  BUF_X1 U18552 ( .A(n25442), .Z(n25447) );
  BUF_X1 U18553 ( .A(n25403), .Z(n25408) );
  BUF_X1 U18554 ( .A(n25480), .Z(n25483) );
  BUF_X1 U18555 ( .A(n25480), .Z(n25484) );
  BUF_X1 U18556 ( .A(n25481), .Z(n25485) );
  BUF_X1 U18557 ( .A(n25481), .Z(n25486) );
  BUF_X1 U18558 ( .A(n25762), .Z(n25765) );
  BUF_X1 U18559 ( .A(n25762), .Z(n25766) );
  BUF_X1 U18560 ( .A(n25763), .Z(n25767) );
  BUF_X1 U18561 ( .A(n25763), .Z(n25768) );
  BUF_X1 U18562 ( .A(n25454), .Z(n25457) );
  BUF_X1 U18563 ( .A(n25454), .Z(n25458) );
  BUF_X1 U18564 ( .A(n25455), .Z(n25459) );
  BUF_X1 U18565 ( .A(n25376), .Z(n25379) );
  BUF_X1 U18566 ( .A(n25376), .Z(n25380) );
  BUF_X1 U18567 ( .A(n25377), .Z(n25381) );
  BUF_X1 U18568 ( .A(n25455), .Z(n25460) );
  BUF_X1 U18569 ( .A(n25377), .Z(n25382) );
  BUF_X1 U18570 ( .A(n25531), .Z(n25534) );
  BUF_X1 U18571 ( .A(n25531), .Z(n25535) );
  BUF_X1 U18572 ( .A(n25532), .Z(n25536) );
  BUF_X1 U18573 ( .A(n25532), .Z(n25537) );
  BUF_X1 U18574 ( .A(n25724), .Z(n25727) );
  BUF_X1 U18575 ( .A(n25724), .Z(n25728) );
  BUF_X1 U18576 ( .A(n25725), .Z(n25729) );
  BUF_X1 U18577 ( .A(n25725), .Z(n25730) );
  BUF_X1 U18578 ( .A(n25647), .Z(n25650) );
  BUF_X1 U18579 ( .A(n25647), .Z(n25651) );
  BUF_X1 U18580 ( .A(n25648), .Z(n25652) );
  BUF_X1 U18581 ( .A(n25648), .Z(n25653) );
  BUF_X1 U18582 ( .A(n25415), .Z(n25418) );
  BUF_X1 U18583 ( .A(n25415), .Z(n25419) );
  BUF_X1 U18584 ( .A(n25416), .Z(n25420) );
  BUF_X1 U18585 ( .A(n25389), .Z(n25392) );
  BUF_X1 U18586 ( .A(n25389), .Z(n25393) );
  BUF_X1 U18587 ( .A(n25390), .Z(n25394) );
  BUF_X1 U18588 ( .A(n25621), .Z(n25624) );
  BUF_X1 U18589 ( .A(n25621), .Z(n25625) );
  BUF_X1 U18590 ( .A(n25622), .Z(n25626) );
  BUF_X1 U18591 ( .A(n25622), .Z(n25627) );
  BUF_X1 U18592 ( .A(n25544), .Z(n25547) );
  BUF_X1 U18593 ( .A(n25544), .Z(n25548) );
  BUF_X1 U18594 ( .A(n25545), .Z(n25549) );
  BUF_X1 U18595 ( .A(n25545), .Z(n25550) );
  BUF_X1 U18596 ( .A(n25518), .Z(n25521) );
  BUF_X1 U18597 ( .A(n25518), .Z(n25522) );
  BUF_X1 U18598 ( .A(n25519), .Z(n25523) );
  BUF_X1 U18599 ( .A(n25519), .Z(n25524) );
  BUF_X1 U18600 ( .A(n25416), .Z(n25421) );
  BUF_X1 U18601 ( .A(n25390), .Z(n25395) );
  BUF_X1 U18602 ( .A(n25737), .Z(n25740) );
  BUF_X1 U18603 ( .A(n25737), .Z(n25741) );
  BUF_X1 U18604 ( .A(n25738), .Z(n25742) );
  BUF_X1 U18605 ( .A(n25738), .Z(n25743) );
  BUF_X1 U18606 ( .A(n25428), .Z(n25431) );
  BUF_X1 U18607 ( .A(n25428), .Z(n25432) );
  BUF_X1 U18608 ( .A(n25429), .Z(n25433) );
  BUF_X1 U18609 ( .A(n25429), .Z(n25434) );
  BUF_X1 U18610 ( .A(n25493), .Z(n25496) );
  BUF_X1 U18611 ( .A(n25493), .Z(n25497) );
  BUF_X1 U18612 ( .A(n25494), .Z(n25498) );
  BUF_X1 U18613 ( .A(n25494), .Z(n25499) );
  BUF_X1 U18614 ( .A(n25608), .Z(n25611) );
  BUF_X1 U18615 ( .A(n25608), .Z(n25612) );
  BUF_X1 U18616 ( .A(n25609), .Z(n25613) );
  BUF_X1 U18617 ( .A(n25609), .Z(n25614) );
  BUF_X1 U18618 ( .A(n25660), .Z(n25663) );
  BUF_X1 U18619 ( .A(n25660), .Z(n25664) );
  BUF_X1 U18620 ( .A(n25661), .Z(n25665) );
  BUF_X1 U18621 ( .A(n25661), .Z(n25666) );
  BUF_X1 U18622 ( .A(n25673), .Z(n25676) );
  BUF_X1 U18623 ( .A(n25673), .Z(n25677) );
  BUF_X1 U18624 ( .A(n25674), .Z(n25678) );
  BUF_X1 U18625 ( .A(n25674), .Z(n25679) );
  BUF_X1 U18626 ( .A(n25698), .Z(n25701) );
  BUF_X1 U18627 ( .A(n25698), .Z(n25702) );
  BUF_X1 U18628 ( .A(n25699), .Z(n25703) );
  BUF_X1 U18629 ( .A(n25699), .Z(n25704) );
  BUF_X1 U18630 ( .A(n25711), .Z(n25714) );
  BUF_X1 U18631 ( .A(n25711), .Z(n25715) );
  BUF_X1 U18632 ( .A(n25712), .Z(n25716) );
  BUF_X1 U18633 ( .A(n25712), .Z(n25717) );
  BUF_X1 U18634 ( .A(n21478), .Z(n25775) );
  BUF_X1 U18635 ( .A(n21478), .Z(n25776) );
  BUF_X1 U18636 ( .A(n21478), .Z(n25777) );
  BUF_X1 U18637 ( .A(n21478), .Z(n25778) );
  BUF_X1 U18638 ( .A(n21478), .Z(n25779) );
  BUF_X1 U18639 ( .A(n21483), .Z(n25756) );
  BUF_X1 U18640 ( .A(n21483), .Z(n25757) );
  BUF_X1 U18641 ( .A(n21483), .Z(n25758) );
  BUF_X1 U18642 ( .A(n21483), .Z(n25759) );
  BUF_X1 U18643 ( .A(n21483), .Z(n25760) );
  BUF_X1 U18644 ( .A(n21555), .Z(n25370) );
  BUF_X1 U18645 ( .A(n21555), .Z(n25371) );
  BUF_X1 U18646 ( .A(n21555), .Z(n25372) );
  BUF_X1 U18647 ( .A(n21555), .Z(n25373) );
  BUF_X1 U18648 ( .A(n21555), .Z(n25374) );
  BUF_X1 U18649 ( .A(n21486), .Z(n25744) );
  BUF_X1 U18650 ( .A(n21486), .Z(n25745) );
  BUF_X1 U18651 ( .A(n21486), .Z(n25746) );
  BUF_X1 U18652 ( .A(n21486), .Z(n25747) );
  BUF_X1 U18653 ( .A(n21486), .Z(n25748) );
  BUF_X1 U18654 ( .A(n21516), .Z(n25589) );
  BUF_X1 U18655 ( .A(n21516), .Z(n25590) );
  BUF_X1 U18656 ( .A(n21516), .Z(n25591) );
  BUF_X1 U18657 ( .A(n21516), .Z(n25592) );
  BUF_X1 U18658 ( .A(n21516), .Z(n25593) );
  BUF_X1 U18659 ( .A(n21523), .Z(n25551) );
  BUF_X1 U18660 ( .A(n21523), .Z(n25552) );
  BUF_X1 U18661 ( .A(n21523), .Z(n25553) );
  BUF_X1 U18662 ( .A(n21523), .Z(n25554) );
  BUF_X1 U18663 ( .A(n21523), .Z(n25555) );
  BUF_X1 U18664 ( .A(n21539), .Z(n25461) );
  BUF_X1 U18665 ( .A(n21539), .Z(n25462) );
  BUF_X1 U18666 ( .A(n21539), .Z(n25463) );
  BUF_X1 U18667 ( .A(n21539), .Z(n25464) );
  BUF_X1 U18668 ( .A(n21539), .Z(n25465) );
  BUF_X1 U18669 ( .A(n21509), .Z(n25628) );
  BUF_X1 U18670 ( .A(n21509), .Z(n25629) );
  BUF_X1 U18671 ( .A(n21509), .Z(n25630) );
  BUF_X1 U18672 ( .A(n21509), .Z(n25631) );
  BUF_X1 U18673 ( .A(n21509), .Z(n25632) );
  BUF_X1 U18674 ( .A(n21544), .Z(n25435) );
  BUF_X1 U18675 ( .A(n21544), .Z(n25436) );
  BUF_X1 U18676 ( .A(n21544), .Z(n25437) );
  BUF_X1 U18677 ( .A(n21544), .Z(n25438) );
  BUF_X1 U18678 ( .A(n21544), .Z(n25439) );
  BUF_X1 U18679 ( .A(n21551), .Z(n25396) );
  BUF_X1 U18680 ( .A(n21551), .Z(n25397) );
  BUF_X1 U18681 ( .A(n21551), .Z(n25398) );
  BUF_X1 U18682 ( .A(n21551), .Z(n25399) );
  BUF_X1 U18683 ( .A(n21551), .Z(n25400) );
  BUF_X1 U18684 ( .A(n21537), .Z(n25474) );
  BUF_X1 U18685 ( .A(n21537), .Z(n25475) );
  BUF_X1 U18686 ( .A(n21537), .Z(n25476) );
  BUF_X1 U18687 ( .A(n21537), .Z(n25477) );
  BUF_X1 U18688 ( .A(n21537), .Z(n25478) );
  BUF_X1 U18689 ( .A(n21520), .Z(n25564) );
  BUF_X1 U18690 ( .A(n21520), .Z(n25565) );
  BUF_X1 U18691 ( .A(n21520), .Z(n25566) );
  BUF_X1 U18692 ( .A(n21520), .Z(n25567) );
  BUF_X1 U18693 ( .A(n21520), .Z(n25568) );
  BUF_X1 U18694 ( .A(n21542), .Z(n25448) );
  BUF_X1 U18695 ( .A(n21542), .Z(n25449) );
  BUF_X1 U18696 ( .A(n21542), .Z(n25450) );
  BUF_X1 U18697 ( .A(n21542), .Z(n25451) );
  BUF_X1 U18698 ( .A(n21542), .Z(n25452) );
  BUF_X1 U18699 ( .A(n21527), .Z(n25525) );
  BUF_X1 U18700 ( .A(n21527), .Z(n25526) );
  BUF_X1 U18701 ( .A(n21527), .Z(n25527) );
  BUF_X1 U18702 ( .A(n21527), .Z(n25528) );
  BUF_X1 U18703 ( .A(n21527), .Z(n25529) );
  BUF_X1 U18704 ( .A(n21493), .Z(n25718) );
  BUF_X1 U18705 ( .A(n21493), .Z(n25719) );
  BUF_X1 U18706 ( .A(n21493), .Z(n25720) );
  BUF_X1 U18707 ( .A(n21493), .Z(n25721) );
  BUF_X1 U18708 ( .A(n21493), .Z(n25722) );
  BUF_X1 U18709 ( .A(n21507), .Z(n25641) );
  BUF_X1 U18710 ( .A(n21507), .Z(n25642) );
  BUF_X1 U18711 ( .A(n21507), .Z(n25643) );
  BUF_X1 U18712 ( .A(n21507), .Z(n25644) );
  BUF_X1 U18713 ( .A(n21507), .Z(n25645) );
  BUF_X1 U18714 ( .A(n21548), .Z(n25409) );
  BUF_X1 U18715 ( .A(n21548), .Z(n25410) );
  BUF_X1 U18716 ( .A(n21548), .Z(n25411) );
  BUF_X1 U18717 ( .A(n21548), .Z(n25412) );
  BUF_X1 U18718 ( .A(n21548), .Z(n25413) );
  BUF_X1 U18719 ( .A(n21553), .Z(n25383) );
  BUF_X1 U18720 ( .A(n21553), .Z(n25384) );
  BUF_X1 U18721 ( .A(n21553), .Z(n25385) );
  BUF_X1 U18722 ( .A(n21553), .Z(n25386) );
  BUF_X1 U18723 ( .A(n21553), .Z(n25387) );
  BUF_X1 U18724 ( .A(n21511), .Z(n25615) );
  BUF_X1 U18725 ( .A(n21511), .Z(n25616) );
  BUF_X1 U18726 ( .A(n21511), .Z(n25617) );
  BUF_X1 U18727 ( .A(n21511), .Z(n25618) );
  BUF_X1 U18728 ( .A(n21511), .Z(n25619) );
  BUF_X1 U18729 ( .A(n21525), .Z(n25538) );
  BUF_X1 U18730 ( .A(n21525), .Z(n25539) );
  BUF_X1 U18731 ( .A(n21525), .Z(n25540) );
  BUF_X1 U18732 ( .A(n21525), .Z(n25541) );
  BUF_X1 U18733 ( .A(n21525), .Z(n25542) );
  BUF_X1 U18734 ( .A(n21530), .Z(n25512) );
  BUF_X1 U18735 ( .A(n21530), .Z(n25513) );
  BUF_X1 U18736 ( .A(n21530), .Z(n25514) );
  BUF_X1 U18737 ( .A(n21530), .Z(n25515) );
  BUF_X1 U18738 ( .A(n21530), .Z(n25516) );
  BUF_X1 U18739 ( .A(n21489), .Z(n25731) );
  BUF_X1 U18740 ( .A(n21489), .Z(n25732) );
  BUF_X1 U18741 ( .A(n21489), .Z(n25733) );
  BUF_X1 U18742 ( .A(n21489), .Z(n25734) );
  BUF_X1 U18743 ( .A(n21489), .Z(n25735) );
  BUF_X1 U18744 ( .A(n21546), .Z(n25422) );
  BUF_X1 U18745 ( .A(n21546), .Z(n25423) );
  BUF_X1 U18746 ( .A(n21546), .Z(n25424) );
  BUF_X1 U18747 ( .A(n21546), .Z(n25425) );
  BUF_X1 U18748 ( .A(n21546), .Z(n25426) );
  BUF_X1 U18749 ( .A(n21518), .Z(n25577) );
  BUF_X1 U18750 ( .A(n21518), .Z(n25578) );
  BUF_X1 U18751 ( .A(n21518), .Z(n25579) );
  BUF_X1 U18752 ( .A(n21518), .Z(n25580) );
  BUF_X1 U18753 ( .A(n21518), .Z(n25581) );
  BUF_X1 U18754 ( .A(n21533), .Z(n25500) );
  BUF_X1 U18755 ( .A(n21533), .Z(n25501) );
  BUF_X1 U18756 ( .A(n21533), .Z(n25502) );
  BUF_X1 U18757 ( .A(n21533), .Z(n25503) );
  BUF_X1 U18758 ( .A(n21533), .Z(n25504) );
  BUF_X1 U18759 ( .A(n21500), .Z(n25680) );
  BUF_X1 U18760 ( .A(n21500), .Z(n25681) );
  BUF_X1 U18761 ( .A(n21500), .Z(n25682) );
  BUF_X1 U18762 ( .A(n21500), .Z(n25683) );
  BUF_X1 U18763 ( .A(n21500), .Z(n25684) );
  BUF_X1 U18764 ( .A(n21535), .Z(n25487) );
  BUF_X1 U18765 ( .A(n21535), .Z(n25488) );
  BUF_X1 U18766 ( .A(n21535), .Z(n25489) );
  BUF_X1 U18767 ( .A(n21535), .Z(n25490) );
  BUF_X1 U18768 ( .A(n21535), .Z(n25491) );
  BUF_X1 U18769 ( .A(n21514), .Z(n25602) );
  BUF_X1 U18770 ( .A(n21514), .Z(n25603) );
  BUF_X1 U18771 ( .A(n21514), .Z(n25604) );
  BUF_X1 U18772 ( .A(n21514), .Z(n25605) );
  BUF_X1 U18773 ( .A(n21514), .Z(n25606) );
  BUF_X1 U18774 ( .A(n21505), .Z(n25654) );
  BUF_X1 U18775 ( .A(n21505), .Z(n25655) );
  BUF_X1 U18776 ( .A(n21505), .Z(n25656) );
  BUF_X1 U18777 ( .A(n21505), .Z(n25657) );
  BUF_X1 U18778 ( .A(n21505), .Z(n25658) );
  BUF_X1 U18779 ( .A(n21502), .Z(n25667) );
  BUF_X1 U18780 ( .A(n21502), .Z(n25668) );
  BUF_X1 U18781 ( .A(n21502), .Z(n25669) );
  BUF_X1 U18782 ( .A(n21502), .Z(n25670) );
  BUF_X1 U18783 ( .A(n21502), .Z(n25671) );
  BUF_X1 U18784 ( .A(n21498), .Z(n25692) );
  BUF_X1 U18785 ( .A(n21498), .Z(n25693) );
  BUF_X1 U18786 ( .A(n21498), .Z(n25694) );
  BUF_X1 U18787 ( .A(n21498), .Z(n25695) );
  BUF_X1 U18788 ( .A(n21498), .Z(n25696) );
  BUF_X1 U18789 ( .A(n21496), .Z(n25705) );
  BUF_X1 U18790 ( .A(n21496), .Z(n25706) );
  BUF_X1 U18791 ( .A(n21496), .Z(n25707) );
  BUF_X1 U18792 ( .A(n21496), .Z(n25708) );
  BUF_X1 U18793 ( .A(n21496), .Z(n25709) );
  BUF_X1 U18794 ( .A(n21479), .Z(n25769) );
  BUF_X1 U18795 ( .A(n21519), .Z(n25570) );
  BUF_X1 U18796 ( .A(n21519), .Z(n25571) );
  OAI21_X1 U18797 ( .B1(n21480), .B2(n21481), .A(n25973), .ZN(n21478) );
  BUF_X1 U18798 ( .A(n22777), .Z(n25082) );
  BUF_X1 U18799 ( .A(n22777), .Z(n25083) );
  BUF_X1 U18800 ( .A(n22777), .Z(n25084) );
  BUF_X1 U18801 ( .A(n22777), .Z(n25085) );
  BUF_X1 U18802 ( .A(n22777), .Z(n25086) );
  BUF_X1 U18803 ( .A(n21580), .Z(n25280) );
  BUF_X1 U18804 ( .A(n21580), .Z(n25281) );
  BUF_X1 U18805 ( .A(n21580), .Z(n25282) );
  BUF_X1 U18806 ( .A(n21580), .Z(n25283) );
  BUF_X1 U18807 ( .A(n21580), .Z(n25284) );
  BUF_X1 U18808 ( .A(n22787), .Z(n25052) );
  BUF_X1 U18809 ( .A(n22787), .Z(n25053) );
  BUF_X1 U18810 ( .A(n22787), .Z(n25054) );
  BUF_X1 U18811 ( .A(n22787), .Z(n25055) );
  BUF_X1 U18812 ( .A(n22787), .Z(n25056) );
  BUF_X1 U18813 ( .A(n21590), .Z(n25250) );
  BUF_X1 U18814 ( .A(n21590), .Z(n25251) );
  BUF_X1 U18815 ( .A(n21590), .Z(n25252) );
  BUF_X1 U18816 ( .A(n21590), .Z(n25253) );
  BUF_X1 U18817 ( .A(n21590), .Z(n25254) );
  BUF_X1 U18818 ( .A(n22767), .Z(n25130) );
  BUF_X1 U18819 ( .A(n22767), .Z(n25131) );
  BUF_X1 U18820 ( .A(n22767), .Z(n25132) );
  BUF_X1 U18821 ( .A(n22767), .Z(n25133) );
  BUF_X1 U18822 ( .A(n22767), .Z(n25134) );
  BUF_X1 U18823 ( .A(n21570), .Z(n25328) );
  BUF_X1 U18824 ( .A(n21570), .Z(n25329) );
  BUF_X1 U18825 ( .A(n21570), .Z(n25330) );
  BUF_X1 U18826 ( .A(n21570), .Z(n25331) );
  BUF_X1 U18827 ( .A(n21570), .Z(n25332) );
  BUF_X1 U18828 ( .A(n22762), .Z(n25154) );
  BUF_X1 U18829 ( .A(n22772), .Z(n25106) );
  BUF_X1 U18830 ( .A(n22792), .Z(n25028) );
  BUF_X1 U18831 ( .A(n22797), .Z(n25004) );
  BUF_X1 U18832 ( .A(n22802), .Z(n24980) );
  BUF_X1 U18833 ( .A(n22762), .Z(n25155) );
  BUF_X1 U18834 ( .A(n22772), .Z(n25107) );
  BUF_X1 U18835 ( .A(n22792), .Z(n25029) );
  BUF_X1 U18836 ( .A(n22797), .Z(n25005) );
  BUF_X1 U18837 ( .A(n22802), .Z(n24981) );
  BUF_X1 U18838 ( .A(n22762), .Z(n25156) );
  BUF_X1 U18839 ( .A(n22772), .Z(n25108) );
  BUF_X1 U18840 ( .A(n22792), .Z(n25030) );
  BUF_X1 U18841 ( .A(n22797), .Z(n25006) );
  BUF_X1 U18842 ( .A(n22802), .Z(n24982) );
  BUF_X1 U18843 ( .A(n22762), .Z(n25157) );
  BUF_X1 U18844 ( .A(n22772), .Z(n25109) );
  BUF_X1 U18845 ( .A(n22792), .Z(n25031) );
  BUF_X1 U18846 ( .A(n22797), .Z(n25007) );
  BUF_X1 U18847 ( .A(n22802), .Z(n24983) );
  BUF_X1 U18848 ( .A(n22762), .Z(n25158) );
  BUF_X1 U18849 ( .A(n22772), .Z(n25110) );
  BUF_X1 U18850 ( .A(n22792), .Z(n25032) );
  BUF_X1 U18851 ( .A(n22797), .Z(n25008) );
  BUF_X1 U18852 ( .A(n22802), .Z(n24984) );
  BUF_X1 U18853 ( .A(n21565), .Z(n25352) );
  BUF_X1 U18854 ( .A(n21575), .Z(n25304) );
  BUF_X1 U18855 ( .A(n21595), .Z(n25226) );
  BUF_X1 U18856 ( .A(n21600), .Z(n25202) );
  BUF_X1 U18857 ( .A(n21605), .Z(n25178) );
  BUF_X1 U18858 ( .A(n21565), .Z(n25353) );
  BUF_X1 U18859 ( .A(n21575), .Z(n25305) );
  BUF_X1 U18860 ( .A(n21595), .Z(n25227) );
  BUF_X1 U18861 ( .A(n21600), .Z(n25203) );
  BUF_X1 U18862 ( .A(n21605), .Z(n25179) );
  BUF_X1 U18863 ( .A(n21565), .Z(n25354) );
  BUF_X1 U18864 ( .A(n21575), .Z(n25306) );
  BUF_X1 U18865 ( .A(n21595), .Z(n25228) );
  BUF_X1 U18866 ( .A(n21600), .Z(n25204) );
  BUF_X1 U18867 ( .A(n21605), .Z(n25180) );
  BUF_X1 U18868 ( .A(n21565), .Z(n25355) );
  BUF_X1 U18869 ( .A(n21575), .Z(n25307) );
  BUF_X1 U18870 ( .A(n21595), .Z(n25229) );
  BUF_X1 U18871 ( .A(n21600), .Z(n25205) );
  BUF_X1 U18872 ( .A(n21605), .Z(n25181) );
  BUF_X1 U18873 ( .A(n21565), .Z(n25356) );
  BUF_X1 U18874 ( .A(n21575), .Z(n25308) );
  BUF_X1 U18875 ( .A(n21595), .Z(n25230) );
  BUF_X1 U18876 ( .A(n21600), .Z(n25206) );
  BUF_X1 U18877 ( .A(n21605), .Z(n25182) );
  BUF_X1 U18878 ( .A(n22759), .Z(n25167) );
  BUF_X1 U18879 ( .A(n22769), .Z(n25119) );
  BUF_X1 U18880 ( .A(n22764), .Z(n25143) );
  BUF_X1 U18881 ( .A(n22789), .Z(n25041) );
  BUF_X1 U18882 ( .A(n22759), .Z(n25168) );
  BUF_X1 U18883 ( .A(n22769), .Z(n25120) );
  BUF_X1 U18884 ( .A(n22764), .Z(n25144) );
  BUF_X1 U18885 ( .A(n22789), .Z(n25042) );
  BUF_X1 U18886 ( .A(n22759), .Z(n25169) );
  BUF_X1 U18887 ( .A(n22769), .Z(n25121) );
  BUF_X1 U18888 ( .A(n22764), .Z(n25145) );
  BUF_X1 U18889 ( .A(n22789), .Z(n25043) );
  BUF_X1 U18890 ( .A(n22759), .Z(n25170) );
  BUF_X1 U18891 ( .A(n22769), .Z(n25122) );
  BUF_X1 U18892 ( .A(n22764), .Z(n25146) );
  BUF_X1 U18893 ( .A(n22789), .Z(n25044) );
  BUF_X1 U18894 ( .A(n21562), .Z(n25365) );
  BUF_X1 U18895 ( .A(n21572), .Z(n25317) );
  BUF_X1 U18896 ( .A(n21567), .Z(n25341) );
  BUF_X1 U18897 ( .A(n21592), .Z(n25239) );
  BUF_X1 U18898 ( .A(n21562), .Z(n25366) );
  BUF_X1 U18899 ( .A(n21572), .Z(n25318) );
  BUF_X1 U18900 ( .A(n21567), .Z(n25342) );
  BUF_X1 U18901 ( .A(n21592), .Z(n25240) );
  BUF_X1 U18902 ( .A(n21562), .Z(n25367) );
  BUF_X1 U18903 ( .A(n21572), .Z(n25319) );
  BUF_X1 U18904 ( .A(n21567), .Z(n25343) );
  BUF_X1 U18905 ( .A(n21592), .Z(n25241) );
  BUF_X1 U18906 ( .A(n21562), .Z(n25368) );
  BUF_X1 U18907 ( .A(n21572), .Z(n25320) );
  BUF_X1 U18908 ( .A(n21567), .Z(n25344) );
  BUF_X1 U18909 ( .A(n21592), .Z(n25242) );
  BUF_X1 U18910 ( .A(n22774), .Z(n25095) );
  BUF_X1 U18911 ( .A(n22794), .Z(n25017) );
  BUF_X1 U18912 ( .A(n22774), .Z(n25096) );
  BUF_X1 U18913 ( .A(n22774), .Z(n25097) );
  BUF_X1 U18914 ( .A(n22799), .Z(n24993) );
  BUF_X1 U18915 ( .A(n22794), .Z(n25018) );
  BUF_X1 U18916 ( .A(n22794), .Z(n25019) );
  BUF_X1 U18917 ( .A(n22774), .Z(n25098) );
  BUF_X1 U18918 ( .A(n22794), .Z(n25020) );
  BUF_X1 U18919 ( .A(n21577), .Z(n25293) );
  BUF_X1 U18920 ( .A(n21577), .Z(n25294) );
  BUF_X1 U18921 ( .A(n21577), .Z(n25296) );
  BUF_X1 U18922 ( .A(n22784), .Z(n25065) );
  BUF_X1 U18923 ( .A(n22784), .Z(n25066) );
  BUF_X1 U18924 ( .A(n22799), .Z(n24994) );
  BUF_X1 U18925 ( .A(n22784), .Z(n25067) );
  BUF_X1 U18926 ( .A(n22799), .Z(n24995) );
  BUF_X1 U18927 ( .A(n22784), .Z(n25068) );
  BUF_X1 U18928 ( .A(n22799), .Z(n24996) );
  BUF_X1 U18929 ( .A(n21587), .Z(n25263) );
  BUF_X1 U18930 ( .A(n21597), .Z(n25215) );
  BUF_X1 U18931 ( .A(n21577), .Z(n25295) );
  BUF_X1 U18932 ( .A(n21602), .Z(n25191) );
  BUF_X1 U18933 ( .A(n21587), .Z(n25264) );
  BUF_X1 U18934 ( .A(n21597), .Z(n25216) );
  BUF_X1 U18935 ( .A(n21602), .Z(n25192) );
  BUF_X1 U18936 ( .A(n21587), .Z(n25265) );
  BUF_X1 U18937 ( .A(n21597), .Z(n25217) );
  BUF_X1 U18938 ( .A(n21602), .Z(n25193) );
  BUF_X1 U18939 ( .A(n21587), .Z(n25266) );
  BUF_X1 U18940 ( .A(n21597), .Z(n25218) );
  BUF_X1 U18941 ( .A(n21602), .Z(n25194) );
  BUF_X1 U18942 ( .A(n22778), .Z(n25076) );
  BUF_X1 U18943 ( .A(n22778), .Z(n25077) );
  BUF_X1 U18944 ( .A(n22778), .Z(n25078) );
  BUF_X1 U18945 ( .A(n22778), .Z(n25079) );
  BUF_X1 U18946 ( .A(n22778), .Z(n25080) );
  BUF_X1 U18947 ( .A(n21581), .Z(n25274) );
  BUF_X1 U18948 ( .A(n21581), .Z(n25275) );
  BUF_X1 U18949 ( .A(n21581), .Z(n25276) );
  BUF_X1 U18950 ( .A(n21581), .Z(n25277) );
  BUF_X1 U18951 ( .A(n21581), .Z(n25278) );
  BUF_X1 U18952 ( .A(n22773), .Z(n25100) );
  BUF_X1 U18953 ( .A(n22768), .Z(n25124) );
  BUF_X1 U18954 ( .A(n22793), .Z(n25022) );
  BUF_X1 U18955 ( .A(n22803), .Z(n24974) );
  BUF_X1 U18956 ( .A(n22773), .Z(n25101) );
  BUF_X1 U18957 ( .A(n22768), .Z(n25125) );
  BUF_X1 U18958 ( .A(n22793), .Z(n25023) );
  BUF_X1 U18959 ( .A(n22803), .Z(n24975) );
  BUF_X1 U18960 ( .A(n22773), .Z(n25102) );
  BUF_X1 U18961 ( .A(n22768), .Z(n25126) );
  BUF_X1 U18962 ( .A(n22793), .Z(n25024) );
  BUF_X1 U18963 ( .A(n22803), .Z(n24976) );
  BUF_X1 U18964 ( .A(n22773), .Z(n25103) );
  BUF_X1 U18965 ( .A(n22768), .Z(n25127) );
  BUF_X1 U18966 ( .A(n22793), .Z(n25025) );
  BUF_X1 U18967 ( .A(n22803), .Z(n24977) );
  BUF_X1 U18968 ( .A(n22773), .Z(n25104) );
  BUF_X1 U18969 ( .A(n22768), .Z(n25128) );
  BUF_X1 U18970 ( .A(n22793), .Z(n25026) );
  BUF_X1 U18971 ( .A(n22803), .Z(n24978) );
  BUF_X1 U18972 ( .A(n21576), .Z(n25298) );
  BUF_X1 U18973 ( .A(n21571), .Z(n25322) );
  BUF_X1 U18974 ( .A(n21596), .Z(n25220) );
  BUF_X1 U18975 ( .A(n21606), .Z(n25172) );
  BUF_X1 U18976 ( .A(n21576), .Z(n25299) );
  BUF_X1 U18977 ( .A(n21571), .Z(n25323) );
  BUF_X1 U18978 ( .A(n21596), .Z(n25221) );
  BUF_X1 U18979 ( .A(n21606), .Z(n25173) );
  BUF_X1 U18980 ( .A(n21576), .Z(n25300) );
  BUF_X1 U18981 ( .A(n21571), .Z(n25324) );
  BUF_X1 U18982 ( .A(n21596), .Z(n25222) );
  BUF_X1 U18983 ( .A(n21606), .Z(n25174) );
  BUF_X1 U18984 ( .A(n21576), .Z(n25301) );
  BUF_X1 U18985 ( .A(n21571), .Z(n25325) );
  BUF_X1 U18986 ( .A(n21596), .Z(n25223) );
  BUF_X1 U18987 ( .A(n21606), .Z(n25175) );
  BUF_X1 U18988 ( .A(n21576), .Z(n25302) );
  BUF_X1 U18989 ( .A(n21571), .Z(n25326) );
  BUF_X1 U18990 ( .A(n21596), .Z(n25224) );
  BUF_X1 U18991 ( .A(n21606), .Z(n25176) );
  BUF_X1 U18992 ( .A(n22763), .Z(n25148) );
  BUF_X1 U18993 ( .A(n22763), .Z(n25149) );
  BUF_X1 U18994 ( .A(n22763), .Z(n25150) );
  BUF_X1 U18995 ( .A(n22763), .Z(n25151) );
  BUF_X1 U18996 ( .A(n22763), .Z(n25152) );
  BUF_X1 U18997 ( .A(n21566), .Z(n25346) );
  BUF_X1 U18998 ( .A(n21566), .Z(n25347) );
  BUF_X1 U18999 ( .A(n21566), .Z(n25348) );
  BUF_X1 U19000 ( .A(n21566), .Z(n25349) );
  BUF_X1 U19001 ( .A(n21566), .Z(n25350) );
  BUF_X1 U19002 ( .A(n22779), .Z(n25070) );
  BUF_X1 U19003 ( .A(n22779), .Z(n25071) );
  BUF_X1 U19004 ( .A(n22779), .Z(n25072) );
  BUF_X1 U19005 ( .A(n22779), .Z(n25073) );
  BUF_X1 U19006 ( .A(n22779), .Z(n25074) );
  BUF_X1 U19007 ( .A(n21582), .Z(n25268) );
  BUF_X1 U19008 ( .A(n21582), .Z(n25269) );
  BUF_X1 U19009 ( .A(n21582), .Z(n25270) );
  BUF_X1 U19010 ( .A(n21582), .Z(n25271) );
  BUF_X1 U19011 ( .A(n21582), .Z(n25272) );
  NAND2_X1 U19012 ( .A1(n25978), .A2(n25764), .ZN(n21483) );
  NAND2_X1 U19013 ( .A1(n25978), .A2(n25378), .ZN(n21555) );
  NAND2_X1 U19014 ( .A1(n25978), .A2(n25750), .ZN(n21486) );
  BUF_X1 U19015 ( .A(n21517), .Z(n25583) );
  BUF_X1 U19016 ( .A(n21532), .Z(n25506) );
  BUF_X1 U19017 ( .A(n21485), .Z(n25750) );
  BUF_X1 U19018 ( .A(n21499), .Z(n25686) );
  BUF_X1 U19019 ( .A(n21517), .Z(n25584) );
  BUF_X1 U19020 ( .A(n21517), .Z(n25585) );
  BUF_X1 U19021 ( .A(n21517), .Z(n25586) );
  BUF_X1 U19022 ( .A(n21517), .Z(n25587) );
  BUF_X1 U19023 ( .A(n21532), .Z(n25507) );
  BUF_X1 U19024 ( .A(n21532), .Z(n25508) );
  BUF_X1 U19025 ( .A(n21532), .Z(n25509) );
  BUF_X1 U19026 ( .A(n21532), .Z(n25510) );
  BUF_X1 U19027 ( .A(n21485), .Z(n25751) );
  BUF_X1 U19028 ( .A(n21485), .Z(n25752) );
  BUF_X1 U19029 ( .A(n21485), .Z(n25753) );
  BUF_X1 U19030 ( .A(n21485), .Z(n25754) );
  BUF_X1 U19031 ( .A(n21499), .Z(n25687) );
  BUF_X1 U19032 ( .A(n21499), .Z(n25688) );
  BUF_X1 U19033 ( .A(n21499), .Z(n25689) );
  BUF_X1 U19034 ( .A(n21499), .Z(n25690) );
  NAND2_X1 U19035 ( .A1(n25975), .A2(n25546), .ZN(n21525) );
  NAND2_X1 U19036 ( .A1(n25975), .A2(n25520), .ZN(n21530) );
  NAND2_X1 U19037 ( .A1(n25975), .A2(n25506), .ZN(n21533) );
  NAND2_X1 U19038 ( .A1(n25975), .A2(n25495), .ZN(n21535) );
  NAND2_X1 U19039 ( .A1(n25976), .A2(n25597), .ZN(n21516) );
  NAND2_X1 U19040 ( .A1(n25976), .A2(n25559), .ZN(n21523) );
  NAND2_X1 U19041 ( .A1(n25976), .A2(n25469), .ZN(n21539) );
  NAND2_X1 U19042 ( .A1(n25976), .A2(n25636), .ZN(n21509) );
  NAND2_X1 U19043 ( .A1(n25976), .A2(n25443), .ZN(n21544) );
  NAND2_X1 U19044 ( .A1(n25977), .A2(n25404), .ZN(n21551) );
  NAND2_X1 U19045 ( .A1(n25976), .A2(n25482), .ZN(n21537) );
  NAND2_X1 U19046 ( .A1(n25976), .A2(n25572), .ZN(n21520) );
  NAND2_X1 U19047 ( .A1(n25977), .A2(n25456), .ZN(n21542) );
  NAND2_X1 U19048 ( .A1(n25976), .A2(n25533), .ZN(n21527) );
  NAND2_X1 U19049 ( .A1(n25977), .A2(n25726), .ZN(n21493) );
  NAND2_X1 U19050 ( .A1(n25976), .A2(n25649), .ZN(n21507) );
  NAND2_X1 U19051 ( .A1(n25976), .A2(n25623), .ZN(n21511) );
  NAND2_X1 U19052 ( .A1(n25977), .A2(n25417), .ZN(n21548) );
  NAND2_X1 U19053 ( .A1(n25977), .A2(n25391), .ZN(n21553) );
  NAND2_X1 U19054 ( .A1(n25977), .A2(n25739), .ZN(n21489) );
  NAND2_X1 U19055 ( .A1(n25977), .A2(n25430), .ZN(n21546) );
  NAND2_X1 U19056 ( .A1(n25976), .A2(n25583), .ZN(n21518) );
  NAND2_X1 U19057 ( .A1(n25977), .A2(n25686), .ZN(n21500) );
  NAND2_X1 U19058 ( .A1(n25976), .A2(n25610), .ZN(n21514) );
  NAND2_X1 U19059 ( .A1(n25977), .A2(n25662), .ZN(n21505) );
  NAND2_X1 U19060 ( .A1(n25977), .A2(n25675), .ZN(n21502) );
  NAND2_X1 U19061 ( .A1(n25977), .A2(n25700), .ZN(n21498) );
  NAND2_X1 U19062 ( .A1(n25977), .A2(n25713), .ZN(n21496) );
  BUF_X1 U19063 ( .A(n22775), .Z(n25088) );
  BUF_X1 U19064 ( .A(n22760), .Z(n25160) );
  BUF_X1 U19065 ( .A(n22765), .Z(n25136) );
  BUF_X1 U19066 ( .A(n22795), .Z(n25010) );
  BUF_X1 U19067 ( .A(n22775), .Z(n25089) );
  BUF_X1 U19068 ( .A(n22760), .Z(n25161) );
  BUF_X1 U19069 ( .A(n22765), .Z(n25137) );
  BUF_X1 U19070 ( .A(n22795), .Z(n25011) );
  BUF_X1 U19071 ( .A(n22760), .Z(n25162) );
  BUF_X1 U19072 ( .A(n22795), .Z(n25012) );
  BUF_X1 U19073 ( .A(n22785), .Z(n25059) );
  BUF_X1 U19074 ( .A(n22775), .Z(n25090) );
  BUF_X1 U19075 ( .A(n22765), .Z(n25138) );
  BUF_X1 U19076 ( .A(n22775), .Z(n25091) );
  BUF_X1 U19077 ( .A(n22760), .Z(n25163) );
  BUF_X1 U19078 ( .A(n22765), .Z(n25139) );
  BUF_X1 U19079 ( .A(n22795), .Z(n25013) );
  BUF_X1 U19080 ( .A(n22765), .Z(n25140) );
  BUF_X1 U19081 ( .A(n22795), .Z(n25014) );
  BUF_X1 U19082 ( .A(n21578), .Z(n25286) );
  BUF_X1 U19083 ( .A(n21563), .Z(n25358) );
  BUF_X1 U19084 ( .A(n21568), .Z(n25334) );
  BUF_X1 U19085 ( .A(n21598), .Z(n25208) );
  BUF_X1 U19086 ( .A(n21563), .Z(n25359) );
  BUF_X1 U19087 ( .A(n21568), .Z(n25335) );
  BUF_X1 U19088 ( .A(n21598), .Z(n25209) );
  BUF_X1 U19089 ( .A(n21563), .Z(n25360) );
  BUF_X1 U19090 ( .A(n21568), .Z(n25336) );
  BUF_X1 U19091 ( .A(n21598), .Z(n25210) );
  BUF_X1 U19092 ( .A(n21563), .Z(n25361) );
  BUF_X1 U19093 ( .A(n21598), .Z(n25211) );
  BUF_X1 U19094 ( .A(n21563), .Z(n25362) );
  BUF_X1 U19095 ( .A(n21568), .Z(n25338) );
  BUF_X1 U19096 ( .A(n21598), .Z(n25212) );
  BUF_X1 U19097 ( .A(n22790), .Z(n25034) );
  BUF_X1 U19098 ( .A(n22785), .Z(n25058) );
  BUF_X1 U19099 ( .A(n22790), .Z(n25035) );
  BUF_X1 U19100 ( .A(n22785), .Z(n25060) );
  BUF_X1 U19101 ( .A(n22790), .Z(n25037) );
  BUF_X1 U19102 ( .A(n22785), .Z(n25061) );
  BUF_X1 U19103 ( .A(n22775), .Z(n25092) );
  BUF_X1 U19104 ( .A(n22760), .Z(n25164) );
  BUF_X1 U19105 ( .A(n22790), .Z(n25038) );
  BUF_X1 U19106 ( .A(n22785), .Z(n25062) );
  BUF_X1 U19107 ( .A(n21593), .Z(n25232) );
  BUF_X1 U19108 ( .A(n21588), .Z(n25256) );
  BUF_X1 U19109 ( .A(n21578), .Z(n25287) );
  BUF_X1 U19110 ( .A(n21568), .Z(n25337) );
  BUF_X1 U19111 ( .A(n22790), .Z(n25036) );
  BUF_X1 U19112 ( .A(n21593), .Z(n25233) );
  BUF_X1 U19113 ( .A(n21588), .Z(n25257) );
  BUF_X1 U19114 ( .A(n21578), .Z(n25288) );
  BUF_X1 U19115 ( .A(n21593), .Z(n25234) );
  BUF_X1 U19116 ( .A(n21588), .Z(n25258) );
  BUF_X1 U19117 ( .A(n21578), .Z(n25289) );
  BUF_X1 U19118 ( .A(n21593), .Z(n25235) );
  BUF_X1 U19119 ( .A(n21588), .Z(n25259) );
  BUF_X1 U19120 ( .A(n21578), .Z(n25290) );
  BUF_X1 U19121 ( .A(n21593), .Z(n25236) );
  BUF_X1 U19122 ( .A(n21588), .Z(n25260) );
  BUF_X1 U19123 ( .A(n22770), .Z(n25112) );
  BUF_X1 U19124 ( .A(n22800), .Z(n24986) );
  BUF_X1 U19125 ( .A(n22770), .Z(n25113) );
  BUF_X1 U19126 ( .A(n22800), .Z(n24987) );
  BUF_X1 U19127 ( .A(n22770), .Z(n25114) );
  BUF_X1 U19128 ( .A(n22800), .Z(n24988) );
  BUF_X1 U19129 ( .A(n22770), .Z(n25115) );
  BUF_X1 U19130 ( .A(n22800), .Z(n24989) );
  BUF_X1 U19131 ( .A(n22770), .Z(n25116) );
  BUF_X1 U19132 ( .A(n22800), .Z(n24990) );
  BUF_X1 U19133 ( .A(n21573), .Z(n25310) );
  BUF_X1 U19134 ( .A(n21603), .Z(n25184) );
  BUF_X1 U19135 ( .A(n21573), .Z(n25311) );
  BUF_X1 U19136 ( .A(n21603), .Z(n25185) );
  BUF_X1 U19137 ( .A(n21573), .Z(n25312) );
  BUF_X1 U19138 ( .A(n21603), .Z(n25186) );
  BUF_X1 U19139 ( .A(n21573), .Z(n25313) );
  BUF_X1 U19140 ( .A(n21603), .Z(n25187) );
  BUF_X1 U19141 ( .A(n21573), .Z(n25314) );
  BUF_X1 U19142 ( .A(n21603), .Z(n25188) );
  BUF_X1 U19143 ( .A(n22759), .Z(n25166) );
  BUF_X1 U19144 ( .A(n22764), .Z(n25142) );
  BUF_X1 U19145 ( .A(n22789), .Z(n25040) );
  BUF_X1 U19146 ( .A(n21562), .Z(n25364) );
  BUF_X1 U19147 ( .A(n21567), .Z(n25340) );
  BUF_X1 U19148 ( .A(n21592), .Z(n25238) );
  BUF_X1 U19149 ( .A(n22769), .Z(n25118) );
  BUF_X1 U19150 ( .A(n21572), .Z(n25316) );
  BUF_X1 U19151 ( .A(n22774), .Z(n25094) );
  BUF_X1 U19152 ( .A(n22794), .Z(n25016) );
  BUF_X1 U19153 ( .A(n21577), .Z(n25292) );
  BUF_X1 U19154 ( .A(n21597), .Z(n25214) );
  BUF_X1 U19155 ( .A(n22784), .Z(n25064) );
  BUF_X1 U19156 ( .A(n22799), .Z(n24992) );
  BUF_X1 U19157 ( .A(n21587), .Z(n25262) );
  BUF_X1 U19158 ( .A(n21602), .Z(n25190) );
  NAND2_X1 U19159 ( .A1(n25978), .A2(n25775), .ZN(n21479) );
  OAI21_X1 U19160 ( .B1(n21481), .B2(n21521), .A(n25974), .ZN(n21519) );
  AND2_X1 U19161 ( .A1(n23946), .A2(n23928), .ZN(n22798) );
  AND2_X1 U19162 ( .A1(n22749), .A2(n22731), .ZN(n21601) );
  BUF_X1 U19163 ( .A(n21482), .Z(n25762) );
  BUF_X1 U19164 ( .A(n21488), .Z(n25737) );
  BUF_X1 U19165 ( .A(n21515), .Z(n25595) );
  BUF_X1 U19166 ( .A(n21522), .Z(n25557) );
  BUF_X1 U19167 ( .A(n21538), .Z(n25467) );
  BUF_X1 U19168 ( .A(n21508), .Z(n25634) );
  BUF_X1 U19169 ( .A(n21543), .Z(n25441) );
  BUF_X1 U19170 ( .A(n21550), .Z(n25402) );
  BUF_X1 U19171 ( .A(n21536), .Z(n25480) );
  BUF_X1 U19172 ( .A(n21541), .Z(n25454) );
  BUF_X1 U19173 ( .A(n21554), .Z(n25376) );
  BUF_X1 U19174 ( .A(n21526), .Z(n25531) );
  BUF_X1 U19175 ( .A(n21492), .Z(n25724) );
  BUF_X1 U19176 ( .A(n21506), .Z(n25647) );
  BUF_X1 U19177 ( .A(n21547), .Z(n25415) );
  BUF_X1 U19178 ( .A(n21552), .Z(n25389) );
  BUF_X1 U19179 ( .A(n21510), .Z(n25621) );
  BUF_X1 U19180 ( .A(n21524), .Z(n25544) );
  BUF_X1 U19181 ( .A(n21529), .Z(n25518) );
  BUF_X1 U19182 ( .A(n21545), .Z(n25428) );
  BUF_X1 U19183 ( .A(n21534), .Z(n25493) );
  BUF_X1 U19184 ( .A(n21513), .Z(n25608) );
  BUF_X1 U19185 ( .A(n21504), .Z(n25660) );
  BUF_X1 U19186 ( .A(n21501), .Z(n25673) );
  BUF_X1 U19187 ( .A(n21497), .Z(n25698) );
  BUF_X1 U19188 ( .A(n21495), .Z(n25711) );
  BUF_X1 U19189 ( .A(n21482), .Z(n25763) );
  BUF_X1 U19190 ( .A(n21488), .Z(n25738) );
  BUF_X1 U19191 ( .A(n21515), .Z(n25596) );
  BUF_X1 U19192 ( .A(n21522), .Z(n25558) );
  BUF_X1 U19193 ( .A(n21538), .Z(n25468) );
  BUF_X1 U19194 ( .A(n21508), .Z(n25635) );
  BUF_X1 U19195 ( .A(n21543), .Z(n25442) );
  BUF_X1 U19196 ( .A(n21550), .Z(n25403) );
  BUF_X1 U19197 ( .A(n21536), .Z(n25481) );
  BUF_X1 U19198 ( .A(n21541), .Z(n25455) );
  BUF_X1 U19199 ( .A(n21554), .Z(n25377) );
  BUF_X1 U19200 ( .A(n21526), .Z(n25532) );
  BUF_X1 U19201 ( .A(n21492), .Z(n25725) );
  BUF_X1 U19202 ( .A(n21506), .Z(n25648) );
  BUF_X1 U19203 ( .A(n21510), .Z(n25622) );
  BUF_X1 U19204 ( .A(n21524), .Z(n25545) );
  BUF_X1 U19205 ( .A(n21529), .Z(n25519) );
  BUF_X1 U19206 ( .A(n21547), .Z(n25416) );
  BUF_X1 U19207 ( .A(n21552), .Z(n25390) );
  BUF_X1 U19208 ( .A(n21545), .Z(n25429) );
  BUF_X1 U19209 ( .A(n21534), .Z(n25494) );
  BUF_X1 U19210 ( .A(n21513), .Z(n25609) );
  BUF_X1 U19211 ( .A(n21504), .Z(n25661) );
  BUF_X1 U19212 ( .A(n21501), .Z(n25674) );
  BUF_X1 U19213 ( .A(n21497), .Z(n25699) );
  BUF_X1 U19214 ( .A(n21495), .Z(n25712) );
  OAI22_X1 U19215 ( .A1(n25563), .A2(n21353), .B1(n25962), .B2(n25556), .ZN(
        n6395) );
  OAI22_X1 U19216 ( .A1(n25563), .A2(n21352), .B1(n25965), .B2(n25556), .ZN(
        n6396) );
  OAI22_X1 U19217 ( .A1(n25563), .A2(n21351), .B1(n25968), .B2(n25556), .ZN(
        n6397) );
  OAI22_X1 U19218 ( .A1(n25563), .A2(n21350), .B1(n25971), .B2(n25556), .ZN(
        n6398) );
  OAI22_X1 U19219 ( .A1(n25640), .A2(n21225), .B1(n25961), .B2(n25633), .ZN(
        n6779) );
  OAI22_X1 U19220 ( .A1(n25640), .A2(n21224), .B1(n25964), .B2(n25633), .ZN(
        n6780) );
  OAI22_X1 U19221 ( .A1(n25640), .A2(n21223), .B1(n25967), .B2(n25633), .ZN(
        n6781) );
  OAI22_X1 U19222 ( .A1(n25640), .A2(n21222), .B1(n25970), .B2(n25633), .ZN(
        n6782) );
  OAI22_X1 U19223 ( .A1(n25447), .A2(n21101), .B1(n25963), .B2(n25440), .ZN(
        n5819) );
  OAI22_X1 U19224 ( .A1(n25447), .A2(n21100), .B1(n25966), .B2(n25440), .ZN(
        n5820) );
  OAI22_X1 U19225 ( .A1(n25447), .A2(n21099), .B1(n25969), .B2(n25440), .ZN(
        n5821) );
  OAI22_X1 U19226 ( .A1(n25447), .A2(n21098), .B1(n25972), .B2(n25440), .ZN(
        n5822) );
  OAI22_X1 U19227 ( .A1(n25408), .A2(n21097), .B1(n25963), .B2(n25401), .ZN(
        n5627) );
  OAI22_X1 U19228 ( .A1(n25408), .A2(n21096), .B1(n25966), .B2(n25401), .ZN(
        n5628) );
  OAI22_X1 U19229 ( .A1(n25408), .A2(n21095), .B1(n25969), .B2(n25401), .ZN(
        n5629) );
  OAI22_X1 U19230 ( .A1(n25408), .A2(n21094), .B1(n25972), .B2(n25401), .ZN(
        n5630) );
  OAI22_X1 U19231 ( .A1(n25768), .A2(n20969), .B1(n25961), .B2(n25761), .ZN(
        n7419) );
  OAI22_X1 U19232 ( .A1(n25768), .A2(n20968), .B1(n25964), .B2(n25761), .ZN(
        n7420) );
  OAI22_X1 U19233 ( .A1(n25768), .A2(n20967), .B1(n25967), .B2(n25761), .ZN(
        n7421) );
  OAI22_X1 U19234 ( .A1(n25768), .A2(n20966), .B1(n25970), .B2(n25761), .ZN(
        n7422) );
  OAI22_X1 U19235 ( .A1(n25537), .A2(n20713), .B1(n25962), .B2(n25530), .ZN(
        n6267) );
  OAI22_X1 U19236 ( .A1(n25537), .A2(n20712), .B1(n25965), .B2(n25530), .ZN(
        n6268) );
  OAI22_X1 U19237 ( .A1(n25537), .A2(n20711), .B1(n25968), .B2(n25530), .ZN(
        n6269) );
  OAI22_X1 U19238 ( .A1(n25537), .A2(n20710), .B1(n25971), .B2(n25530), .ZN(
        n6270) );
  OAI22_X1 U19239 ( .A1(n25730), .A2(n20649), .B1(n25961), .B2(n25723), .ZN(
        n7227) );
  OAI22_X1 U19240 ( .A1(n25730), .A2(n20648), .B1(n25964), .B2(n25723), .ZN(
        n7228) );
  OAI22_X1 U19241 ( .A1(n25730), .A2(n20647), .B1(n25967), .B2(n25723), .ZN(
        n7229) );
  OAI22_X1 U19242 ( .A1(n25730), .A2(n20646), .B1(n25970), .B2(n25723), .ZN(
        n7230) );
  OAI22_X1 U19243 ( .A1(n25627), .A2(n20401), .B1(n25962), .B2(n25620), .ZN(
        n6715) );
  OAI22_X1 U19244 ( .A1(n25627), .A2(n20400), .B1(n25965), .B2(n25620), .ZN(
        n6716) );
  OAI22_X1 U19245 ( .A1(n25627), .A2(n20399), .B1(n25968), .B2(n25620), .ZN(
        n6717) );
  OAI22_X1 U19246 ( .A1(n25627), .A2(n20398), .B1(n25971), .B2(n25620), .ZN(
        n6718) );
  OAI22_X1 U19247 ( .A1(n25550), .A2(n20337), .B1(n25962), .B2(n25543), .ZN(
        n6331) );
  OAI22_X1 U19248 ( .A1(n25550), .A2(n20336), .B1(n25965), .B2(n25543), .ZN(
        n6332) );
  OAI22_X1 U19249 ( .A1(n25550), .A2(n20335), .B1(n25968), .B2(n25543), .ZN(
        n6333) );
  OAI22_X1 U19250 ( .A1(n25550), .A2(n20334), .B1(n25971), .B2(n25543), .ZN(
        n6334) );
  OAI22_X1 U19251 ( .A1(n25524), .A2(n20273), .B1(n25962), .B2(n25517), .ZN(
        n6203) );
  OAI22_X1 U19252 ( .A1(n25524), .A2(n20272), .B1(n25965), .B2(n25517), .ZN(
        n6204) );
  OAI22_X1 U19253 ( .A1(n25524), .A2(n20271), .B1(n25968), .B2(n25517), .ZN(
        n6205) );
  OAI22_X1 U19254 ( .A1(n25524), .A2(n20270), .B1(n25971), .B2(n25517), .ZN(
        n6206) );
  OAI22_X1 U19255 ( .A1(n25434), .A2(n20137), .B1(n25963), .B2(n25427), .ZN(
        n5755) );
  OAI22_X1 U19256 ( .A1(n25434), .A2(n20136), .B1(n25966), .B2(n25427), .ZN(
        n5756) );
  OAI22_X1 U19257 ( .A1(n25434), .A2(n20135), .B1(n25969), .B2(n25427), .ZN(
        n5757) );
  OAI22_X1 U19258 ( .A1(n25434), .A2(n20134), .B1(n25972), .B2(n25427), .ZN(
        n5758) );
  OAI22_X1 U19259 ( .A1(n25666), .A2(n20133), .B1(n25970), .B2(n25659), .ZN(
        n6910) );
  OAI22_X1 U19260 ( .A1(n25614), .A2(n19816), .B1(n25962), .B2(n25607), .ZN(
        n6651) );
  OAI22_X1 U19261 ( .A1(n25614), .A2(n19815), .B1(n25965), .B2(n25607), .ZN(
        n6652) );
  OAI22_X1 U19262 ( .A1(n25614), .A2(n19814), .B1(n25968), .B2(n25607), .ZN(
        n6653) );
  OAI22_X1 U19263 ( .A1(n25614), .A2(n19813), .B1(n25971), .B2(n25607), .ZN(
        n6654) );
  OAI22_X1 U19264 ( .A1(n25666), .A2(n19752), .B1(n25961), .B2(n25659), .ZN(
        n6907) );
  OAI22_X1 U19265 ( .A1(n25666), .A2(n19751), .B1(n25964), .B2(n25659), .ZN(
        n6908) );
  OAI22_X1 U19266 ( .A1(n25666), .A2(n19750), .B1(n25967), .B2(n25659), .ZN(
        n6909) );
  OAI22_X1 U19267 ( .A1(n25717), .A2(n19561), .B1(n25961), .B2(n25710), .ZN(
        n7163) );
  OAI22_X1 U19268 ( .A1(n25717), .A2(n19560), .B1(n25964), .B2(n25710), .ZN(
        n7164) );
  OAI22_X1 U19269 ( .A1(n25717), .A2(n19559), .B1(n25967), .B2(n25710), .ZN(
        n7165) );
  OAI22_X1 U19270 ( .A1(n25717), .A2(n19558), .B1(n25970), .B2(n25710), .ZN(
        n7166) );
  OAI22_X1 U19271 ( .A1(n25443), .A2(n21221), .B1(n25783), .B2(n25435), .ZN(
        n5759) );
  OAI22_X1 U19272 ( .A1(n25443), .A2(n21220), .B1(n25786), .B2(n25435), .ZN(
        n5760) );
  OAI22_X1 U19273 ( .A1(n25443), .A2(n21219), .B1(n25789), .B2(n25435), .ZN(
        n5761) );
  OAI22_X1 U19274 ( .A1(n25443), .A2(n21218), .B1(n25792), .B2(n25435), .ZN(
        n5762) );
  OAI22_X1 U19275 ( .A1(n25443), .A2(n21217), .B1(n25795), .B2(n25435), .ZN(
        n5763) );
  OAI22_X1 U19276 ( .A1(n25443), .A2(n21216), .B1(n25798), .B2(n25435), .ZN(
        n5764) );
  OAI22_X1 U19277 ( .A1(n25443), .A2(n21215), .B1(n25801), .B2(n25435), .ZN(
        n5765) );
  OAI22_X1 U19278 ( .A1(n25443), .A2(n21214), .B1(n25804), .B2(n25435), .ZN(
        n5766) );
  OAI22_X1 U19279 ( .A1(n25443), .A2(n21213), .B1(n25807), .B2(n25435), .ZN(
        n5767) );
  OAI22_X1 U19280 ( .A1(n25443), .A2(n21212), .B1(n25810), .B2(n25435), .ZN(
        n5768) );
  OAI22_X1 U19281 ( .A1(n25443), .A2(n21211), .B1(n25813), .B2(n25435), .ZN(
        n5769) );
  OAI22_X1 U19282 ( .A1(n25443), .A2(n21210), .B1(n25816), .B2(n25435), .ZN(
        n5770) );
  OAI22_X1 U19283 ( .A1(n25444), .A2(n21209), .B1(n25819), .B2(n25436), .ZN(
        n5771) );
  OAI22_X1 U19284 ( .A1(n25444), .A2(n21208), .B1(n25822), .B2(n25436), .ZN(
        n5772) );
  OAI22_X1 U19285 ( .A1(n25444), .A2(n21207), .B1(n25825), .B2(n25436), .ZN(
        n5773) );
  OAI22_X1 U19286 ( .A1(n25444), .A2(n21206), .B1(n25828), .B2(n25436), .ZN(
        n5774) );
  OAI22_X1 U19287 ( .A1(n25444), .A2(n21205), .B1(n25831), .B2(n25436), .ZN(
        n5775) );
  OAI22_X1 U19288 ( .A1(n25444), .A2(n21204), .B1(n25834), .B2(n25436), .ZN(
        n5776) );
  OAI22_X1 U19289 ( .A1(n25444), .A2(n21203), .B1(n25837), .B2(n25436), .ZN(
        n5777) );
  OAI22_X1 U19290 ( .A1(n25444), .A2(n21202), .B1(n25840), .B2(n25436), .ZN(
        n5778) );
  OAI22_X1 U19291 ( .A1(n25444), .A2(n21201), .B1(n25843), .B2(n25436), .ZN(
        n5779) );
  OAI22_X1 U19292 ( .A1(n25444), .A2(n21200), .B1(n25846), .B2(n25436), .ZN(
        n5780) );
  OAI22_X1 U19293 ( .A1(n25444), .A2(n21199), .B1(n25849), .B2(n25436), .ZN(
        n5781) );
  OAI22_X1 U19294 ( .A1(n25444), .A2(n21198), .B1(n25852), .B2(n25436), .ZN(
        n5782) );
  OAI22_X1 U19295 ( .A1(n25444), .A2(n21197), .B1(n25855), .B2(n25437), .ZN(
        n5783) );
  OAI22_X1 U19296 ( .A1(n25445), .A2(n21196), .B1(n25858), .B2(n25437), .ZN(
        n5784) );
  OAI22_X1 U19297 ( .A1(n25445), .A2(n21195), .B1(n25861), .B2(n25437), .ZN(
        n5785) );
  OAI22_X1 U19298 ( .A1(n25445), .A2(n21194), .B1(n25864), .B2(n25437), .ZN(
        n5786) );
  OAI22_X1 U19299 ( .A1(n25445), .A2(n21193), .B1(n25867), .B2(n25437), .ZN(
        n5787) );
  OAI22_X1 U19300 ( .A1(n25445), .A2(n21192), .B1(n25870), .B2(n25437), .ZN(
        n5788) );
  OAI22_X1 U19301 ( .A1(n25445), .A2(n21191), .B1(n25873), .B2(n25437), .ZN(
        n5789) );
  OAI22_X1 U19302 ( .A1(n25445), .A2(n21190), .B1(n25876), .B2(n25437), .ZN(
        n5790) );
  OAI22_X1 U19303 ( .A1(n25445), .A2(n21189), .B1(n25879), .B2(n25437), .ZN(
        n5791) );
  OAI22_X1 U19304 ( .A1(n25445), .A2(n21188), .B1(n25882), .B2(n25437), .ZN(
        n5792) );
  OAI22_X1 U19305 ( .A1(n25445), .A2(n21187), .B1(n25885), .B2(n25437), .ZN(
        n5793) );
  OAI22_X1 U19306 ( .A1(n25445), .A2(n21186), .B1(n25888), .B2(n25437), .ZN(
        n5794) );
  OAI22_X1 U19307 ( .A1(n25445), .A2(n21185), .B1(n25891), .B2(n25438), .ZN(
        n5795) );
  OAI22_X1 U19308 ( .A1(n25445), .A2(n21184), .B1(n25894), .B2(n25438), .ZN(
        n5796) );
  OAI22_X1 U19309 ( .A1(n25446), .A2(n21183), .B1(n25897), .B2(n25438), .ZN(
        n5797) );
  OAI22_X1 U19310 ( .A1(n25446), .A2(n21182), .B1(n25900), .B2(n25438), .ZN(
        n5798) );
  OAI22_X1 U19311 ( .A1(n25446), .A2(n21181), .B1(n25903), .B2(n25438), .ZN(
        n5799) );
  OAI22_X1 U19312 ( .A1(n25446), .A2(n21180), .B1(n25906), .B2(n25438), .ZN(
        n5800) );
  OAI22_X1 U19313 ( .A1(n25446), .A2(n21179), .B1(n25909), .B2(n25438), .ZN(
        n5801) );
  OAI22_X1 U19314 ( .A1(n25446), .A2(n21178), .B1(n25912), .B2(n25438), .ZN(
        n5802) );
  OAI22_X1 U19315 ( .A1(n25446), .A2(n21177), .B1(n25915), .B2(n25438), .ZN(
        n5803) );
  OAI22_X1 U19316 ( .A1(n25446), .A2(n21176), .B1(n25918), .B2(n25438), .ZN(
        n5804) );
  OAI22_X1 U19317 ( .A1(n25446), .A2(n21175), .B1(n25921), .B2(n25438), .ZN(
        n5805) );
  OAI22_X1 U19318 ( .A1(n25446), .A2(n21174), .B1(n25924), .B2(n25438), .ZN(
        n5806) );
  OAI22_X1 U19319 ( .A1(n25446), .A2(n21173), .B1(n25927), .B2(n25439), .ZN(
        n5807) );
  OAI22_X1 U19320 ( .A1(n25446), .A2(n21172), .B1(n25930), .B2(n25439), .ZN(
        n5808) );
  OAI22_X1 U19321 ( .A1(n25446), .A2(n21171), .B1(n25933), .B2(n25439), .ZN(
        n5809) );
  OAI22_X1 U19322 ( .A1(n25447), .A2(n21170), .B1(n25936), .B2(n25439), .ZN(
        n5810) );
  OAI22_X1 U19323 ( .A1(n25447), .A2(n21169), .B1(n25939), .B2(n25439), .ZN(
        n5811) );
  OAI22_X1 U19324 ( .A1(n25447), .A2(n21168), .B1(n25942), .B2(n25439), .ZN(
        n5812) );
  OAI22_X1 U19325 ( .A1(n25447), .A2(n21167), .B1(n25945), .B2(n25439), .ZN(
        n5813) );
  OAI22_X1 U19326 ( .A1(n25447), .A2(n21166), .B1(n25948), .B2(n25439), .ZN(
        n5814) );
  OAI22_X1 U19327 ( .A1(n25447), .A2(n21165), .B1(n25951), .B2(n25439), .ZN(
        n5815) );
  OAI22_X1 U19328 ( .A1(n25447), .A2(n21164), .B1(n25954), .B2(n25439), .ZN(
        n5816) );
  OAI22_X1 U19329 ( .A1(n25447), .A2(n21163), .B1(n25957), .B2(n25439), .ZN(
        n5817) );
  OAI22_X1 U19330 ( .A1(n25447), .A2(n21162), .B1(n25960), .B2(n25439), .ZN(
        n5818) );
  OAI22_X1 U19331 ( .A1(n25404), .A2(n21161), .B1(n25783), .B2(n25396), .ZN(
        n5567) );
  OAI22_X1 U19332 ( .A1(n25404), .A2(n21160), .B1(n25786), .B2(n25396), .ZN(
        n5568) );
  OAI22_X1 U19333 ( .A1(n25404), .A2(n21159), .B1(n25789), .B2(n25396), .ZN(
        n5569) );
  OAI22_X1 U19334 ( .A1(n25404), .A2(n21158), .B1(n25792), .B2(n25396), .ZN(
        n5570) );
  OAI22_X1 U19335 ( .A1(n25404), .A2(n21157), .B1(n25795), .B2(n25396), .ZN(
        n5571) );
  OAI22_X1 U19336 ( .A1(n25404), .A2(n21156), .B1(n25798), .B2(n25396), .ZN(
        n5572) );
  OAI22_X1 U19337 ( .A1(n25404), .A2(n21155), .B1(n25801), .B2(n25396), .ZN(
        n5573) );
  OAI22_X1 U19338 ( .A1(n25404), .A2(n21154), .B1(n25804), .B2(n25396), .ZN(
        n5574) );
  OAI22_X1 U19339 ( .A1(n25404), .A2(n21153), .B1(n25807), .B2(n25396), .ZN(
        n5575) );
  OAI22_X1 U19340 ( .A1(n25404), .A2(n21152), .B1(n25810), .B2(n25396), .ZN(
        n5576) );
  OAI22_X1 U19341 ( .A1(n25404), .A2(n21151), .B1(n25813), .B2(n25396), .ZN(
        n5577) );
  OAI22_X1 U19342 ( .A1(n25404), .A2(n21150), .B1(n25816), .B2(n25396), .ZN(
        n5578) );
  OAI22_X1 U19343 ( .A1(n25405), .A2(n21149), .B1(n25819), .B2(n25397), .ZN(
        n5579) );
  OAI22_X1 U19344 ( .A1(n25405), .A2(n21148), .B1(n25822), .B2(n25397), .ZN(
        n5580) );
  OAI22_X1 U19345 ( .A1(n25405), .A2(n21147), .B1(n25825), .B2(n25397), .ZN(
        n5581) );
  OAI22_X1 U19346 ( .A1(n25405), .A2(n21146), .B1(n25828), .B2(n25397), .ZN(
        n5582) );
  OAI22_X1 U19347 ( .A1(n25405), .A2(n21145), .B1(n25831), .B2(n25397), .ZN(
        n5583) );
  OAI22_X1 U19348 ( .A1(n25405), .A2(n21144), .B1(n25834), .B2(n25397), .ZN(
        n5584) );
  OAI22_X1 U19349 ( .A1(n25405), .A2(n21143), .B1(n25837), .B2(n25397), .ZN(
        n5585) );
  OAI22_X1 U19350 ( .A1(n25405), .A2(n21142), .B1(n25840), .B2(n25397), .ZN(
        n5586) );
  OAI22_X1 U19351 ( .A1(n25405), .A2(n21141), .B1(n25843), .B2(n25397), .ZN(
        n5587) );
  OAI22_X1 U19352 ( .A1(n25405), .A2(n21140), .B1(n25846), .B2(n25397), .ZN(
        n5588) );
  OAI22_X1 U19353 ( .A1(n25405), .A2(n21139), .B1(n25849), .B2(n25397), .ZN(
        n5589) );
  OAI22_X1 U19354 ( .A1(n25405), .A2(n21138), .B1(n25852), .B2(n25397), .ZN(
        n5590) );
  OAI22_X1 U19355 ( .A1(n25405), .A2(n21137), .B1(n25855), .B2(n25398), .ZN(
        n5591) );
  OAI22_X1 U19356 ( .A1(n25406), .A2(n21136), .B1(n25858), .B2(n25398), .ZN(
        n5592) );
  OAI22_X1 U19357 ( .A1(n25406), .A2(n21135), .B1(n25861), .B2(n25398), .ZN(
        n5593) );
  OAI22_X1 U19358 ( .A1(n25406), .A2(n21134), .B1(n25864), .B2(n25398), .ZN(
        n5594) );
  OAI22_X1 U19359 ( .A1(n25406), .A2(n21133), .B1(n25867), .B2(n25398), .ZN(
        n5595) );
  OAI22_X1 U19360 ( .A1(n25406), .A2(n21132), .B1(n25870), .B2(n25398), .ZN(
        n5596) );
  OAI22_X1 U19361 ( .A1(n25406), .A2(n21131), .B1(n25873), .B2(n25398), .ZN(
        n5597) );
  OAI22_X1 U19362 ( .A1(n25406), .A2(n21130), .B1(n25876), .B2(n25398), .ZN(
        n5598) );
  OAI22_X1 U19363 ( .A1(n25406), .A2(n21129), .B1(n25879), .B2(n25398), .ZN(
        n5599) );
  OAI22_X1 U19364 ( .A1(n25406), .A2(n21128), .B1(n25882), .B2(n25398), .ZN(
        n5600) );
  OAI22_X1 U19365 ( .A1(n25406), .A2(n21127), .B1(n25885), .B2(n25398), .ZN(
        n5601) );
  OAI22_X1 U19366 ( .A1(n25406), .A2(n21126), .B1(n25888), .B2(n25398), .ZN(
        n5602) );
  OAI22_X1 U19367 ( .A1(n25406), .A2(n21125), .B1(n25891), .B2(n25399), .ZN(
        n5603) );
  OAI22_X1 U19368 ( .A1(n25406), .A2(n21124), .B1(n25894), .B2(n25399), .ZN(
        n5604) );
  OAI22_X1 U19369 ( .A1(n25407), .A2(n21123), .B1(n25897), .B2(n25399), .ZN(
        n5605) );
  OAI22_X1 U19370 ( .A1(n25407), .A2(n21122), .B1(n25900), .B2(n25399), .ZN(
        n5606) );
  OAI22_X1 U19371 ( .A1(n25407), .A2(n21121), .B1(n25903), .B2(n25399), .ZN(
        n5607) );
  OAI22_X1 U19372 ( .A1(n25407), .A2(n21120), .B1(n25906), .B2(n25399), .ZN(
        n5608) );
  OAI22_X1 U19373 ( .A1(n25407), .A2(n21119), .B1(n25909), .B2(n25399), .ZN(
        n5609) );
  OAI22_X1 U19374 ( .A1(n25407), .A2(n21118), .B1(n25912), .B2(n25399), .ZN(
        n5610) );
  OAI22_X1 U19375 ( .A1(n25407), .A2(n21117), .B1(n25915), .B2(n25399), .ZN(
        n5611) );
  OAI22_X1 U19376 ( .A1(n25407), .A2(n21116), .B1(n25918), .B2(n25399), .ZN(
        n5612) );
  OAI22_X1 U19377 ( .A1(n25407), .A2(n21115), .B1(n25921), .B2(n25399), .ZN(
        n5613) );
  OAI22_X1 U19378 ( .A1(n25407), .A2(n21114), .B1(n25924), .B2(n25399), .ZN(
        n5614) );
  OAI22_X1 U19379 ( .A1(n25407), .A2(n21113), .B1(n25927), .B2(n25400), .ZN(
        n5615) );
  OAI22_X1 U19380 ( .A1(n25407), .A2(n21112), .B1(n25930), .B2(n25400), .ZN(
        n5616) );
  OAI22_X1 U19381 ( .A1(n25407), .A2(n21111), .B1(n25933), .B2(n25400), .ZN(
        n5617) );
  OAI22_X1 U19382 ( .A1(n25408), .A2(n21110), .B1(n25936), .B2(n25400), .ZN(
        n5618) );
  OAI22_X1 U19383 ( .A1(n25408), .A2(n21109), .B1(n25939), .B2(n25400), .ZN(
        n5619) );
  OAI22_X1 U19384 ( .A1(n25408), .A2(n21108), .B1(n25942), .B2(n25400), .ZN(
        n5620) );
  OAI22_X1 U19385 ( .A1(n25408), .A2(n21107), .B1(n25945), .B2(n25400), .ZN(
        n5621) );
  OAI22_X1 U19386 ( .A1(n25408), .A2(n21106), .B1(n25948), .B2(n25400), .ZN(
        n5622) );
  OAI22_X1 U19387 ( .A1(n25408), .A2(n21105), .B1(n25951), .B2(n25400), .ZN(
        n5623) );
  OAI22_X1 U19388 ( .A1(n25408), .A2(n21104), .B1(n25954), .B2(n25400), .ZN(
        n5624) );
  OAI22_X1 U19389 ( .A1(n25408), .A2(n21103), .B1(n25957), .B2(n25400), .ZN(
        n5625) );
  OAI22_X1 U19390 ( .A1(n25408), .A2(n21102), .B1(n25960), .B2(n25400), .ZN(
        n5626) );
  OAI22_X1 U19391 ( .A1(n25430), .A2(n20197), .B1(n25783), .B2(n25422), .ZN(
        n5695) );
  OAI22_X1 U19392 ( .A1(n25430), .A2(n20196), .B1(n25786), .B2(n25422), .ZN(
        n5696) );
  OAI22_X1 U19393 ( .A1(n25430), .A2(n20195), .B1(n25789), .B2(n25422), .ZN(
        n5697) );
  OAI22_X1 U19394 ( .A1(n25430), .A2(n20194), .B1(n25792), .B2(n25422), .ZN(
        n5698) );
  OAI22_X1 U19395 ( .A1(n25430), .A2(n20193), .B1(n25795), .B2(n25422), .ZN(
        n5699) );
  OAI22_X1 U19396 ( .A1(n25430), .A2(n20192), .B1(n25798), .B2(n25422), .ZN(
        n5700) );
  OAI22_X1 U19397 ( .A1(n25430), .A2(n20191), .B1(n25801), .B2(n25422), .ZN(
        n5701) );
  OAI22_X1 U19398 ( .A1(n25430), .A2(n20190), .B1(n25804), .B2(n25422), .ZN(
        n5702) );
  OAI22_X1 U19399 ( .A1(n25430), .A2(n20189), .B1(n25807), .B2(n25422), .ZN(
        n5703) );
  OAI22_X1 U19400 ( .A1(n25430), .A2(n20188), .B1(n25810), .B2(n25422), .ZN(
        n5704) );
  OAI22_X1 U19401 ( .A1(n25430), .A2(n20187), .B1(n25813), .B2(n25422), .ZN(
        n5705) );
  OAI22_X1 U19402 ( .A1(n25430), .A2(n20186), .B1(n25816), .B2(n25422), .ZN(
        n5706) );
  OAI22_X1 U19403 ( .A1(n25431), .A2(n20185), .B1(n25819), .B2(n25423), .ZN(
        n5707) );
  OAI22_X1 U19404 ( .A1(n25431), .A2(n20184), .B1(n25822), .B2(n25423), .ZN(
        n5708) );
  OAI22_X1 U19405 ( .A1(n25431), .A2(n20183), .B1(n25825), .B2(n25423), .ZN(
        n5709) );
  OAI22_X1 U19406 ( .A1(n25431), .A2(n20182), .B1(n25828), .B2(n25423), .ZN(
        n5710) );
  OAI22_X1 U19407 ( .A1(n25431), .A2(n20181), .B1(n25831), .B2(n25423), .ZN(
        n5711) );
  OAI22_X1 U19408 ( .A1(n25431), .A2(n20180), .B1(n25834), .B2(n25423), .ZN(
        n5712) );
  OAI22_X1 U19409 ( .A1(n25431), .A2(n20179), .B1(n25837), .B2(n25423), .ZN(
        n5713) );
  OAI22_X1 U19410 ( .A1(n25431), .A2(n20178), .B1(n25840), .B2(n25423), .ZN(
        n5714) );
  OAI22_X1 U19411 ( .A1(n25431), .A2(n20177), .B1(n25843), .B2(n25423), .ZN(
        n5715) );
  OAI22_X1 U19412 ( .A1(n25431), .A2(n20176), .B1(n25846), .B2(n25423), .ZN(
        n5716) );
  OAI22_X1 U19413 ( .A1(n25431), .A2(n20175), .B1(n25849), .B2(n25423), .ZN(
        n5717) );
  OAI22_X1 U19414 ( .A1(n25431), .A2(n20174), .B1(n25852), .B2(n25423), .ZN(
        n5718) );
  OAI22_X1 U19415 ( .A1(n25431), .A2(n20173), .B1(n25855), .B2(n25424), .ZN(
        n5719) );
  OAI22_X1 U19416 ( .A1(n25432), .A2(n20172), .B1(n25858), .B2(n25424), .ZN(
        n5720) );
  OAI22_X1 U19417 ( .A1(n25432), .A2(n20171), .B1(n25861), .B2(n25424), .ZN(
        n5721) );
  OAI22_X1 U19418 ( .A1(n25432), .A2(n20170), .B1(n25864), .B2(n25424), .ZN(
        n5722) );
  OAI22_X1 U19419 ( .A1(n25432), .A2(n20169), .B1(n25867), .B2(n25424), .ZN(
        n5723) );
  OAI22_X1 U19420 ( .A1(n25432), .A2(n20168), .B1(n25870), .B2(n25424), .ZN(
        n5724) );
  OAI22_X1 U19421 ( .A1(n25432), .A2(n20167), .B1(n25873), .B2(n25424), .ZN(
        n5725) );
  OAI22_X1 U19422 ( .A1(n25432), .A2(n20166), .B1(n25876), .B2(n25424), .ZN(
        n5726) );
  OAI22_X1 U19423 ( .A1(n25432), .A2(n20165), .B1(n25879), .B2(n25424), .ZN(
        n5727) );
  OAI22_X1 U19424 ( .A1(n25432), .A2(n20164), .B1(n25882), .B2(n25424), .ZN(
        n5728) );
  OAI22_X1 U19425 ( .A1(n25432), .A2(n20163), .B1(n25885), .B2(n25424), .ZN(
        n5729) );
  OAI22_X1 U19426 ( .A1(n25432), .A2(n20162), .B1(n25888), .B2(n25424), .ZN(
        n5730) );
  OAI22_X1 U19427 ( .A1(n25432), .A2(n20161), .B1(n25891), .B2(n25425), .ZN(
        n5731) );
  OAI22_X1 U19428 ( .A1(n25432), .A2(n20160), .B1(n25894), .B2(n25425), .ZN(
        n5732) );
  OAI22_X1 U19429 ( .A1(n25433), .A2(n20159), .B1(n25897), .B2(n25425), .ZN(
        n5733) );
  OAI22_X1 U19430 ( .A1(n25433), .A2(n20158), .B1(n25900), .B2(n25425), .ZN(
        n5734) );
  OAI22_X1 U19431 ( .A1(n25433), .A2(n20157), .B1(n25903), .B2(n25425), .ZN(
        n5735) );
  OAI22_X1 U19432 ( .A1(n25433), .A2(n20156), .B1(n25906), .B2(n25425), .ZN(
        n5736) );
  OAI22_X1 U19433 ( .A1(n25433), .A2(n20155), .B1(n25909), .B2(n25425), .ZN(
        n5737) );
  OAI22_X1 U19434 ( .A1(n25433), .A2(n20154), .B1(n25912), .B2(n25425), .ZN(
        n5738) );
  OAI22_X1 U19435 ( .A1(n25433), .A2(n20153), .B1(n25915), .B2(n25425), .ZN(
        n5739) );
  OAI22_X1 U19436 ( .A1(n25433), .A2(n20152), .B1(n25918), .B2(n25425), .ZN(
        n5740) );
  OAI22_X1 U19437 ( .A1(n25433), .A2(n20151), .B1(n25921), .B2(n25425), .ZN(
        n5741) );
  OAI22_X1 U19438 ( .A1(n25433), .A2(n20150), .B1(n25924), .B2(n25425), .ZN(
        n5742) );
  OAI22_X1 U19439 ( .A1(n25433), .A2(n20149), .B1(n25927), .B2(n25426), .ZN(
        n5743) );
  OAI22_X1 U19440 ( .A1(n25433), .A2(n20148), .B1(n25930), .B2(n25426), .ZN(
        n5744) );
  OAI22_X1 U19441 ( .A1(n25433), .A2(n20147), .B1(n25933), .B2(n25426), .ZN(
        n5745) );
  OAI22_X1 U19442 ( .A1(n25434), .A2(n20146), .B1(n25936), .B2(n25426), .ZN(
        n5746) );
  OAI22_X1 U19443 ( .A1(n25434), .A2(n20145), .B1(n25939), .B2(n25426), .ZN(
        n5747) );
  OAI22_X1 U19444 ( .A1(n25434), .A2(n20144), .B1(n25942), .B2(n25426), .ZN(
        n5748) );
  OAI22_X1 U19445 ( .A1(n25434), .A2(n20143), .B1(n25945), .B2(n25426), .ZN(
        n5749) );
  OAI22_X1 U19446 ( .A1(n25434), .A2(n20142), .B1(n25948), .B2(n25426), .ZN(
        n5750) );
  OAI22_X1 U19447 ( .A1(n25434), .A2(n20141), .B1(n25951), .B2(n25426), .ZN(
        n5751) );
  OAI22_X1 U19448 ( .A1(n25434), .A2(n20140), .B1(n25954), .B2(n25426), .ZN(
        n5752) );
  OAI22_X1 U19449 ( .A1(n25434), .A2(n20139), .B1(n25957), .B2(n25426), .ZN(
        n5753) );
  OAI22_X1 U19450 ( .A1(n25434), .A2(n20138), .B1(n25960), .B2(n25426), .ZN(
        n5754) );
  OAI22_X1 U19451 ( .A1(n25559), .A2(n21413), .B1(n25782), .B2(n25551), .ZN(
        n6335) );
  OAI22_X1 U19452 ( .A1(n25559), .A2(n21412), .B1(n25785), .B2(n25551), .ZN(
        n6336) );
  OAI22_X1 U19453 ( .A1(n25559), .A2(n21411), .B1(n25788), .B2(n25551), .ZN(
        n6337) );
  OAI22_X1 U19454 ( .A1(n25559), .A2(n21410), .B1(n25791), .B2(n25551), .ZN(
        n6338) );
  OAI22_X1 U19455 ( .A1(n25559), .A2(n21409), .B1(n25794), .B2(n25551), .ZN(
        n6339) );
  OAI22_X1 U19456 ( .A1(n25559), .A2(n21408), .B1(n25797), .B2(n25551), .ZN(
        n6340) );
  OAI22_X1 U19457 ( .A1(n25559), .A2(n21407), .B1(n25800), .B2(n25551), .ZN(
        n6341) );
  OAI22_X1 U19458 ( .A1(n25559), .A2(n21406), .B1(n25803), .B2(n25551), .ZN(
        n6342) );
  OAI22_X1 U19459 ( .A1(n25559), .A2(n21405), .B1(n25806), .B2(n25551), .ZN(
        n6343) );
  OAI22_X1 U19460 ( .A1(n25559), .A2(n21404), .B1(n25809), .B2(n25551), .ZN(
        n6344) );
  OAI22_X1 U19461 ( .A1(n25559), .A2(n21403), .B1(n25812), .B2(n25551), .ZN(
        n6345) );
  OAI22_X1 U19462 ( .A1(n25559), .A2(n21402), .B1(n25815), .B2(n25551), .ZN(
        n6346) );
  OAI22_X1 U19463 ( .A1(n25560), .A2(n21401), .B1(n25818), .B2(n25552), .ZN(
        n6347) );
  OAI22_X1 U19464 ( .A1(n25560), .A2(n21400), .B1(n25821), .B2(n25552), .ZN(
        n6348) );
  OAI22_X1 U19465 ( .A1(n25560), .A2(n21399), .B1(n25824), .B2(n25552), .ZN(
        n6349) );
  OAI22_X1 U19466 ( .A1(n25560), .A2(n21398), .B1(n25827), .B2(n25552), .ZN(
        n6350) );
  OAI22_X1 U19467 ( .A1(n25560), .A2(n21397), .B1(n25830), .B2(n25552), .ZN(
        n6351) );
  OAI22_X1 U19468 ( .A1(n25560), .A2(n21396), .B1(n25833), .B2(n25552), .ZN(
        n6352) );
  OAI22_X1 U19469 ( .A1(n25560), .A2(n21395), .B1(n25836), .B2(n25552), .ZN(
        n6353) );
  OAI22_X1 U19470 ( .A1(n25560), .A2(n21394), .B1(n25839), .B2(n25552), .ZN(
        n6354) );
  OAI22_X1 U19471 ( .A1(n25560), .A2(n21393), .B1(n25842), .B2(n25552), .ZN(
        n6355) );
  OAI22_X1 U19472 ( .A1(n25560), .A2(n21392), .B1(n25845), .B2(n25552), .ZN(
        n6356) );
  OAI22_X1 U19473 ( .A1(n25560), .A2(n21391), .B1(n25848), .B2(n25552), .ZN(
        n6357) );
  OAI22_X1 U19474 ( .A1(n25560), .A2(n21390), .B1(n25851), .B2(n25552), .ZN(
        n6358) );
  OAI22_X1 U19475 ( .A1(n25560), .A2(n21389), .B1(n25854), .B2(n25553), .ZN(
        n6359) );
  OAI22_X1 U19476 ( .A1(n25561), .A2(n21388), .B1(n25857), .B2(n25553), .ZN(
        n6360) );
  OAI22_X1 U19477 ( .A1(n25561), .A2(n21387), .B1(n25860), .B2(n25553), .ZN(
        n6361) );
  OAI22_X1 U19478 ( .A1(n25561), .A2(n21386), .B1(n25863), .B2(n25553), .ZN(
        n6362) );
  OAI22_X1 U19479 ( .A1(n25561), .A2(n21385), .B1(n25866), .B2(n25553), .ZN(
        n6363) );
  OAI22_X1 U19480 ( .A1(n25561), .A2(n21384), .B1(n25869), .B2(n25553), .ZN(
        n6364) );
  OAI22_X1 U19481 ( .A1(n25561), .A2(n21383), .B1(n25872), .B2(n25553), .ZN(
        n6365) );
  OAI22_X1 U19482 ( .A1(n25561), .A2(n21382), .B1(n25875), .B2(n25553), .ZN(
        n6366) );
  OAI22_X1 U19483 ( .A1(n25561), .A2(n21381), .B1(n25878), .B2(n25553), .ZN(
        n6367) );
  OAI22_X1 U19484 ( .A1(n25561), .A2(n21380), .B1(n25881), .B2(n25553), .ZN(
        n6368) );
  OAI22_X1 U19485 ( .A1(n25561), .A2(n21379), .B1(n25884), .B2(n25553), .ZN(
        n6369) );
  OAI22_X1 U19486 ( .A1(n25561), .A2(n21378), .B1(n25887), .B2(n25553), .ZN(
        n6370) );
  OAI22_X1 U19487 ( .A1(n25561), .A2(n21377), .B1(n25890), .B2(n25554), .ZN(
        n6371) );
  OAI22_X1 U19488 ( .A1(n25561), .A2(n21376), .B1(n25893), .B2(n25554), .ZN(
        n6372) );
  OAI22_X1 U19489 ( .A1(n25562), .A2(n21375), .B1(n25896), .B2(n25554), .ZN(
        n6373) );
  OAI22_X1 U19490 ( .A1(n25562), .A2(n21374), .B1(n25899), .B2(n25554), .ZN(
        n6374) );
  OAI22_X1 U19491 ( .A1(n25562), .A2(n21373), .B1(n25902), .B2(n25554), .ZN(
        n6375) );
  OAI22_X1 U19492 ( .A1(n25562), .A2(n21372), .B1(n25905), .B2(n25554), .ZN(
        n6376) );
  OAI22_X1 U19493 ( .A1(n25562), .A2(n21371), .B1(n25908), .B2(n25554), .ZN(
        n6377) );
  OAI22_X1 U19494 ( .A1(n25562), .A2(n21370), .B1(n25911), .B2(n25554), .ZN(
        n6378) );
  OAI22_X1 U19495 ( .A1(n25562), .A2(n21369), .B1(n25914), .B2(n25554), .ZN(
        n6379) );
  OAI22_X1 U19496 ( .A1(n25562), .A2(n21368), .B1(n25917), .B2(n25554), .ZN(
        n6380) );
  OAI22_X1 U19497 ( .A1(n25562), .A2(n21367), .B1(n25920), .B2(n25554), .ZN(
        n6381) );
  OAI22_X1 U19498 ( .A1(n25562), .A2(n21366), .B1(n25923), .B2(n25554), .ZN(
        n6382) );
  OAI22_X1 U19499 ( .A1(n25562), .A2(n21365), .B1(n25926), .B2(n25555), .ZN(
        n6383) );
  OAI22_X1 U19500 ( .A1(n25562), .A2(n21364), .B1(n25929), .B2(n25555), .ZN(
        n6384) );
  OAI22_X1 U19501 ( .A1(n25562), .A2(n21363), .B1(n25932), .B2(n25555), .ZN(
        n6385) );
  OAI22_X1 U19502 ( .A1(n25563), .A2(n21362), .B1(n25935), .B2(n25555), .ZN(
        n6386) );
  OAI22_X1 U19503 ( .A1(n25563), .A2(n21361), .B1(n25938), .B2(n25555), .ZN(
        n6387) );
  OAI22_X1 U19504 ( .A1(n25563), .A2(n21360), .B1(n25941), .B2(n25555), .ZN(
        n6388) );
  OAI22_X1 U19505 ( .A1(n25563), .A2(n21359), .B1(n25944), .B2(n25555), .ZN(
        n6389) );
  OAI22_X1 U19506 ( .A1(n25563), .A2(n21358), .B1(n25947), .B2(n25555), .ZN(
        n6390) );
  OAI22_X1 U19507 ( .A1(n25563), .A2(n21357), .B1(n25950), .B2(n25555), .ZN(
        n6391) );
  OAI22_X1 U19508 ( .A1(n25563), .A2(n21356), .B1(n25953), .B2(n25555), .ZN(
        n6392) );
  OAI22_X1 U19509 ( .A1(n25563), .A2(n21355), .B1(n25956), .B2(n25555), .ZN(
        n6393) );
  OAI22_X1 U19510 ( .A1(n25563), .A2(n21354), .B1(n25959), .B2(n25555), .ZN(
        n6394) );
  OAI22_X1 U19511 ( .A1(n25636), .A2(n21285), .B1(n25781), .B2(n25628), .ZN(
        n6719) );
  OAI22_X1 U19512 ( .A1(n25636), .A2(n21284), .B1(n25784), .B2(n25628), .ZN(
        n6720) );
  OAI22_X1 U19513 ( .A1(n25636), .A2(n21283), .B1(n25787), .B2(n25628), .ZN(
        n6721) );
  OAI22_X1 U19514 ( .A1(n25636), .A2(n21282), .B1(n25790), .B2(n25628), .ZN(
        n6722) );
  OAI22_X1 U19515 ( .A1(n25636), .A2(n21281), .B1(n25793), .B2(n25628), .ZN(
        n6723) );
  OAI22_X1 U19516 ( .A1(n25636), .A2(n21280), .B1(n25796), .B2(n25628), .ZN(
        n6724) );
  OAI22_X1 U19517 ( .A1(n25636), .A2(n21279), .B1(n25799), .B2(n25628), .ZN(
        n6725) );
  OAI22_X1 U19518 ( .A1(n25636), .A2(n21278), .B1(n25802), .B2(n25628), .ZN(
        n6726) );
  OAI22_X1 U19519 ( .A1(n25636), .A2(n21277), .B1(n25805), .B2(n25628), .ZN(
        n6727) );
  OAI22_X1 U19520 ( .A1(n25636), .A2(n21276), .B1(n25808), .B2(n25628), .ZN(
        n6728) );
  OAI22_X1 U19521 ( .A1(n25636), .A2(n21275), .B1(n25811), .B2(n25628), .ZN(
        n6729) );
  OAI22_X1 U19522 ( .A1(n25636), .A2(n21274), .B1(n25814), .B2(n25628), .ZN(
        n6730) );
  OAI22_X1 U19523 ( .A1(n25637), .A2(n21273), .B1(n25817), .B2(n25629), .ZN(
        n6731) );
  OAI22_X1 U19524 ( .A1(n25637), .A2(n21272), .B1(n25820), .B2(n25629), .ZN(
        n6732) );
  OAI22_X1 U19525 ( .A1(n25637), .A2(n21271), .B1(n25823), .B2(n25629), .ZN(
        n6733) );
  OAI22_X1 U19526 ( .A1(n25637), .A2(n21270), .B1(n25826), .B2(n25629), .ZN(
        n6734) );
  OAI22_X1 U19527 ( .A1(n25637), .A2(n21269), .B1(n25829), .B2(n25629), .ZN(
        n6735) );
  OAI22_X1 U19528 ( .A1(n25637), .A2(n21268), .B1(n25832), .B2(n25629), .ZN(
        n6736) );
  OAI22_X1 U19529 ( .A1(n25637), .A2(n21267), .B1(n25835), .B2(n25629), .ZN(
        n6737) );
  OAI22_X1 U19530 ( .A1(n25637), .A2(n21266), .B1(n25838), .B2(n25629), .ZN(
        n6738) );
  OAI22_X1 U19531 ( .A1(n25637), .A2(n21265), .B1(n25841), .B2(n25629), .ZN(
        n6739) );
  OAI22_X1 U19532 ( .A1(n25637), .A2(n21264), .B1(n25844), .B2(n25629), .ZN(
        n6740) );
  OAI22_X1 U19533 ( .A1(n25637), .A2(n21263), .B1(n25847), .B2(n25629), .ZN(
        n6741) );
  OAI22_X1 U19534 ( .A1(n25637), .A2(n21262), .B1(n25850), .B2(n25629), .ZN(
        n6742) );
  OAI22_X1 U19535 ( .A1(n25637), .A2(n21261), .B1(n25853), .B2(n25630), .ZN(
        n6743) );
  OAI22_X1 U19536 ( .A1(n25638), .A2(n21260), .B1(n25856), .B2(n25630), .ZN(
        n6744) );
  OAI22_X1 U19537 ( .A1(n25638), .A2(n21259), .B1(n25859), .B2(n25630), .ZN(
        n6745) );
  OAI22_X1 U19538 ( .A1(n25638), .A2(n21258), .B1(n25862), .B2(n25630), .ZN(
        n6746) );
  OAI22_X1 U19539 ( .A1(n25638), .A2(n21257), .B1(n25865), .B2(n25630), .ZN(
        n6747) );
  OAI22_X1 U19540 ( .A1(n25638), .A2(n21256), .B1(n25868), .B2(n25630), .ZN(
        n6748) );
  OAI22_X1 U19541 ( .A1(n25638), .A2(n21255), .B1(n25871), .B2(n25630), .ZN(
        n6749) );
  OAI22_X1 U19542 ( .A1(n25638), .A2(n21254), .B1(n25874), .B2(n25630), .ZN(
        n6750) );
  OAI22_X1 U19543 ( .A1(n25638), .A2(n21253), .B1(n25877), .B2(n25630), .ZN(
        n6751) );
  OAI22_X1 U19544 ( .A1(n25638), .A2(n21252), .B1(n25880), .B2(n25630), .ZN(
        n6752) );
  OAI22_X1 U19545 ( .A1(n25638), .A2(n21251), .B1(n25883), .B2(n25630), .ZN(
        n6753) );
  OAI22_X1 U19546 ( .A1(n25638), .A2(n21250), .B1(n25886), .B2(n25630), .ZN(
        n6754) );
  OAI22_X1 U19547 ( .A1(n25638), .A2(n21249), .B1(n25889), .B2(n25631), .ZN(
        n6755) );
  OAI22_X1 U19548 ( .A1(n25638), .A2(n21248), .B1(n25892), .B2(n25631), .ZN(
        n6756) );
  OAI22_X1 U19549 ( .A1(n25639), .A2(n21247), .B1(n25895), .B2(n25631), .ZN(
        n6757) );
  OAI22_X1 U19550 ( .A1(n25639), .A2(n21246), .B1(n25898), .B2(n25631), .ZN(
        n6758) );
  OAI22_X1 U19551 ( .A1(n25639), .A2(n21245), .B1(n25901), .B2(n25631), .ZN(
        n6759) );
  OAI22_X1 U19552 ( .A1(n25639), .A2(n21244), .B1(n25904), .B2(n25631), .ZN(
        n6760) );
  OAI22_X1 U19553 ( .A1(n25639), .A2(n21243), .B1(n25907), .B2(n25631), .ZN(
        n6761) );
  OAI22_X1 U19554 ( .A1(n25639), .A2(n21242), .B1(n25910), .B2(n25631), .ZN(
        n6762) );
  OAI22_X1 U19555 ( .A1(n25639), .A2(n21241), .B1(n25913), .B2(n25631), .ZN(
        n6763) );
  OAI22_X1 U19556 ( .A1(n25639), .A2(n21240), .B1(n25916), .B2(n25631), .ZN(
        n6764) );
  OAI22_X1 U19557 ( .A1(n25639), .A2(n21239), .B1(n25919), .B2(n25631), .ZN(
        n6765) );
  OAI22_X1 U19558 ( .A1(n25639), .A2(n21238), .B1(n25922), .B2(n25631), .ZN(
        n6766) );
  OAI22_X1 U19559 ( .A1(n25639), .A2(n21237), .B1(n25925), .B2(n25632), .ZN(
        n6767) );
  OAI22_X1 U19560 ( .A1(n25639), .A2(n21236), .B1(n25928), .B2(n25632), .ZN(
        n6768) );
  OAI22_X1 U19561 ( .A1(n25639), .A2(n21235), .B1(n25931), .B2(n25632), .ZN(
        n6769) );
  OAI22_X1 U19562 ( .A1(n25640), .A2(n21234), .B1(n25934), .B2(n25632), .ZN(
        n6770) );
  OAI22_X1 U19563 ( .A1(n25640), .A2(n21233), .B1(n25937), .B2(n25632), .ZN(
        n6771) );
  OAI22_X1 U19564 ( .A1(n25640), .A2(n21232), .B1(n25940), .B2(n25632), .ZN(
        n6772) );
  OAI22_X1 U19565 ( .A1(n25640), .A2(n21231), .B1(n25943), .B2(n25632), .ZN(
        n6773) );
  OAI22_X1 U19566 ( .A1(n25640), .A2(n21230), .B1(n25946), .B2(n25632), .ZN(
        n6774) );
  OAI22_X1 U19567 ( .A1(n25640), .A2(n21229), .B1(n25949), .B2(n25632), .ZN(
        n6775) );
  OAI22_X1 U19568 ( .A1(n25640), .A2(n21228), .B1(n25952), .B2(n25632), .ZN(
        n6776) );
  OAI22_X1 U19569 ( .A1(n25640), .A2(n21227), .B1(n25955), .B2(n25632), .ZN(
        n6777) );
  OAI22_X1 U19570 ( .A1(n25640), .A2(n21226), .B1(n25958), .B2(n25632), .ZN(
        n6778) );
  OAI22_X1 U19571 ( .A1(n25764), .A2(n21029), .B1(n25781), .B2(n25756), .ZN(
        n7359) );
  OAI22_X1 U19572 ( .A1(n25764), .A2(n21028), .B1(n25784), .B2(n25756), .ZN(
        n7360) );
  OAI22_X1 U19573 ( .A1(n25764), .A2(n21027), .B1(n25787), .B2(n25756), .ZN(
        n7361) );
  OAI22_X1 U19574 ( .A1(n25764), .A2(n21026), .B1(n25790), .B2(n25756), .ZN(
        n7362) );
  OAI22_X1 U19575 ( .A1(n25764), .A2(n21025), .B1(n25793), .B2(n25756), .ZN(
        n7363) );
  OAI22_X1 U19576 ( .A1(n25764), .A2(n21024), .B1(n25796), .B2(n25756), .ZN(
        n7364) );
  OAI22_X1 U19577 ( .A1(n25764), .A2(n21023), .B1(n25799), .B2(n25756), .ZN(
        n7365) );
  OAI22_X1 U19578 ( .A1(n25764), .A2(n21022), .B1(n25802), .B2(n25756), .ZN(
        n7366) );
  OAI22_X1 U19579 ( .A1(n25764), .A2(n21021), .B1(n25805), .B2(n25756), .ZN(
        n7367) );
  OAI22_X1 U19580 ( .A1(n25764), .A2(n21020), .B1(n25808), .B2(n25756), .ZN(
        n7368) );
  OAI22_X1 U19581 ( .A1(n25764), .A2(n21019), .B1(n25811), .B2(n25756), .ZN(
        n7369) );
  OAI22_X1 U19582 ( .A1(n25764), .A2(n21018), .B1(n25814), .B2(n25756), .ZN(
        n7370) );
  OAI22_X1 U19583 ( .A1(n25765), .A2(n21017), .B1(n25817), .B2(n25757), .ZN(
        n7371) );
  OAI22_X1 U19584 ( .A1(n25765), .A2(n21016), .B1(n25820), .B2(n25757), .ZN(
        n7372) );
  OAI22_X1 U19585 ( .A1(n25765), .A2(n21015), .B1(n25823), .B2(n25757), .ZN(
        n7373) );
  OAI22_X1 U19586 ( .A1(n25765), .A2(n21014), .B1(n25826), .B2(n25757), .ZN(
        n7374) );
  OAI22_X1 U19587 ( .A1(n25765), .A2(n21013), .B1(n25829), .B2(n25757), .ZN(
        n7375) );
  OAI22_X1 U19588 ( .A1(n25765), .A2(n21012), .B1(n25832), .B2(n25757), .ZN(
        n7376) );
  OAI22_X1 U19589 ( .A1(n25765), .A2(n21011), .B1(n25835), .B2(n25757), .ZN(
        n7377) );
  OAI22_X1 U19590 ( .A1(n25765), .A2(n21010), .B1(n25838), .B2(n25757), .ZN(
        n7378) );
  OAI22_X1 U19591 ( .A1(n25765), .A2(n21009), .B1(n25841), .B2(n25757), .ZN(
        n7379) );
  OAI22_X1 U19592 ( .A1(n25765), .A2(n21008), .B1(n25844), .B2(n25757), .ZN(
        n7380) );
  OAI22_X1 U19593 ( .A1(n25765), .A2(n21007), .B1(n25847), .B2(n25757), .ZN(
        n7381) );
  OAI22_X1 U19594 ( .A1(n25765), .A2(n21006), .B1(n25850), .B2(n25757), .ZN(
        n7382) );
  OAI22_X1 U19595 ( .A1(n25765), .A2(n21005), .B1(n25853), .B2(n25758), .ZN(
        n7383) );
  OAI22_X1 U19596 ( .A1(n25766), .A2(n21004), .B1(n25856), .B2(n25758), .ZN(
        n7384) );
  OAI22_X1 U19597 ( .A1(n25766), .A2(n21003), .B1(n25859), .B2(n25758), .ZN(
        n7385) );
  OAI22_X1 U19598 ( .A1(n25766), .A2(n21002), .B1(n25862), .B2(n25758), .ZN(
        n7386) );
  OAI22_X1 U19599 ( .A1(n25766), .A2(n21001), .B1(n25865), .B2(n25758), .ZN(
        n7387) );
  OAI22_X1 U19600 ( .A1(n25766), .A2(n21000), .B1(n25868), .B2(n25758), .ZN(
        n7388) );
  OAI22_X1 U19601 ( .A1(n25766), .A2(n20999), .B1(n25871), .B2(n25758), .ZN(
        n7389) );
  OAI22_X1 U19602 ( .A1(n25766), .A2(n20998), .B1(n25874), .B2(n25758), .ZN(
        n7390) );
  OAI22_X1 U19603 ( .A1(n25766), .A2(n20997), .B1(n25877), .B2(n25758), .ZN(
        n7391) );
  OAI22_X1 U19604 ( .A1(n25766), .A2(n20996), .B1(n25880), .B2(n25758), .ZN(
        n7392) );
  OAI22_X1 U19605 ( .A1(n25766), .A2(n20995), .B1(n25883), .B2(n25758), .ZN(
        n7393) );
  OAI22_X1 U19606 ( .A1(n25766), .A2(n20994), .B1(n25886), .B2(n25758), .ZN(
        n7394) );
  OAI22_X1 U19607 ( .A1(n25766), .A2(n20993), .B1(n25889), .B2(n25759), .ZN(
        n7395) );
  OAI22_X1 U19608 ( .A1(n25766), .A2(n20992), .B1(n25892), .B2(n25759), .ZN(
        n7396) );
  OAI22_X1 U19609 ( .A1(n25767), .A2(n20991), .B1(n25895), .B2(n25759), .ZN(
        n7397) );
  OAI22_X1 U19610 ( .A1(n25767), .A2(n20990), .B1(n25898), .B2(n25759), .ZN(
        n7398) );
  OAI22_X1 U19611 ( .A1(n25767), .A2(n20989), .B1(n25901), .B2(n25759), .ZN(
        n7399) );
  OAI22_X1 U19612 ( .A1(n25767), .A2(n20988), .B1(n25904), .B2(n25759), .ZN(
        n7400) );
  OAI22_X1 U19613 ( .A1(n25767), .A2(n20987), .B1(n25907), .B2(n25759), .ZN(
        n7401) );
  OAI22_X1 U19614 ( .A1(n25767), .A2(n20986), .B1(n25910), .B2(n25759), .ZN(
        n7402) );
  OAI22_X1 U19615 ( .A1(n25767), .A2(n20985), .B1(n25913), .B2(n25759), .ZN(
        n7403) );
  OAI22_X1 U19616 ( .A1(n25767), .A2(n20984), .B1(n25916), .B2(n25759), .ZN(
        n7404) );
  OAI22_X1 U19617 ( .A1(n25767), .A2(n20983), .B1(n25919), .B2(n25759), .ZN(
        n7405) );
  OAI22_X1 U19618 ( .A1(n25767), .A2(n20982), .B1(n25922), .B2(n25759), .ZN(
        n7406) );
  OAI22_X1 U19619 ( .A1(n25767), .A2(n20981), .B1(n25925), .B2(n25760), .ZN(
        n7407) );
  OAI22_X1 U19620 ( .A1(n25767), .A2(n20980), .B1(n25928), .B2(n25760), .ZN(
        n7408) );
  OAI22_X1 U19621 ( .A1(n25767), .A2(n20979), .B1(n25931), .B2(n25760), .ZN(
        n7409) );
  OAI22_X1 U19622 ( .A1(n25768), .A2(n20978), .B1(n25934), .B2(n25760), .ZN(
        n7410) );
  OAI22_X1 U19623 ( .A1(n25768), .A2(n20977), .B1(n25937), .B2(n25760), .ZN(
        n7411) );
  OAI22_X1 U19624 ( .A1(n25768), .A2(n20976), .B1(n25940), .B2(n25760), .ZN(
        n7412) );
  OAI22_X1 U19625 ( .A1(n25768), .A2(n20975), .B1(n25943), .B2(n25760), .ZN(
        n7413) );
  OAI22_X1 U19626 ( .A1(n25768), .A2(n20974), .B1(n25946), .B2(n25760), .ZN(
        n7414) );
  OAI22_X1 U19627 ( .A1(n25768), .A2(n20973), .B1(n25949), .B2(n25760), .ZN(
        n7415) );
  OAI22_X1 U19628 ( .A1(n25768), .A2(n20972), .B1(n25952), .B2(n25760), .ZN(
        n7416) );
  OAI22_X1 U19629 ( .A1(n25768), .A2(n20971), .B1(n25955), .B2(n25760), .ZN(
        n7417) );
  OAI22_X1 U19630 ( .A1(n25768), .A2(n20970), .B1(n25958), .B2(n25760), .ZN(
        n7418) );
  OAI22_X1 U19631 ( .A1(n25533), .A2(n20773), .B1(n25782), .B2(n25525), .ZN(
        n6207) );
  OAI22_X1 U19632 ( .A1(n25533), .A2(n20772), .B1(n25785), .B2(n25525), .ZN(
        n6208) );
  OAI22_X1 U19633 ( .A1(n25533), .A2(n20771), .B1(n25788), .B2(n25525), .ZN(
        n6209) );
  OAI22_X1 U19634 ( .A1(n25533), .A2(n20770), .B1(n25791), .B2(n25525), .ZN(
        n6210) );
  OAI22_X1 U19635 ( .A1(n25533), .A2(n20769), .B1(n25794), .B2(n25525), .ZN(
        n6211) );
  OAI22_X1 U19636 ( .A1(n25533), .A2(n20768), .B1(n25797), .B2(n25525), .ZN(
        n6212) );
  OAI22_X1 U19637 ( .A1(n25533), .A2(n20767), .B1(n25800), .B2(n25525), .ZN(
        n6213) );
  OAI22_X1 U19638 ( .A1(n25533), .A2(n20766), .B1(n25803), .B2(n25525), .ZN(
        n6214) );
  OAI22_X1 U19639 ( .A1(n25533), .A2(n20765), .B1(n25806), .B2(n25525), .ZN(
        n6215) );
  OAI22_X1 U19640 ( .A1(n25533), .A2(n20764), .B1(n25809), .B2(n25525), .ZN(
        n6216) );
  OAI22_X1 U19641 ( .A1(n25533), .A2(n20763), .B1(n25812), .B2(n25525), .ZN(
        n6217) );
  OAI22_X1 U19642 ( .A1(n25533), .A2(n20762), .B1(n25815), .B2(n25525), .ZN(
        n6218) );
  OAI22_X1 U19643 ( .A1(n25534), .A2(n20761), .B1(n25818), .B2(n25526), .ZN(
        n6219) );
  OAI22_X1 U19644 ( .A1(n25534), .A2(n20760), .B1(n25821), .B2(n25526), .ZN(
        n6220) );
  OAI22_X1 U19645 ( .A1(n25534), .A2(n20759), .B1(n25824), .B2(n25526), .ZN(
        n6221) );
  OAI22_X1 U19646 ( .A1(n25534), .A2(n20758), .B1(n25827), .B2(n25526), .ZN(
        n6222) );
  OAI22_X1 U19647 ( .A1(n25534), .A2(n20757), .B1(n25830), .B2(n25526), .ZN(
        n6223) );
  OAI22_X1 U19648 ( .A1(n25534), .A2(n20756), .B1(n25833), .B2(n25526), .ZN(
        n6224) );
  OAI22_X1 U19649 ( .A1(n25534), .A2(n20755), .B1(n25836), .B2(n25526), .ZN(
        n6225) );
  OAI22_X1 U19650 ( .A1(n25534), .A2(n20754), .B1(n25839), .B2(n25526), .ZN(
        n6226) );
  OAI22_X1 U19651 ( .A1(n25534), .A2(n20753), .B1(n25842), .B2(n25526), .ZN(
        n6227) );
  OAI22_X1 U19652 ( .A1(n25534), .A2(n20752), .B1(n25845), .B2(n25526), .ZN(
        n6228) );
  OAI22_X1 U19653 ( .A1(n25534), .A2(n20751), .B1(n25848), .B2(n25526), .ZN(
        n6229) );
  OAI22_X1 U19654 ( .A1(n25534), .A2(n20750), .B1(n25851), .B2(n25526), .ZN(
        n6230) );
  OAI22_X1 U19655 ( .A1(n25534), .A2(n20749), .B1(n25854), .B2(n25527), .ZN(
        n6231) );
  OAI22_X1 U19656 ( .A1(n25535), .A2(n20748), .B1(n25857), .B2(n25527), .ZN(
        n6232) );
  OAI22_X1 U19657 ( .A1(n25535), .A2(n20747), .B1(n25860), .B2(n25527), .ZN(
        n6233) );
  OAI22_X1 U19658 ( .A1(n25535), .A2(n20746), .B1(n25863), .B2(n25527), .ZN(
        n6234) );
  OAI22_X1 U19659 ( .A1(n25535), .A2(n20745), .B1(n25866), .B2(n25527), .ZN(
        n6235) );
  OAI22_X1 U19660 ( .A1(n25535), .A2(n20744), .B1(n25869), .B2(n25527), .ZN(
        n6236) );
  OAI22_X1 U19661 ( .A1(n25535), .A2(n20743), .B1(n25872), .B2(n25527), .ZN(
        n6237) );
  OAI22_X1 U19662 ( .A1(n25535), .A2(n20742), .B1(n25875), .B2(n25527), .ZN(
        n6238) );
  OAI22_X1 U19663 ( .A1(n25535), .A2(n20741), .B1(n25878), .B2(n25527), .ZN(
        n6239) );
  OAI22_X1 U19664 ( .A1(n25535), .A2(n20740), .B1(n25881), .B2(n25527), .ZN(
        n6240) );
  OAI22_X1 U19665 ( .A1(n25535), .A2(n20739), .B1(n25884), .B2(n25527), .ZN(
        n6241) );
  OAI22_X1 U19666 ( .A1(n25535), .A2(n20738), .B1(n25887), .B2(n25527), .ZN(
        n6242) );
  OAI22_X1 U19667 ( .A1(n25535), .A2(n20737), .B1(n25890), .B2(n25528), .ZN(
        n6243) );
  OAI22_X1 U19668 ( .A1(n25535), .A2(n20736), .B1(n25893), .B2(n25528), .ZN(
        n6244) );
  OAI22_X1 U19669 ( .A1(n25536), .A2(n20735), .B1(n25896), .B2(n25528), .ZN(
        n6245) );
  OAI22_X1 U19670 ( .A1(n25536), .A2(n20734), .B1(n25899), .B2(n25528), .ZN(
        n6246) );
  OAI22_X1 U19671 ( .A1(n25536), .A2(n20733), .B1(n25902), .B2(n25528), .ZN(
        n6247) );
  OAI22_X1 U19672 ( .A1(n25536), .A2(n20732), .B1(n25905), .B2(n25528), .ZN(
        n6248) );
  OAI22_X1 U19673 ( .A1(n25536), .A2(n20731), .B1(n25908), .B2(n25528), .ZN(
        n6249) );
  OAI22_X1 U19674 ( .A1(n25536), .A2(n20730), .B1(n25911), .B2(n25528), .ZN(
        n6250) );
  OAI22_X1 U19675 ( .A1(n25536), .A2(n20729), .B1(n25914), .B2(n25528), .ZN(
        n6251) );
  OAI22_X1 U19676 ( .A1(n25536), .A2(n20728), .B1(n25917), .B2(n25528), .ZN(
        n6252) );
  OAI22_X1 U19677 ( .A1(n25536), .A2(n20727), .B1(n25920), .B2(n25528), .ZN(
        n6253) );
  OAI22_X1 U19678 ( .A1(n25536), .A2(n20726), .B1(n25923), .B2(n25528), .ZN(
        n6254) );
  OAI22_X1 U19679 ( .A1(n25536), .A2(n20725), .B1(n25926), .B2(n25529), .ZN(
        n6255) );
  OAI22_X1 U19680 ( .A1(n25536), .A2(n20724), .B1(n25929), .B2(n25529), .ZN(
        n6256) );
  OAI22_X1 U19681 ( .A1(n25536), .A2(n20723), .B1(n25932), .B2(n25529), .ZN(
        n6257) );
  OAI22_X1 U19682 ( .A1(n25537), .A2(n20722), .B1(n25935), .B2(n25529), .ZN(
        n6258) );
  OAI22_X1 U19683 ( .A1(n25537), .A2(n20721), .B1(n25938), .B2(n25529), .ZN(
        n6259) );
  OAI22_X1 U19684 ( .A1(n25537), .A2(n20720), .B1(n25941), .B2(n25529), .ZN(
        n6260) );
  OAI22_X1 U19685 ( .A1(n25537), .A2(n20719), .B1(n25944), .B2(n25529), .ZN(
        n6261) );
  OAI22_X1 U19686 ( .A1(n25537), .A2(n20718), .B1(n25947), .B2(n25529), .ZN(
        n6262) );
  OAI22_X1 U19687 ( .A1(n25537), .A2(n20717), .B1(n25950), .B2(n25529), .ZN(
        n6263) );
  OAI22_X1 U19688 ( .A1(n25537), .A2(n20716), .B1(n25953), .B2(n25529), .ZN(
        n6264) );
  OAI22_X1 U19689 ( .A1(n25537), .A2(n20715), .B1(n25956), .B2(n25529), .ZN(
        n6265) );
  OAI22_X1 U19690 ( .A1(n25537), .A2(n20714), .B1(n25959), .B2(n25529), .ZN(
        n6266) );
  OAI22_X1 U19691 ( .A1(n25726), .A2(n20709), .B1(n25781), .B2(n25718), .ZN(
        n7167) );
  OAI22_X1 U19692 ( .A1(n25726), .A2(n20708), .B1(n25784), .B2(n25718), .ZN(
        n7168) );
  OAI22_X1 U19693 ( .A1(n25726), .A2(n20707), .B1(n25787), .B2(n25718), .ZN(
        n7169) );
  OAI22_X1 U19694 ( .A1(n25726), .A2(n20706), .B1(n25790), .B2(n25718), .ZN(
        n7170) );
  OAI22_X1 U19695 ( .A1(n25726), .A2(n20705), .B1(n25793), .B2(n25718), .ZN(
        n7171) );
  OAI22_X1 U19696 ( .A1(n25726), .A2(n20704), .B1(n25796), .B2(n25718), .ZN(
        n7172) );
  OAI22_X1 U19697 ( .A1(n25726), .A2(n20703), .B1(n25799), .B2(n25718), .ZN(
        n7173) );
  OAI22_X1 U19698 ( .A1(n25726), .A2(n20702), .B1(n25802), .B2(n25718), .ZN(
        n7174) );
  OAI22_X1 U19699 ( .A1(n25726), .A2(n20701), .B1(n25805), .B2(n25718), .ZN(
        n7175) );
  OAI22_X1 U19700 ( .A1(n25726), .A2(n20700), .B1(n25808), .B2(n25718), .ZN(
        n7176) );
  OAI22_X1 U19701 ( .A1(n25726), .A2(n20699), .B1(n25811), .B2(n25718), .ZN(
        n7177) );
  OAI22_X1 U19702 ( .A1(n25726), .A2(n20698), .B1(n25814), .B2(n25718), .ZN(
        n7178) );
  OAI22_X1 U19703 ( .A1(n25727), .A2(n20697), .B1(n25817), .B2(n25719), .ZN(
        n7179) );
  OAI22_X1 U19704 ( .A1(n25727), .A2(n20696), .B1(n25820), .B2(n25719), .ZN(
        n7180) );
  OAI22_X1 U19705 ( .A1(n25727), .A2(n20695), .B1(n25823), .B2(n25719), .ZN(
        n7181) );
  OAI22_X1 U19706 ( .A1(n25727), .A2(n20694), .B1(n25826), .B2(n25719), .ZN(
        n7182) );
  OAI22_X1 U19707 ( .A1(n25727), .A2(n20693), .B1(n25829), .B2(n25719), .ZN(
        n7183) );
  OAI22_X1 U19708 ( .A1(n25727), .A2(n20692), .B1(n25832), .B2(n25719), .ZN(
        n7184) );
  OAI22_X1 U19709 ( .A1(n25727), .A2(n20691), .B1(n25835), .B2(n25719), .ZN(
        n7185) );
  OAI22_X1 U19710 ( .A1(n25727), .A2(n20690), .B1(n25838), .B2(n25719), .ZN(
        n7186) );
  OAI22_X1 U19711 ( .A1(n25727), .A2(n20689), .B1(n25841), .B2(n25719), .ZN(
        n7187) );
  OAI22_X1 U19712 ( .A1(n25727), .A2(n20688), .B1(n25844), .B2(n25719), .ZN(
        n7188) );
  OAI22_X1 U19713 ( .A1(n25727), .A2(n20687), .B1(n25847), .B2(n25719), .ZN(
        n7189) );
  OAI22_X1 U19714 ( .A1(n25727), .A2(n20686), .B1(n25850), .B2(n25719), .ZN(
        n7190) );
  OAI22_X1 U19715 ( .A1(n25727), .A2(n20685), .B1(n25853), .B2(n25720), .ZN(
        n7191) );
  OAI22_X1 U19716 ( .A1(n25728), .A2(n20684), .B1(n25856), .B2(n25720), .ZN(
        n7192) );
  OAI22_X1 U19717 ( .A1(n25728), .A2(n20683), .B1(n25859), .B2(n25720), .ZN(
        n7193) );
  OAI22_X1 U19718 ( .A1(n25728), .A2(n20682), .B1(n25862), .B2(n25720), .ZN(
        n7194) );
  OAI22_X1 U19719 ( .A1(n25728), .A2(n20681), .B1(n25865), .B2(n25720), .ZN(
        n7195) );
  OAI22_X1 U19720 ( .A1(n25728), .A2(n20680), .B1(n25868), .B2(n25720), .ZN(
        n7196) );
  OAI22_X1 U19721 ( .A1(n25728), .A2(n20679), .B1(n25871), .B2(n25720), .ZN(
        n7197) );
  OAI22_X1 U19722 ( .A1(n25728), .A2(n20678), .B1(n25874), .B2(n25720), .ZN(
        n7198) );
  OAI22_X1 U19723 ( .A1(n25728), .A2(n20677), .B1(n25877), .B2(n25720), .ZN(
        n7199) );
  OAI22_X1 U19724 ( .A1(n25728), .A2(n20676), .B1(n25880), .B2(n25720), .ZN(
        n7200) );
  OAI22_X1 U19725 ( .A1(n25728), .A2(n20675), .B1(n25883), .B2(n25720), .ZN(
        n7201) );
  OAI22_X1 U19726 ( .A1(n25728), .A2(n20674), .B1(n25886), .B2(n25720), .ZN(
        n7202) );
  OAI22_X1 U19727 ( .A1(n25728), .A2(n20673), .B1(n25889), .B2(n25721), .ZN(
        n7203) );
  OAI22_X1 U19728 ( .A1(n25728), .A2(n20672), .B1(n25892), .B2(n25721), .ZN(
        n7204) );
  OAI22_X1 U19729 ( .A1(n25729), .A2(n20671), .B1(n25895), .B2(n25721), .ZN(
        n7205) );
  OAI22_X1 U19730 ( .A1(n25729), .A2(n20670), .B1(n25898), .B2(n25721), .ZN(
        n7206) );
  OAI22_X1 U19731 ( .A1(n25729), .A2(n20669), .B1(n25901), .B2(n25721), .ZN(
        n7207) );
  OAI22_X1 U19732 ( .A1(n25729), .A2(n20668), .B1(n25904), .B2(n25721), .ZN(
        n7208) );
  OAI22_X1 U19733 ( .A1(n25729), .A2(n20667), .B1(n25907), .B2(n25721), .ZN(
        n7209) );
  OAI22_X1 U19734 ( .A1(n25729), .A2(n20666), .B1(n25910), .B2(n25721), .ZN(
        n7210) );
  OAI22_X1 U19735 ( .A1(n25729), .A2(n20665), .B1(n25913), .B2(n25721), .ZN(
        n7211) );
  OAI22_X1 U19736 ( .A1(n25729), .A2(n20664), .B1(n25916), .B2(n25721), .ZN(
        n7212) );
  OAI22_X1 U19737 ( .A1(n25729), .A2(n20663), .B1(n25919), .B2(n25721), .ZN(
        n7213) );
  OAI22_X1 U19738 ( .A1(n25729), .A2(n20662), .B1(n25922), .B2(n25721), .ZN(
        n7214) );
  OAI22_X1 U19739 ( .A1(n25729), .A2(n20661), .B1(n25925), .B2(n25722), .ZN(
        n7215) );
  OAI22_X1 U19740 ( .A1(n25729), .A2(n20660), .B1(n25928), .B2(n25722), .ZN(
        n7216) );
  OAI22_X1 U19741 ( .A1(n25729), .A2(n20659), .B1(n25931), .B2(n25722), .ZN(
        n7217) );
  OAI22_X1 U19742 ( .A1(n25730), .A2(n20658), .B1(n25934), .B2(n25722), .ZN(
        n7218) );
  OAI22_X1 U19743 ( .A1(n25730), .A2(n20657), .B1(n25937), .B2(n25722), .ZN(
        n7219) );
  OAI22_X1 U19744 ( .A1(n25730), .A2(n20656), .B1(n25940), .B2(n25722), .ZN(
        n7220) );
  OAI22_X1 U19745 ( .A1(n25730), .A2(n20655), .B1(n25943), .B2(n25722), .ZN(
        n7221) );
  OAI22_X1 U19746 ( .A1(n25730), .A2(n20654), .B1(n25946), .B2(n25722), .ZN(
        n7222) );
  OAI22_X1 U19747 ( .A1(n25730), .A2(n20653), .B1(n25949), .B2(n25722), .ZN(
        n7223) );
  OAI22_X1 U19748 ( .A1(n25730), .A2(n20652), .B1(n25952), .B2(n25722), .ZN(
        n7224) );
  OAI22_X1 U19749 ( .A1(n25730), .A2(n20651), .B1(n25955), .B2(n25722), .ZN(
        n7225) );
  OAI22_X1 U19750 ( .A1(n25730), .A2(n20650), .B1(n25958), .B2(n25722), .ZN(
        n7226) );
  OAI22_X1 U19751 ( .A1(n25623), .A2(n20461), .B1(n25782), .B2(n25615), .ZN(
        n6655) );
  OAI22_X1 U19752 ( .A1(n25623), .A2(n20460), .B1(n25785), .B2(n25615), .ZN(
        n6656) );
  OAI22_X1 U19753 ( .A1(n25623), .A2(n20459), .B1(n25788), .B2(n25615), .ZN(
        n6657) );
  OAI22_X1 U19754 ( .A1(n25623), .A2(n20458), .B1(n25791), .B2(n25615), .ZN(
        n6658) );
  OAI22_X1 U19755 ( .A1(n25623), .A2(n20457), .B1(n25794), .B2(n25615), .ZN(
        n6659) );
  OAI22_X1 U19756 ( .A1(n25623), .A2(n20456), .B1(n25797), .B2(n25615), .ZN(
        n6660) );
  OAI22_X1 U19757 ( .A1(n25623), .A2(n20455), .B1(n25800), .B2(n25615), .ZN(
        n6661) );
  OAI22_X1 U19758 ( .A1(n25623), .A2(n20454), .B1(n25803), .B2(n25615), .ZN(
        n6662) );
  OAI22_X1 U19759 ( .A1(n25623), .A2(n20453), .B1(n25806), .B2(n25615), .ZN(
        n6663) );
  OAI22_X1 U19760 ( .A1(n25623), .A2(n20452), .B1(n25809), .B2(n25615), .ZN(
        n6664) );
  OAI22_X1 U19761 ( .A1(n25623), .A2(n20451), .B1(n25812), .B2(n25615), .ZN(
        n6665) );
  OAI22_X1 U19762 ( .A1(n25623), .A2(n20450), .B1(n25815), .B2(n25615), .ZN(
        n6666) );
  OAI22_X1 U19763 ( .A1(n25624), .A2(n20449), .B1(n25818), .B2(n25616), .ZN(
        n6667) );
  OAI22_X1 U19764 ( .A1(n25624), .A2(n20448), .B1(n25821), .B2(n25616), .ZN(
        n6668) );
  OAI22_X1 U19765 ( .A1(n25624), .A2(n20447), .B1(n25824), .B2(n25616), .ZN(
        n6669) );
  OAI22_X1 U19766 ( .A1(n25624), .A2(n20446), .B1(n25827), .B2(n25616), .ZN(
        n6670) );
  OAI22_X1 U19767 ( .A1(n25624), .A2(n20445), .B1(n25830), .B2(n25616), .ZN(
        n6671) );
  OAI22_X1 U19768 ( .A1(n25624), .A2(n20444), .B1(n25833), .B2(n25616), .ZN(
        n6672) );
  OAI22_X1 U19769 ( .A1(n25624), .A2(n20443), .B1(n25836), .B2(n25616), .ZN(
        n6673) );
  OAI22_X1 U19770 ( .A1(n25624), .A2(n20442), .B1(n25839), .B2(n25616), .ZN(
        n6674) );
  OAI22_X1 U19771 ( .A1(n25624), .A2(n20441), .B1(n25842), .B2(n25616), .ZN(
        n6675) );
  OAI22_X1 U19772 ( .A1(n25624), .A2(n20440), .B1(n25845), .B2(n25616), .ZN(
        n6676) );
  OAI22_X1 U19773 ( .A1(n25624), .A2(n20439), .B1(n25848), .B2(n25616), .ZN(
        n6677) );
  OAI22_X1 U19774 ( .A1(n25624), .A2(n20438), .B1(n25851), .B2(n25616), .ZN(
        n6678) );
  OAI22_X1 U19775 ( .A1(n25624), .A2(n20437), .B1(n25854), .B2(n25617), .ZN(
        n6679) );
  OAI22_X1 U19776 ( .A1(n25625), .A2(n20436), .B1(n25857), .B2(n25617), .ZN(
        n6680) );
  OAI22_X1 U19777 ( .A1(n25625), .A2(n20435), .B1(n25860), .B2(n25617), .ZN(
        n6681) );
  OAI22_X1 U19778 ( .A1(n25625), .A2(n20434), .B1(n25863), .B2(n25617), .ZN(
        n6682) );
  OAI22_X1 U19779 ( .A1(n25625), .A2(n20433), .B1(n25866), .B2(n25617), .ZN(
        n6683) );
  OAI22_X1 U19780 ( .A1(n25625), .A2(n20432), .B1(n25869), .B2(n25617), .ZN(
        n6684) );
  OAI22_X1 U19781 ( .A1(n25625), .A2(n20431), .B1(n25872), .B2(n25617), .ZN(
        n6685) );
  OAI22_X1 U19782 ( .A1(n25625), .A2(n20430), .B1(n25875), .B2(n25617), .ZN(
        n6686) );
  OAI22_X1 U19783 ( .A1(n25625), .A2(n20429), .B1(n25878), .B2(n25617), .ZN(
        n6687) );
  OAI22_X1 U19784 ( .A1(n25625), .A2(n20428), .B1(n25881), .B2(n25617), .ZN(
        n6688) );
  OAI22_X1 U19785 ( .A1(n25625), .A2(n20427), .B1(n25884), .B2(n25617), .ZN(
        n6689) );
  OAI22_X1 U19786 ( .A1(n25625), .A2(n20426), .B1(n25887), .B2(n25617), .ZN(
        n6690) );
  OAI22_X1 U19787 ( .A1(n25625), .A2(n20425), .B1(n25890), .B2(n25618), .ZN(
        n6691) );
  OAI22_X1 U19788 ( .A1(n25625), .A2(n20424), .B1(n25893), .B2(n25618), .ZN(
        n6692) );
  OAI22_X1 U19789 ( .A1(n25626), .A2(n20423), .B1(n25896), .B2(n25618), .ZN(
        n6693) );
  OAI22_X1 U19790 ( .A1(n25626), .A2(n20422), .B1(n25899), .B2(n25618), .ZN(
        n6694) );
  OAI22_X1 U19791 ( .A1(n25626), .A2(n20421), .B1(n25902), .B2(n25618), .ZN(
        n6695) );
  OAI22_X1 U19792 ( .A1(n25626), .A2(n20420), .B1(n25905), .B2(n25618), .ZN(
        n6696) );
  OAI22_X1 U19793 ( .A1(n25626), .A2(n20419), .B1(n25908), .B2(n25618), .ZN(
        n6697) );
  OAI22_X1 U19794 ( .A1(n25626), .A2(n20418), .B1(n25911), .B2(n25618), .ZN(
        n6698) );
  OAI22_X1 U19795 ( .A1(n25626), .A2(n20417), .B1(n25914), .B2(n25618), .ZN(
        n6699) );
  OAI22_X1 U19796 ( .A1(n25626), .A2(n20416), .B1(n25917), .B2(n25618), .ZN(
        n6700) );
  OAI22_X1 U19797 ( .A1(n25626), .A2(n20415), .B1(n25920), .B2(n25618), .ZN(
        n6701) );
  OAI22_X1 U19798 ( .A1(n25626), .A2(n20414), .B1(n25923), .B2(n25618), .ZN(
        n6702) );
  OAI22_X1 U19799 ( .A1(n25626), .A2(n20413), .B1(n25926), .B2(n25619), .ZN(
        n6703) );
  OAI22_X1 U19800 ( .A1(n25626), .A2(n20412), .B1(n25929), .B2(n25619), .ZN(
        n6704) );
  OAI22_X1 U19801 ( .A1(n25626), .A2(n20411), .B1(n25932), .B2(n25619), .ZN(
        n6705) );
  OAI22_X1 U19802 ( .A1(n25627), .A2(n20410), .B1(n25935), .B2(n25619), .ZN(
        n6706) );
  OAI22_X1 U19803 ( .A1(n25627), .A2(n20409), .B1(n25938), .B2(n25619), .ZN(
        n6707) );
  OAI22_X1 U19804 ( .A1(n25627), .A2(n20408), .B1(n25941), .B2(n25619), .ZN(
        n6708) );
  OAI22_X1 U19805 ( .A1(n25627), .A2(n20407), .B1(n25944), .B2(n25619), .ZN(
        n6709) );
  OAI22_X1 U19806 ( .A1(n25627), .A2(n20406), .B1(n25947), .B2(n25619), .ZN(
        n6710) );
  OAI22_X1 U19807 ( .A1(n25627), .A2(n20405), .B1(n25950), .B2(n25619), .ZN(
        n6711) );
  OAI22_X1 U19808 ( .A1(n25627), .A2(n20404), .B1(n25953), .B2(n25619), .ZN(
        n6712) );
  OAI22_X1 U19809 ( .A1(n25627), .A2(n20403), .B1(n25956), .B2(n25619), .ZN(
        n6713) );
  OAI22_X1 U19810 ( .A1(n25627), .A2(n20402), .B1(n25959), .B2(n25619), .ZN(
        n6714) );
  OAI22_X1 U19811 ( .A1(n25546), .A2(n20397), .B1(n25782), .B2(n25538), .ZN(
        n6271) );
  OAI22_X1 U19812 ( .A1(n25546), .A2(n20396), .B1(n25785), .B2(n25538), .ZN(
        n6272) );
  OAI22_X1 U19813 ( .A1(n25546), .A2(n20395), .B1(n25788), .B2(n25538), .ZN(
        n6273) );
  OAI22_X1 U19814 ( .A1(n25546), .A2(n20394), .B1(n25791), .B2(n25538), .ZN(
        n6274) );
  OAI22_X1 U19815 ( .A1(n25546), .A2(n20393), .B1(n25794), .B2(n25538), .ZN(
        n6275) );
  OAI22_X1 U19816 ( .A1(n25546), .A2(n20392), .B1(n25797), .B2(n25538), .ZN(
        n6276) );
  OAI22_X1 U19817 ( .A1(n25546), .A2(n20391), .B1(n25800), .B2(n25538), .ZN(
        n6277) );
  OAI22_X1 U19818 ( .A1(n25546), .A2(n20390), .B1(n25803), .B2(n25538), .ZN(
        n6278) );
  OAI22_X1 U19819 ( .A1(n25546), .A2(n20389), .B1(n25806), .B2(n25538), .ZN(
        n6279) );
  OAI22_X1 U19820 ( .A1(n25546), .A2(n20388), .B1(n25809), .B2(n25538), .ZN(
        n6280) );
  OAI22_X1 U19821 ( .A1(n25546), .A2(n20387), .B1(n25812), .B2(n25538), .ZN(
        n6281) );
  OAI22_X1 U19822 ( .A1(n25546), .A2(n20386), .B1(n25815), .B2(n25538), .ZN(
        n6282) );
  OAI22_X1 U19823 ( .A1(n25547), .A2(n20385), .B1(n25818), .B2(n25539), .ZN(
        n6283) );
  OAI22_X1 U19824 ( .A1(n25547), .A2(n20384), .B1(n25821), .B2(n25539), .ZN(
        n6284) );
  OAI22_X1 U19825 ( .A1(n25547), .A2(n20383), .B1(n25824), .B2(n25539), .ZN(
        n6285) );
  OAI22_X1 U19826 ( .A1(n25547), .A2(n20382), .B1(n25827), .B2(n25539), .ZN(
        n6286) );
  OAI22_X1 U19827 ( .A1(n25547), .A2(n20381), .B1(n25830), .B2(n25539), .ZN(
        n6287) );
  OAI22_X1 U19828 ( .A1(n25547), .A2(n20380), .B1(n25833), .B2(n25539), .ZN(
        n6288) );
  OAI22_X1 U19829 ( .A1(n25547), .A2(n20379), .B1(n25836), .B2(n25539), .ZN(
        n6289) );
  OAI22_X1 U19830 ( .A1(n25547), .A2(n20378), .B1(n25839), .B2(n25539), .ZN(
        n6290) );
  OAI22_X1 U19831 ( .A1(n25547), .A2(n20377), .B1(n25842), .B2(n25539), .ZN(
        n6291) );
  OAI22_X1 U19832 ( .A1(n25547), .A2(n20376), .B1(n25845), .B2(n25539), .ZN(
        n6292) );
  OAI22_X1 U19833 ( .A1(n25547), .A2(n20375), .B1(n25848), .B2(n25539), .ZN(
        n6293) );
  OAI22_X1 U19834 ( .A1(n25547), .A2(n20374), .B1(n25851), .B2(n25539), .ZN(
        n6294) );
  OAI22_X1 U19835 ( .A1(n25547), .A2(n20373), .B1(n25854), .B2(n25540), .ZN(
        n6295) );
  OAI22_X1 U19836 ( .A1(n25548), .A2(n20372), .B1(n25857), .B2(n25540), .ZN(
        n6296) );
  OAI22_X1 U19837 ( .A1(n25548), .A2(n20371), .B1(n25860), .B2(n25540), .ZN(
        n6297) );
  OAI22_X1 U19838 ( .A1(n25548), .A2(n20370), .B1(n25863), .B2(n25540), .ZN(
        n6298) );
  OAI22_X1 U19839 ( .A1(n25548), .A2(n20369), .B1(n25866), .B2(n25540), .ZN(
        n6299) );
  OAI22_X1 U19840 ( .A1(n25548), .A2(n20368), .B1(n25869), .B2(n25540), .ZN(
        n6300) );
  OAI22_X1 U19841 ( .A1(n25548), .A2(n20367), .B1(n25872), .B2(n25540), .ZN(
        n6301) );
  OAI22_X1 U19842 ( .A1(n25548), .A2(n20366), .B1(n25875), .B2(n25540), .ZN(
        n6302) );
  OAI22_X1 U19843 ( .A1(n25548), .A2(n20365), .B1(n25878), .B2(n25540), .ZN(
        n6303) );
  OAI22_X1 U19844 ( .A1(n25548), .A2(n20364), .B1(n25881), .B2(n25540), .ZN(
        n6304) );
  OAI22_X1 U19845 ( .A1(n25548), .A2(n20363), .B1(n25884), .B2(n25540), .ZN(
        n6305) );
  OAI22_X1 U19846 ( .A1(n25548), .A2(n20362), .B1(n25887), .B2(n25540), .ZN(
        n6306) );
  OAI22_X1 U19847 ( .A1(n25548), .A2(n20361), .B1(n25890), .B2(n25541), .ZN(
        n6307) );
  OAI22_X1 U19848 ( .A1(n25548), .A2(n20360), .B1(n25893), .B2(n25541), .ZN(
        n6308) );
  OAI22_X1 U19849 ( .A1(n25549), .A2(n20359), .B1(n25896), .B2(n25541), .ZN(
        n6309) );
  OAI22_X1 U19850 ( .A1(n25549), .A2(n20358), .B1(n25899), .B2(n25541), .ZN(
        n6310) );
  OAI22_X1 U19851 ( .A1(n25549), .A2(n20357), .B1(n25902), .B2(n25541), .ZN(
        n6311) );
  OAI22_X1 U19852 ( .A1(n25549), .A2(n20356), .B1(n25905), .B2(n25541), .ZN(
        n6312) );
  OAI22_X1 U19853 ( .A1(n25549), .A2(n20355), .B1(n25908), .B2(n25541), .ZN(
        n6313) );
  OAI22_X1 U19854 ( .A1(n25549), .A2(n20354), .B1(n25911), .B2(n25541), .ZN(
        n6314) );
  OAI22_X1 U19855 ( .A1(n25549), .A2(n20353), .B1(n25914), .B2(n25541), .ZN(
        n6315) );
  OAI22_X1 U19856 ( .A1(n25549), .A2(n20352), .B1(n25917), .B2(n25541), .ZN(
        n6316) );
  OAI22_X1 U19857 ( .A1(n25549), .A2(n20351), .B1(n25920), .B2(n25541), .ZN(
        n6317) );
  OAI22_X1 U19858 ( .A1(n25549), .A2(n20350), .B1(n25923), .B2(n25541), .ZN(
        n6318) );
  OAI22_X1 U19859 ( .A1(n25549), .A2(n20349), .B1(n25926), .B2(n25542), .ZN(
        n6319) );
  OAI22_X1 U19860 ( .A1(n25549), .A2(n20348), .B1(n25929), .B2(n25542), .ZN(
        n6320) );
  OAI22_X1 U19861 ( .A1(n25549), .A2(n20347), .B1(n25932), .B2(n25542), .ZN(
        n6321) );
  OAI22_X1 U19862 ( .A1(n25550), .A2(n20346), .B1(n25935), .B2(n25542), .ZN(
        n6322) );
  OAI22_X1 U19863 ( .A1(n25550), .A2(n20345), .B1(n25938), .B2(n25542), .ZN(
        n6323) );
  OAI22_X1 U19864 ( .A1(n25550), .A2(n20344), .B1(n25941), .B2(n25542), .ZN(
        n6324) );
  OAI22_X1 U19865 ( .A1(n25550), .A2(n20343), .B1(n25944), .B2(n25542), .ZN(
        n6325) );
  OAI22_X1 U19866 ( .A1(n25550), .A2(n20342), .B1(n25947), .B2(n25542), .ZN(
        n6326) );
  OAI22_X1 U19867 ( .A1(n25550), .A2(n20341), .B1(n25950), .B2(n25542), .ZN(
        n6327) );
  OAI22_X1 U19868 ( .A1(n25550), .A2(n20340), .B1(n25953), .B2(n25542), .ZN(
        n6328) );
  OAI22_X1 U19869 ( .A1(n25550), .A2(n20339), .B1(n25956), .B2(n25542), .ZN(
        n6329) );
  OAI22_X1 U19870 ( .A1(n25550), .A2(n20338), .B1(n25959), .B2(n25542), .ZN(
        n6330) );
  OAI22_X1 U19871 ( .A1(n25520), .A2(n20333), .B1(n25782), .B2(n25512), .ZN(
        n6143) );
  OAI22_X1 U19872 ( .A1(n25520), .A2(n20332), .B1(n25785), .B2(n25512), .ZN(
        n6144) );
  OAI22_X1 U19873 ( .A1(n25520), .A2(n20331), .B1(n25788), .B2(n25512), .ZN(
        n6145) );
  OAI22_X1 U19874 ( .A1(n25520), .A2(n20330), .B1(n25791), .B2(n25512), .ZN(
        n6146) );
  OAI22_X1 U19875 ( .A1(n25520), .A2(n20329), .B1(n25794), .B2(n25512), .ZN(
        n6147) );
  OAI22_X1 U19876 ( .A1(n25520), .A2(n20328), .B1(n25797), .B2(n25512), .ZN(
        n6148) );
  OAI22_X1 U19877 ( .A1(n25520), .A2(n20327), .B1(n25800), .B2(n25512), .ZN(
        n6149) );
  OAI22_X1 U19878 ( .A1(n25520), .A2(n20326), .B1(n25803), .B2(n25512), .ZN(
        n6150) );
  OAI22_X1 U19879 ( .A1(n25520), .A2(n20325), .B1(n25806), .B2(n25512), .ZN(
        n6151) );
  OAI22_X1 U19880 ( .A1(n25520), .A2(n20324), .B1(n25809), .B2(n25512), .ZN(
        n6152) );
  OAI22_X1 U19881 ( .A1(n25520), .A2(n20323), .B1(n25812), .B2(n25512), .ZN(
        n6153) );
  OAI22_X1 U19882 ( .A1(n25520), .A2(n20322), .B1(n25815), .B2(n25512), .ZN(
        n6154) );
  OAI22_X1 U19883 ( .A1(n25521), .A2(n20321), .B1(n25818), .B2(n25513), .ZN(
        n6155) );
  OAI22_X1 U19884 ( .A1(n25521), .A2(n20320), .B1(n25821), .B2(n25513), .ZN(
        n6156) );
  OAI22_X1 U19885 ( .A1(n25521), .A2(n20319), .B1(n25824), .B2(n25513), .ZN(
        n6157) );
  OAI22_X1 U19886 ( .A1(n25521), .A2(n20318), .B1(n25827), .B2(n25513), .ZN(
        n6158) );
  OAI22_X1 U19887 ( .A1(n25521), .A2(n20317), .B1(n25830), .B2(n25513), .ZN(
        n6159) );
  OAI22_X1 U19888 ( .A1(n25521), .A2(n20316), .B1(n25833), .B2(n25513), .ZN(
        n6160) );
  OAI22_X1 U19889 ( .A1(n25521), .A2(n20315), .B1(n25836), .B2(n25513), .ZN(
        n6161) );
  OAI22_X1 U19890 ( .A1(n25521), .A2(n20314), .B1(n25839), .B2(n25513), .ZN(
        n6162) );
  OAI22_X1 U19891 ( .A1(n25521), .A2(n20313), .B1(n25842), .B2(n25513), .ZN(
        n6163) );
  OAI22_X1 U19892 ( .A1(n25521), .A2(n20312), .B1(n25845), .B2(n25513), .ZN(
        n6164) );
  OAI22_X1 U19893 ( .A1(n25521), .A2(n20311), .B1(n25848), .B2(n25513), .ZN(
        n6165) );
  OAI22_X1 U19894 ( .A1(n25521), .A2(n20310), .B1(n25851), .B2(n25513), .ZN(
        n6166) );
  OAI22_X1 U19895 ( .A1(n25521), .A2(n20309), .B1(n25854), .B2(n25514), .ZN(
        n6167) );
  OAI22_X1 U19896 ( .A1(n25522), .A2(n20308), .B1(n25857), .B2(n25514), .ZN(
        n6168) );
  OAI22_X1 U19897 ( .A1(n25522), .A2(n20307), .B1(n25860), .B2(n25514), .ZN(
        n6169) );
  OAI22_X1 U19898 ( .A1(n25522), .A2(n20306), .B1(n25863), .B2(n25514), .ZN(
        n6170) );
  OAI22_X1 U19899 ( .A1(n25522), .A2(n20305), .B1(n25866), .B2(n25514), .ZN(
        n6171) );
  OAI22_X1 U19900 ( .A1(n25522), .A2(n20304), .B1(n25869), .B2(n25514), .ZN(
        n6172) );
  OAI22_X1 U19901 ( .A1(n25522), .A2(n20303), .B1(n25872), .B2(n25514), .ZN(
        n6173) );
  OAI22_X1 U19902 ( .A1(n25522), .A2(n20302), .B1(n25875), .B2(n25514), .ZN(
        n6174) );
  OAI22_X1 U19903 ( .A1(n25522), .A2(n20301), .B1(n25878), .B2(n25514), .ZN(
        n6175) );
  OAI22_X1 U19904 ( .A1(n25522), .A2(n20300), .B1(n25881), .B2(n25514), .ZN(
        n6176) );
  OAI22_X1 U19905 ( .A1(n25522), .A2(n20299), .B1(n25884), .B2(n25514), .ZN(
        n6177) );
  OAI22_X1 U19906 ( .A1(n25522), .A2(n20298), .B1(n25887), .B2(n25514), .ZN(
        n6178) );
  OAI22_X1 U19907 ( .A1(n25522), .A2(n20297), .B1(n25890), .B2(n25515), .ZN(
        n6179) );
  OAI22_X1 U19908 ( .A1(n25522), .A2(n20296), .B1(n25893), .B2(n25515), .ZN(
        n6180) );
  OAI22_X1 U19909 ( .A1(n25523), .A2(n20295), .B1(n25896), .B2(n25515), .ZN(
        n6181) );
  OAI22_X1 U19910 ( .A1(n25523), .A2(n20294), .B1(n25899), .B2(n25515), .ZN(
        n6182) );
  OAI22_X1 U19911 ( .A1(n25523), .A2(n20293), .B1(n25902), .B2(n25515), .ZN(
        n6183) );
  OAI22_X1 U19912 ( .A1(n25523), .A2(n20292), .B1(n25905), .B2(n25515), .ZN(
        n6184) );
  OAI22_X1 U19913 ( .A1(n25523), .A2(n20291), .B1(n25908), .B2(n25515), .ZN(
        n6185) );
  OAI22_X1 U19914 ( .A1(n25523), .A2(n20290), .B1(n25911), .B2(n25515), .ZN(
        n6186) );
  OAI22_X1 U19915 ( .A1(n25523), .A2(n20289), .B1(n25914), .B2(n25515), .ZN(
        n6187) );
  OAI22_X1 U19916 ( .A1(n25523), .A2(n20288), .B1(n25917), .B2(n25515), .ZN(
        n6188) );
  OAI22_X1 U19917 ( .A1(n25523), .A2(n20287), .B1(n25920), .B2(n25515), .ZN(
        n6189) );
  OAI22_X1 U19918 ( .A1(n25523), .A2(n20286), .B1(n25923), .B2(n25515), .ZN(
        n6190) );
  OAI22_X1 U19919 ( .A1(n25523), .A2(n20285), .B1(n25926), .B2(n25516), .ZN(
        n6191) );
  OAI22_X1 U19920 ( .A1(n25523), .A2(n20284), .B1(n25929), .B2(n25516), .ZN(
        n6192) );
  OAI22_X1 U19921 ( .A1(n25523), .A2(n20283), .B1(n25932), .B2(n25516), .ZN(
        n6193) );
  OAI22_X1 U19922 ( .A1(n25524), .A2(n20282), .B1(n25935), .B2(n25516), .ZN(
        n6194) );
  OAI22_X1 U19923 ( .A1(n25524), .A2(n20281), .B1(n25938), .B2(n25516), .ZN(
        n6195) );
  OAI22_X1 U19924 ( .A1(n25524), .A2(n20280), .B1(n25941), .B2(n25516), .ZN(
        n6196) );
  OAI22_X1 U19925 ( .A1(n25524), .A2(n20279), .B1(n25944), .B2(n25516), .ZN(
        n6197) );
  OAI22_X1 U19926 ( .A1(n25524), .A2(n20278), .B1(n25947), .B2(n25516), .ZN(
        n6198) );
  OAI22_X1 U19927 ( .A1(n25524), .A2(n20277), .B1(n25950), .B2(n25516), .ZN(
        n6199) );
  OAI22_X1 U19928 ( .A1(n25524), .A2(n20276), .B1(n25953), .B2(n25516), .ZN(
        n6200) );
  OAI22_X1 U19929 ( .A1(n25524), .A2(n20275), .B1(n25956), .B2(n25516), .ZN(
        n6201) );
  OAI22_X1 U19930 ( .A1(n25524), .A2(n20274), .B1(n25959), .B2(n25516), .ZN(
        n6202) );
  OAI22_X1 U19931 ( .A1(n25610), .A2(n19876), .B1(n25782), .B2(n25602), .ZN(
        n6591) );
  OAI22_X1 U19932 ( .A1(n25610), .A2(n19875), .B1(n25785), .B2(n25602), .ZN(
        n6592) );
  OAI22_X1 U19933 ( .A1(n25610), .A2(n19874), .B1(n25788), .B2(n25602), .ZN(
        n6593) );
  OAI22_X1 U19934 ( .A1(n25610), .A2(n19873), .B1(n25791), .B2(n25602), .ZN(
        n6594) );
  OAI22_X1 U19935 ( .A1(n25610), .A2(n19872), .B1(n25794), .B2(n25602), .ZN(
        n6595) );
  OAI22_X1 U19936 ( .A1(n25610), .A2(n19871), .B1(n25797), .B2(n25602), .ZN(
        n6596) );
  OAI22_X1 U19937 ( .A1(n25610), .A2(n19870), .B1(n25800), .B2(n25602), .ZN(
        n6597) );
  OAI22_X1 U19938 ( .A1(n25610), .A2(n19869), .B1(n25803), .B2(n25602), .ZN(
        n6598) );
  OAI22_X1 U19939 ( .A1(n25610), .A2(n19868), .B1(n25806), .B2(n25602), .ZN(
        n6599) );
  OAI22_X1 U19940 ( .A1(n25610), .A2(n19867), .B1(n25809), .B2(n25602), .ZN(
        n6600) );
  OAI22_X1 U19941 ( .A1(n25610), .A2(n19866), .B1(n25812), .B2(n25602), .ZN(
        n6601) );
  OAI22_X1 U19942 ( .A1(n25610), .A2(n19865), .B1(n25815), .B2(n25602), .ZN(
        n6602) );
  OAI22_X1 U19943 ( .A1(n25611), .A2(n19864), .B1(n25818), .B2(n25603), .ZN(
        n6603) );
  OAI22_X1 U19944 ( .A1(n25611), .A2(n19863), .B1(n25821), .B2(n25603), .ZN(
        n6604) );
  OAI22_X1 U19945 ( .A1(n25611), .A2(n19862), .B1(n25824), .B2(n25603), .ZN(
        n6605) );
  OAI22_X1 U19946 ( .A1(n25611), .A2(n19861), .B1(n25827), .B2(n25603), .ZN(
        n6606) );
  OAI22_X1 U19947 ( .A1(n25611), .A2(n19860), .B1(n25830), .B2(n25603), .ZN(
        n6607) );
  OAI22_X1 U19948 ( .A1(n25611), .A2(n19859), .B1(n25833), .B2(n25603), .ZN(
        n6608) );
  OAI22_X1 U19949 ( .A1(n25611), .A2(n19858), .B1(n25836), .B2(n25603), .ZN(
        n6609) );
  OAI22_X1 U19950 ( .A1(n25611), .A2(n19857), .B1(n25839), .B2(n25603), .ZN(
        n6610) );
  OAI22_X1 U19951 ( .A1(n25611), .A2(n19856), .B1(n25842), .B2(n25603), .ZN(
        n6611) );
  OAI22_X1 U19952 ( .A1(n25611), .A2(n19855), .B1(n25845), .B2(n25603), .ZN(
        n6612) );
  OAI22_X1 U19953 ( .A1(n25611), .A2(n19854), .B1(n25848), .B2(n25603), .ZN(
        n6613) );
  OAI22_X1 U19954 ( .A1(n25611), .A2(n19853), .B1(n25851), .B2(n25603), .ZN(
        n6614) );
  OAI22_X1 U19955 ( .A1(n25611), .A2(n19852), .B1(n25854), .B2(n25604), .ZN(
        n6615) );
  OAI22_X1 U19956 ( .A1(n25612), .A2(n19851), .B1(n25857), .B2(n25604), .ZN(
        n6616) );
  OAI22_X1 U19957 ( .A1(n25612), .A2(n19850), .B1(n25860), .B2(n25604), .ZN(
        n6617) );
  OAI22_X1 U19958 ( .A1(n25612), .A2(n19849), .B1(n25863), .B2(n25604), .ZN(
        n6618) );
  OAI22_X1 U19959 ( .A1(n25612), .A2(n19848), .B1(n25866), .B2(n25604), .ZN(
        n6619) );
  OAI22_X1 U19960 ( .A1(n25612), .A2(n19847), .B1(n25869), .B2(n25604), .ZN(
        n6620) );
  OAI22_X1 U19961 ( .A1(n25612), .A2(n19846), .B1(n25872), .B2(n25604), .ZN(
        n6621) );
  OAI22_X1 U19962 ( .A1(n25612), .A2(n19845), .B1(n25875), .B2(n25604), .ZN(
        n6622) );
  OAI22_X1 U19963 ( .A1(n25612), .A2(n19844), .B1(n25878), .B2(n25604), .ZN(
        n6623) );
  OAI22_X1 U19964 ( .A1(n25612), .A2(n19843), .B1(n25881), .B2(n25604), .ZN(
        n6624) );
  OAI22_X1 U19965 ( .A1(n25612), .A2(n19842), .B1(n25884), .B2(n25604), .ZN(
        n6625) );
  OAI22_X1 U19966 ( .A1(n25612), .A2(n19841), .B1(n25887), .B2(n25604), .ZN(
        n6626) );
  OAI22_X1 U19967 ( .A1(n25612), .A2(n19840), .B1(n25890), .B2(n25605), .ZN(
        n6627) );
  OAI22_X1 U19968 ( .A1(n25612), .A2(n19839), .B1(n25893), .B2(n25605), .ZN(
        n6628) );
  OAI22_X1 U19969 ( .A1(n25613), .A2(n19838), .B1(n25896), .B2(n25605), .ZN(
        n6629) );
  OAI22_X1 U19970 ( .A1(n25613), .A2(n19837), .B1(n25899), .B2(n25605), .ZN(
        n6630) );
  OAI22_X1 U19971 ( .A1(n25613), .A2(n19836), .B1(n25902), .B2(n25605), .ZN(
        n6631) );
  OAI22_X1 U19972 ( .A1(n25613), .A2(n19835), .B1(n25905), .B2(n25605), .ZN(
        n6632) );
  OAI22_X1 U19973 ( .A1(n25613), .A2(n19834), .B1(n25908), .B2(n25605), .ZN(
        n6633) );
  OAI22_X1 U19974 ( .A1(n25613), .A2(n19833), .B1(n25911), .B2(n25605), .ZN(
        n6634) );
  OAI22_X1 U19975 ( .A1(n25613), .A2(n19832), .B1(n25914), .B2(n25605), .ZN(
        n6635) );
  OAI22_X1 U19976 ( .A1(n25613), .A2(n19831), .B1(n25917), .B2(n25605), .ZN(
        n6636) );
  OAI22_X1 U19977 ( .A1(n25613), .A2(n19830), .B1(n25920), .B2(n25605), .ZN(
        n6637) );
  OAI22_X1 U19978 ( .A1(n25613), .A2(n19829), .B1(n25923), .B2(n25605), .ZN(
        n6638) );
  OAI22_X1 U19979 ( .A1(n25613), .A2(n19828), .B1(n25926), .B2(n25606), .ZN(
        n6639) );
  OAI22_X1 U19980 ( .A1(n25613), .A2(n19827), .B1(n25929), .B2(n25606), .ZN(
        n6640) );
  OAI22_X1 U19981 ( .A1(n25613), .A2(n19826), .B1(n25932), .B2(n25606), .ZN(
        n6641) );
  OAI22_X1 U19982 ( .A1(n25614), .A2(n19825), .B1(n25935), .B2(n25606), .ZN(
        n6642) );
  OAI22_X1 U19983 ( .A1(n25614), .A2(n19824), .B1(n25938), .B2(n25606), .ZN(
        n6643) );
  OAI22_X1 U19984 ( .A1(n25614), .A2(n19823), .B1(n25941), .B2(n25606), .ZN(
        n6644) );
  OAI22_X1 U19985 ( .A1(n25614), .A2(n19822), .B1(n25944), .B2(n25606), .ZN(
        n6645) );
  OAI22_X1 U19986 ( .A1(n25614), .A2(n19821), .B1(n25947), .B2(n25606), .ZN(
        n6646) );
  OAI22_X1 U19987 ( .A1(n25614), .A2(n19820), .B1(n25950), .B2(n25606), .ZN(
        n6647) );
  OAI22_X1 U19988 ( .A1(n25614), .A2(n19819), .B1(n25953), .B2(n25606), .ZN(
        n6648) );
  OAI22_X1 U19989 ( .A1(n25614), .A2(n19818), .B1(n25956), .B2(n25606), .ZN(
        n6649) );
  OAI22_X1 U19990 ( .A1(n25614), .A2(n19817), .B1(n25959), .B2(n25606), .ZN(
        n6650) );
  OAI22_X1 U19991 ( .A1(n25662), .A2(n19812), .B1(n25781), .B2(n25654), .ZN(
        n6847) );
  OAI22_X1 U19992 ( .A1(n25662), .A2(n19811), .B1(n25784), .B2(n25654), .ZN(
        n6848) );
  OAI22_X1 U19993 ( .A1(n25662), .A2(n19810), .B1(n25787), .B2(n25654), .ZN(
        n6849) );
  OAI22_X1 U19994 ( .A1(n25662), .A2(n19809), .B1(n25790), .B2(n25654), .ZN(
        n6850) );
  OAI22_X1 U19995 ( .A1(n25662), .A2(n19808), .B1(n25793), .B2(n25654), .ZN(
        n6851) );
  OAI22_X1 U19996 ( .A1(n25662), .A2(n19807), .B1(n25796), .B2(n25654), .ZN(
        n6852) );
  OAI22_X1 U19997 ( .A1(n25662), .A2(n19806), .B1(n25799), .B2(n25654), .ZN(
        n6853) );
  OAI22_X1 U19998 ( .A1(n25662), .A2(n19805), .B1(n25802), .B2(n25654), .ZN(
        n6854) );
  OAI22_X1 U19999 ( .A1(n25662), .A2(n19804), .B1(n25805), .B2(n25654), .ZN(
        n6855) );
  OAI22_X1 U20000 ( .A1(n25662), .A2(n19803), .B1(n25808), .B2(n25654), .ZN(
        n6856) );
  OAI22_X1 U20001 ( .A1(n25662), .A2(n19802), .B1(n25811), .B2(n25654), .ZN(
        n6857) );
  OAI22_X1 U20002 ( .A1(n25662), .A2(n19801), .B1(n25814), .B2(n25654), .ZN(
        n6858) );
  OAI22_X1 U20003 ( .A1(n25663), .A2(n19800), .B1(n25817), .B2(n25655), .ZN(
        n6859) );
  OAI22_X1 U20004 ( .A1(n25663), .A2(n19799), .B1(n25820), .B2(n25655), .ZN(
        n6860) );
  OAI22_X1 U20005 ( .A1(n25663), .A2(n19798), .B1(n25823), .B2(n25655), .ZN(
        n6861) );
  OAI22_X1 U20006 ( .A1(n25663), .A2(n19797), .B1(n25826), .B2(n25655), .ZN(
        n6862) );
  OAI22_X1 U20007 ( .A1(n25663), .A2(n19796), .B1(n25829), .B2(n25655), .ZN(
        n6863) );
  OAI22_X1 U20008 ( .A1(n25663), .A2(n19795), .B1(n25832), .B2(n25655), .ZN(
        n6864) );
  OAI22_X1 U20009 ( .A1(n25663), .A2(n19794), .B1(n25835), .B2(n25655), .ZN(
        n6865) );
  OAI22_X1 U20010 ( .A1(n25663), .A2(n19793), .B1(n25838), .B2(n25655), .ZN(
        n6866) );
  OAI22_X1 U20011 ( .A1(n25663), .A2(n19792), .B1(n25841), .B2(n25655), .ZN(
        n6867) );
  OAI22_X1 U20012 ( .A1(n25663), .A2(n19791), .B1(n25844), .B2(n25655), .ZN(
        n6868) );
  OAI22_X1 U20013 ( .A1(n25663), .A2(n19790), .B1(n25847), .B2(n25655), .ZN(
        n6869) );
  OAI22_X1 U20014 ( .A1(n25663), .A2(n19789), .B1(n25850), .B2(n25655), .ZN(
        n6870) );
  OAI22_X1 U20015 ( .A1(n25663), .A2(n19788), .B1(n25853), .B2(n25656), .ZN(
        n6871) );
  OAI22_X1 U20016 ( .A1(n25664), .A2(n19787), .B1(n25856), .B2(n25656), .ZN(
        n6872) );
  OAI22_X1 U20017 ( .A1(n25664), .A2(n19786), .B1(n25859), .B2(n25656), .ZN(
        n6873) );
  OAI22_X1 U20018 ( .A1(n25664), .A2(n19785), .B1(n25862), .B2(n25656), .ZN(
        n6874) );
  OAI22_X1 U20019 ( .A1(n25664), .A2(n19784), .B1(n25865), .B2(n25656), .ZN(
        n6875) );
  OAI22_X1 U20020 ( .A1(n25664), .A2(n19783), .B1(n25868), .B2(n25656), .ZN(
        n6876) );
  OAI22_X1 U20021 ( .A1(n25664), .A2(n19782), .B1(n25871), .B2(n25656), .ZN(
        n6877) );
  OAI22_X1 U20022 ( .A1(n25664), .A2(n19781), .B1(n25874), .B2(n25656), .ZN(
        n6878) );
  OAI22_X1 U20023 ( .A1(n25664), .A2(n19780), .B1(n25877), .B2(n25656), .ZN(
        n6879) );
  OAI22_X1 U20024 ( .A1(n25664), .A2(n19779), .B1(n25880), .B2(n25656), .ZN(
        n6880) );
  OAI22_X1 U20025 ( .A1(n25664), .A2(n19778), .B1(n25883), .B2(n25656), .ZN(
        n6881) );
  OAI22_X1 U20026 ( .A1(n25664), .A2(n19777), .B1(n25886), .B2(n25656), .ZN(
        n6882) );
  OAI22_X1 U20027 ( .A1(n25664), .A2(n19776), .B1(n25889), .B2(n25657), .ZN(
        n6883) );
  OAI22_X1 U20028 ( .A1(n25664), .A2(n19775), .B1(n25892), .B2(n25657), .ZN(
        n6884) );
  OAI22_X1 U20029 ( .A1(n25665), .A2(n19774), .B1(n25895), .B2(n25657), .ZN(
        n6885) );
  OAI22_X1 U20030 ( .A1(n25665), .A2(n19773), .B1(n25898), .B2(n25657), .ZN(
        n6886) );
  OAI22_X1 U20031 ( .A1(n25665), .A2(n19772), .B1(n25901), .B2(n25657), .ZN(
        n6887) );
  OAI22_X1 U20032 ( .A1(n25665), .A2(n19771), .B1(n25904), .B2(n25657), .ZN(
        n6888) );
  OAI22_X1 U20033 ( .A1(n25665), .A2(n19770), .B1(n25907), .B2(n25657), .ZN(
        n6889) );
  OAI22_X1 U20034 ( .A1(n25665), .A2(n19769), .B1(n25910), .B2(n25657), .ZN(
        n6890) );
  OAI22_X1 U20035 ( .A1(n25665), .A2(n19768), .B1(n25913), .B2(n25657), .ZN(
        n6891) );
  OAI22_X1 U20036 ( .A1(n25665), .A2(n19767), .B1(n25916), .B2(n25657), .ZN(
        n6892) );
  OAI22_X1 U20037 ( .A1(n25665), .A2(n19766), .B1(n25919), .B2(n25657), .ZN(
        n6893) );
  OAI22_X1 U20038 ( .A1(n25665), .A2(n19765), .B1(n25922), .B2(n25657), .ZN(
        n6894) );
  OAI22_X1 U20039 ( .A1(n25665), .A2(n19764), .B1(n25925), .B2(n25658), .ZN(
        n6895) );
  OAI22_X1 U20040 ( .A1(n25665), .A2(n19763), .B1(n25928), .B2(n25658), .ZN(
        n6896) );
  OAI22_X1 U20041 ( .A1(n25665), .A2(n19762), .B1(n25931), .B2(n25658), .ZN(
        n6897) );
  OAI22_X1 U20042 ( .A1(n25666), .A2(n19761), .B1(n25934), .B2(n25658), .ZN(
        n6898) );
  OAI22_X1 U20043 ( .A1(n25666), .A2(n19760), .B1(n25937), .B2(n25658), .ZN(
        n6899) );
  OAI22_X1 U20044 ( .A1(n25666), .A2(n19759), .B1(n25940), .B2(n25658), .ZN(
        n6900) );
  OAI22_X1 U20045 ( .A1(n25666), .A2(n19758), .B1(n25943), .B2(n25658), .ZN(
        n6901) );
  OAI22_X1 U20046 ( .A1(n25666), .A2(n19757), .B1(n25946), .B2(n25658), .ZN(
        n6902) );
  OAI22_X1 U20047 ( .A1(n25666), .A2(n19756), .B1(n25949), .B2(n25658), .ZN(
        n6903) );
  OAI22_X1 U20048 ( .A1(n25666), .A2(n19755), .B1(n25952), .B2(n25658), .ZN(
        n6904) );
  OAI22_X1 U20049 ( .A1(n25666), .A2(n19754), .B1(n25955), .B2(n25658), .ZN(
        n6905) );
  OAI22_X1 U20050 ( .A1(n25666), .A2(n19753), .B1(n25958), .B2(n25658), .ZN(
        n6906) );
  OAI22_X1 U20051 ( .A1(n25713), .A2(n19621), .B1(n25781), .B2(n25705), .ZN(
        n7103) );
  OAI22_X1 U20052 ( .A1(n25713), .A2(n19620), .B1(n25784), .B2(n25705), .ZN(
        n7104) );
  OAI22_X1 U20053 ( .A1(n25713), .A2(n19619), .B1(n25787), .B2(n25705), .ZN(
        n7105) );
  OAI22_X1 U20054 ( .A1(n25713), .A2(n19618), .B1(n25790), .B2(n25705), .ZN(
        n7106) );
  OAI22_X1 U20055 ( .A1(n25713), .A2(n19617), .B1(n25793), .B2(n25705), .ZN(
        n7107) );
  OAI22_X1 U20056 ( .A1(n25713), .A2(n19616), .B1(n25796), .B2(n25705), .ZN(
        n7108) );
  OAI22_X1 U20057 ( .A1(n25713), .A2(n19615), .B1(n25799), .B2(n25705), .ZN(
        n7109) );
  OAI22_X1 U20058 ( .A1(n25713), .A2(n19614), .B1(n25802), .B2(n25705), .ZN(
        n7110) );
  OAI22_X1 U20059 ( .A1(n25713), .A2(n19613), .B1(n25805), .B2(n25705), .ZN(
        n7111) );
  OAI22_X1 U20060 ( .A1(n25713), .A2(n19612), .B1(n25808), .B2(n25705), .ZN(
        n7112) );
  OAI22_X1 U20061 ( .A1(n25713), .A2(n19611), .B1(n25811), .B2(n25705), .ZN(
        n7113) );
  OAI22_X1 U20062 ( .A1(n25713), .A2(n19610), .B1(n25814), .B2(n25705), .ZN(
        n7114) );
  OAI22_X1 U20063 ( .A1(n25714), .A2(n19609), .B1(n25817), .B2(n25706), .ZN(
        n7115) );
  OAI22_X1 U20064 ( .A1(n25714), .A2(n19608), .B1(n25820), .B2(n25706), .ZN(
        n7116) );
  OAI22_X1 U20065 ( .A1(n25714), .A2(n19607), .B1(n25823), .B2(n25706), .ZN(
        n7117) );
  OAI22_X1 U20066 ( .A1(n25714), .A2(n19606), .B1(n25826), .B2(n25706), .ZN(
        n7118) );
  OAI22_X1 U20067 ( .A1(n25714), .A2(n19605), .B1(n25829), .B2(n25706), .ZN(
        n7119) );
  OAI22_X1 U20068 ( .A1(n25714), .A2(n19604), .B1(n25832), .B2(n25706), .ZN(
        n7120) );
  OAI22_X1 U20069 ( .A1(n25714), .A2(n19603), .B1(n25835), .B2(n25706), .ZN(
        n7121) );
  OAI22_X1 U20070 ( .A1(n25714), .A2(n19602), .B1(n25838), .B2(n25706), .ZN(
        n7122) );
  OAI22_X1 U20071 ( .A1(n25714), .A2(n19601), .B1(n25841), .B2(n25706), .ZN(
        n7123) );
  OAI22_X1 U20072 ( .A1(n25714), .A2(n19600), .B1(n25844), .B2(n25706), .ZN(
        n7124) );
  OAI22_X1 U20073 ( .A1(n25714), .A2(n19599), .B1(n25847), .B2(n25706), .ZN(
        n7125) );
  OAI22_X1 U20074 ( .A1(n25714), .A2(n19598), .B1(n25850), .B2(n25706), .ZN(
        n7126) );
  OAI22_X1 U20075 ( .A1(n25714), .A2(n19597), .B1(n25853), .B2(n25707), .ZN(
        n7127) );
  OAI22_X1 U20076 ( .A1(n25715), .A2(n19596), .B1(n25856), .B2(n25707), .ZN(
        n7128) );
  OAI22_X1 U20077 ( .A1(n25715), .A2(n19595), .B1(n25859), .B2(n25707), .ZN(
        n7129) );
  OAI22_X1 U20078 ( .A1(n25715), .A2(n19594), .B1(n25862), .B2(n25707), .ZN(
        n7130) );
  OAI22_X1 U20079 ( .A1(n25715), .A2(n19593), .B1(n25865), .B2(n25707), .ZN(
        n7131) );
  OAI22_X1 U20080 ( .A1(n25715), .A2(n19592), .B1(n25868), .B2(n25707), .ZN(
        n7132) );
  OAI22_X1 U20081 ( .A1(n25715), .A2(n19591), .B1(n25871), .B2(n25707), .ZN(
        n7133) );
  OAI22_X1 U20082 ( .A1(n25715), .A2(n19590), .B1(n25874), .B2(n25707), .ZN(
        n7134) );
  OAI22_X1 U20083 ( .A1(n25715), .A2(n19589), .B1(n25877), .B2(n25707), .ZN(
        n7135) );
  OAI22_X1 U20084 ( .A1(n25715), .A2(n19588), .B1(n25880), .B2(n25707), .ZN(
        n7136) );
  OAI22_X1 U20085 ( .A1(n25715), .A2(n19587), .B1(n25883), .B2(n25707), .ZN(
        n7137) );
  OAI22_X1 U20086 ( .A1(n25715), .A2(n19586), .B1(n25886), .B2(n25707), .ZN(
        n7138) );
  OAI22_X1 U20087 ( .A1(n25715), .A2(n19585), .B1(n25889), .B2(n25708), .ZN(
        n7139) );
  OAI22_X1 U20088 ( .A1(n25715), .A2(n19584), .B1(n25892), .B2(n25708), .ZN(
        n7140) );
  OAI22_X1 U20089 ( .A1(n25716), .A2(n19583), .B1(n25895), .B2(n25708), .ZN(
        n7141) );
  OAI22_X1 U20090 ( .A1(n25716), .A2(n19582), .B1(n25898), .B2(n25708), .ZN(
        n7142) );
  OAI22_X1 U20091 ( .A1(n25716), .A2(n19581), .B1(n25901), .B2(n25708), .ZN(
        n7143) );
  OAI22_X1 U20092 ( .A1(n25716), .A2(n19580), .B1(n25904), .B2(n25708), .ZN(
        n7144) );
  OAI22_X1 U20093 ( .A1(n25716), .A2(n19579), .B1(n25907), .B2(n25708), .ZN(
        n7145) );
  OAI22_X1 U20094 ( .A1(n25716), .A2(n19578), .B1(n25910), .B2(n25708), .ZN(
        n7146) );
  OAI22_X1 U20095 ( .A1(n25716), .A2(n19577), .B1(n25913), .B2(n25708), .ZN(
        n7147) );
  OAI22_X1 U20096 ( .A1(n25716), .A2(n19576), .B1(n25916), .B2(n25708), .ZN(
        n7148) );
  OAI22_X1 U20097 ( .A1(n25716), .A2(n19575), .B1(n25919), .B2(n25708), .ZN(
        n7149) );
  OAI22_X1 U20098 ( .A1(n25716), .A2(n19574), .B1(n25922), .B2(n25708), .ZN(
        n7150) );
  OAI22_X1 U20099 ( .A1(n25716), .A2(n19573), .B1(n25925), .B2(n25709), .ZN(
        n7151) );
  OAI22_X1 U20100 ( .A1(n25716), .A2(n19572), .B1(n25928), .B2(n25709), .ZN(
        n7152) );
  OAI22_X1 U20101 ( .A1(n25716), .A2(n19571), .B1(n25931), .B2(n25709), .ZN(
        n7153) );
  OAI22_X1 U20102 ( .A1(n25717), .A2(n19570), .B1(n25934), .B2(n25709), .ZN(
        n7154) );
  OAI22_X1 U20103 ( .A1(n25717), .A2(n19569), .B1(n25937), .B2(n25709), .ZN(
        n7155) );
  OAI22_X1 U20104 ( .A1(n25717), .A2(n19568), .B1(n25940), .B2(n25709), .ZN(
        n7156) );
  OAI22_X1 U20105 ( .A1(n25717), .A2(n19567), .B1(n25943), .B2(n25709), .ZN(
        n7157) );
  OAI22_X1 U20106 ( .A1(n25717), .A2(n19566), .B1(n25946), .B2(n25709), .ZN(
        n7158) );
  OAI22_X1 U20107 ( .A1(n25717), .A2(n19565), .B1(n25949), .B2(n25709), .ZN(
        n7159) );
  OAI22_X1 U20108 ( .A1(n25717), .A2(n19564), .B1(n25952), .B2(n25709), .ZN(
        n7160) );
  OAI22_X1 U20109 ( .A1(n25717), .A2(n19563), .B1(n25955), .B2(n25709), .ZN(
        n7161) );
  OAI22_X1 U20110 ( .A1(n25717), .A2(n19562), .B1(n25958), .B2(n25709), .ZN(
        n7162) );
  NOR3_X1 U20111 ( .A1(n19492), .A2(n25046), .A3(n19491), .ZN(n23928) );
  NOR3_X1 U20112 ( .A1(n19487), .A2(n25244), .A3(n19486), .ZN(n22731) );
  OAI21_X1 U20113 ( .B1(n21490), .B2(n21512), .A(n25974), .ZN(n21517) );
  OAI21_X1 U20114 ( .B1(n21484), .B2(n21531), .A(n25974), .ZN(n21532) );
  OAI21_X1 U20115 ( .B1(n21490), .B2(n21494), .A(n25973), .ZN(n21499) );
  OAI21_X1 U20116 ( .B1(n21480), .B2(n21487), .A(n25973), .ZN(n21485) );
  BUF_X1 U20117 ( .A(n22788), .Z(n25046) );
  BUF_X1 U20118 ( .A(n21591), .Z(n25244) );
  BUF_X1 U20119 ( .A(n22788), .Z(n25049) );
  BUF_X1 U20120 ( .A(n22788), .Z(n25048) );
  BUF_X1 U20121 ( .A(n22788), .Z(n25047) );
  BUF_X1 U20122 ( .A(n21591), .Z(n25247) );
  BUF_X1 U20123 ( .A(n21591), .Z(n25245) );
  BUF_X1 U20124 ( .A(n21591), .Z(n25246) );
  NOR3_X1 U20125 ( .A1(n19489), .A2(n19493), .A3(n19490), .ZN(n23946) );
  NOR3_X1 U20126 ( .A1(n19484), .A2(n19488), .A3(n19485), .ZN(n22749) );
  NAND2_X1 U20127 ( .A1(n23930), .A2(n23937), .ZN(n22770) );
  NAND2_X1 U20128 ( .A1(n23930), .A2(n23940), .ZN(n22800) );
  NAND2_X1 U20129 ( .A1(n22733), .A2(n22740), .ZN(n21573) );
  NAND2_X1 U20130 ( .A1(n22733), .A2(n22743), .ZN(n21603) );
  NAND2_X1 U20131 ( .A1(n19482), .A2(n19483), .ZN(n21481) );
  BUF_X1 U20132 ( .A(n19478), .Z(n25974) );
  BUF_X1 U20133 ( .A(n19478), .Z(n25973) );
  BUF_X1 U20134 ( .A(n19478), .Z(n25975) );
  NAND2_X1 U20135 ( .A1(n23930), .A2(n23935), .ZN(n22774) );
  NAND2_X1 U20136 ( .A1(n22733), .A2(n22738), .ZN(n21577) );
  BUF_X1 U20137 ( .A(n19478), .Z(n25976) );
  BUF_X1 U20138 ( .A(n19478), .Z(n25977) );
  NAND2_X1 U20139 ( .A1(n23929), .A2(n23930), .ZN(n22760) );
  NAND2_X1 U20140 ( .A1(n23927), .A2(n23930), .ZN(n22765) );
  NAND2_X1 U20141 ( .A1(n23933), .A2(n23930), .ZN(n22795) );
  NAND2_X1 U20142 ( .A1(n22732), .A2(n22733), .ZN(n21563) );
  NAND2_X1 U20143 ( .A1(n22730), .A2(n22733), .ZN(n21568) );
  NAND2_X1 U20144 ( .A1(n22736), .A2(n22733), .ZN(n21598) );
  NAND2_X1 U20145 ( .A1(n23934), .A2(n23939), .ZN(n22784) );
  NAND2_X1 U20146 ( .A1(n23934), .A2(n23940), .ZN(n22799) );
  NAND2_X1 U20147 ( .A1(n22737), .A2(n22742), .ZN(n21587) );
  NAND2_X1 U20148 ( .A1(n22737), .A2(n22743), .ZN(n21602) );
  NAND2_X1 U20149 ( .A1(n23931), .A2(n23940), .ZN(n22794) );
  NAND2_X1 U20150 ( .A1(n22734), .A2(n22743), .ZN(n21597) );
  NAND2_X1 U20151 ( .A1(n23933), .A2(n23934), .ZN(n22790) );
  NAND2_X1 U20152 ( .A1(n23946), .A2(n23934), .ZN(n22785) );
  NAND2_X1 U20153 ( .A1(n22736), .A2(n22737), .ZN(n21593) );
  NAND2_X1 U20154 ( .A1(n22749), .A2(n22737), .ZN(n21588) );
  NAND2_X1 U20155 ( .A1(n23937), .A2(n23931), .ZN(n22775) );
  NAND2_X1 U20156 ( .A1(n22740), .A2(n22734), .ZN(n21578) );
  BUF_X1 U20157 ( .A(n19557), .Z(n25782) );
  BUF_X1 U20158 ( .A(n19556), .Z(n25785) );
  BUF_X1 U20159 ( .A(n19555), .Z(n25788) );
  BUF_X1 U20160 ( .A(n19554), .Z(n25791) );
  BUF_X1 U20161 ( .A(n19553), .Z(n25794) );
  BUF_X1 U20162 ( .A(n19552), .Z(n25797) );
  BUF_X1 U20163 ( .A(n19551), .Z(n25800) );
  BUF_X1 U20164 ( .A(n19550), .Z(n25803) );
  BUF_X1 U20165 ( .A(n19549), .Z(n25806) );
  BUF_X1 U20166 ( .A(n19548), .Z(n25809) );
  BUF_X1 U20167 ( .A(n19547), .Z(n25812) );
  BUF_X1 U20168 ( .A(n19546), .Z(n25815) );
  BUF_X1 U20169 ( .A(n19545), .Z(n25818) );
  BUF_X1 U20170 ( .A(n19544), .Z(n25821) );
  BUF_X1 U20171 ( .A(n19543), .Z(n25824) );
  BUF_X1 U20172 ( .A(n19542), .Z(n25827) );
  BUF_X1 U20173 ( .A(n19541), .Z(n25830) );
  BUF_X1 U20174 ( .A(n19540), .Z(n25833) );
  BUF_X1 U20175 ( .A(n19539), .Z(n25836) );
  BUF_X1 U20176 ( .A(n19538), .Z(n25839) );
  BUF_X1 U20177 ( .A(n19537), .Z(n25842) );
  BUF_X1 U20178 ( .A(n19536), .Z(n25845) );
  BUF_X1 U20179 ( .A(n19535), .Z(n25848) );
  BUF_X1 U20180 ( .A(n19534), .Z(n25851) );
  BUF_X1 U20181 ( .A(n19533), .Z(n25854) );
  BUF_X1 U20182 ( .A(n19532), .Z(n25857) );
  BUF_X1 U20183 ( .A(n19531), .Z(n25860) );
  BUF_X1 U20184 ( .A(n19530), .Z(n25863) );
  BUF_X1 U20185 ( .A(n19529), .Z(n25866) );
  BUF_X1 U20186 ( .A(n19528), .Z(n25869) );
  BUF_X1 U20187 ( .A(n19527), .Z(n25872) );
  BUF_X1 U20188 ( .A(n19526), .Z(n25875) );
  BUF_X1 U20189 ( .A(n19525), .Z(n25878) );
  BUF_X1 U20190 ( .A(n19524), .Z(n25881) );
  BUF_X1 U20191 ( .A(n19523), .Z(n25884) );
  BUF_X1 U20192 ( .A(n19522), .Z(n25887) );
  BUF_X1 U20193 ( .A(n19521), .Z(n25890) );
  BUF_X1 U20194 ( .A(n19520), .Z(n25893) );
  BUF_X1 U20195 ( .A(n19519), .Z(n25896) );
  BUF_X1 U20196 ( .A(n19518), .Z(n25899) );
  BUF_X1 U20197 ( .A(n19517), .Z(n25902) );
  BUF_X1 U20198 ( .A(n19516), .Z(n25905) );
  BUF_X1 U20199 ( .A(n19515), .Z(n25908) );
  BUF_X1 U20200 ( .A(n19514), .Z(n25911) );
  BUF_X1 U20201 ( .A(n19513), .Z(n25914) );
  BUF_X1 U20202 ( .A(n19512), .Z(n25917) );
  BUF_X1 U20203 ( .A(n19511), .Z(n25920) );
  BUF_X1 U20204 ( .A(n19510), .Z(n25923) );
  BUF_X1 U20205 ( .A(n19509), .Z(n25926) );
  BUF_X1 U20206 ( .A(n19508), .Z(n25929) );
  BUF_X1 U20207 ( .A(n19507), .Z(n25932) );
  BUF_X1 U20208 ( .A(n19506), .Z(n25935) );
  BUF_X1 U20209 ( .A(n19505), .Z(n25938) );
  BUF_X1 U20210 ( .A(n19504), .Z(n25941) );
  BUF_X1 U20211 ( .A(n19503), .Z(n25944) );
  BUF_X1 U20212 ( .A(n19502), .Z(n25947) );
  BUF_X1 U20213 ( .A(n19501), .Z(n25950) );
  BUF_X1 U20214 ( .A(n19500), .Z(n25953) );
  BUF_X1 U20215 ( .A(n19499), .Z(n25956) );
  BUF_X1 U20216 ( .A(n19498), .Z(n25959) );
  BUF_X1 U20217 ( .A(n19497), .Z(n25962) );
  BUF_X1 U20218 ( .A(n19496), .Z(n25965) );
  BUF_X1 U20219 ( .A(n19495), .Z(n25968) );
  BUF_X1 U20220 ( .A(n19494), .Z(n25971) );
  BUF_X1 U20221 ( .A(n22788), .Z(n25050) );
  BUF_X1 U20222 ( .A(n21591), .Z(n25248) );
  BUF_X1 U20223 ( .A(n19557), .Z(n25781) );
  BUF_X1 U20224 ( .A(n19556), .Z(n25784) );
  BUF_X1 U20225 ( .A(n19555), .Z(n25787) );
  BUF_X1 U20226 ( .A(n19554), .Z(n25790) );
  BUF_X1 U20227 ( .A(n19553), .Z(n25793) );
  BUF_X1 U20228 ( .A(n19552), .Z(n25796) );
  BUF_X1 U20229 ( .A(n19551), .Z(n25799) );
  BUF_X1 U20230 ( .A(n19550), .Z(n25802) );
  BUF_X1 U20231 ( .A(n19549), .Z(n25805) );
  BUF_X1 U20232 ( .A(n19548), .Z(n25808) );
  BUF_X1 U20233 ( .A(n19547), .Z(n25811) );
  BUF_X1 U20234 ( .A(n19546), .Z(n25814) );
  BUF_X1 U20235 ( .A(n19545), .Z(n25817) );
  BUF_X1 U20236 ( .A(n19544), .Z(n25820) );
  BUF_X1 U20237 ( .A(n19543), .Z(n25823) );
  BUF_X1 U20238 ( .A(n19542), .Z(n25826) );
  BUF_X1 U20239 ( .A(n19541), .Z(n25829) );
  BUF_X1 U20240 ( .A(n19540), .Z(n25832) );
  BUF_X1 U20241 ( .A(n19539), .Z(n25835) );
  BUF_X1 U20242 ( .A(n19538), .Z(n25838) );
  BUF_X1 U20243 ( .A(n19537), .Z(n25841) );
  BUF_X1 U20244 ( .A(n19536), .Z(n25844) );
  BUF_X1 U20245 ( .A(n19535), .Z(n25847) );
  BUF_X1 U20246 ( .A(n19534), .Z(n25850) );
  BUF_X1 U20247 ( .A(n19533), .Z(n25853) );
  BUF_X1 U20248 ( .A(n19532), .Z(n25856) );
  BUF_X1 U20249 ( .A(n19531), .Z(n25859) );
  BUF_X1 U20250 ( .A(n19530), .Z(n25862) );
  BUF_X1 U20251 ( .A(n19529), .Z(n25865) );
  BUF_X1 U20252 ( .A(n19528), .Z(n25868) );
  BUF_X1 U20253 ( .A(n19527), .Z(n25871) );
  BUF_X1 U20254 ( .A(n19526), .Z(n25874) );
  BUF_X1 U20255 ( .A(n19525), .Z(n25877) );
  BUF_X1 U20256 ( .A(n19524), .Z(n25880) );
  BUF_X1 U20257 ( .A(n19523), .Z(n25883) );
  BUF_X1 U20258 ( .A(n19522), .Z(n25886) );
  BUF_X1 U20259 ( .A(n19521), .Z(n25889) );
  BUF_X1 U20260 ( .A(n19520), .Z(n25892) );
  BUF_X1 U20261 ( .A(n19519), .Z(n25895) );
  BUF_X1 U20262 ( .A(n19518), .Z(n25898) );
  BUF_X1 U20263 ( .A(n19517), .Z(n25901) );
  BUF_X1 U20264 ( .A(n19516), .Z(n25904) );
  BUF_X1 U20265 ( .A(n19515), .Z(n25907) );
  BUF_X1 U20266 ( .A(n19514), .Z(n25910) );
  BUF_X1 U20267 ( .A(n19513), .Z(n25913) );
  BUF_X1 U20268 ( .A(n19512), .Z(n25916) );
  BUF_X1 U20269 ( .A(n19511), .Z(n25919) );
  BUF_X1 U20270 ( .A(n19510), .Z(n25922) );
  BUF_X1 U20271 ( .A(n19509), .Z(n25925) );
  BUF_X1 U20272 ( .A(n19508), .Z(n25928) );
  BUF_X1 U20273 ( .A(n19507), .Z(n25931) );
  BUF_X1 U20274 ( .A(n19506), .Z(n25934) );
  BUF_X1 U20275 ( .A(n19505), .Z(n25937) );
  BUF_X1 U20276 ( .A(n19504), .Z(n25940) );
  BUF_X1 U20277 ( .A(n19503), .Z(n25943) );
  BUF_X1 U20278 ( .A(n19502), .Z(n25946) );
  BUF_X1 U20279 ( .A(n19501), .Z(n25949) );
  BUF_X1 U20280 ( .A(n19500), .Z(n25952) );
  BUF_X1 U20281 ( .A(n19499), .Z(n25955) );
  BUF_X1 U20282 ( .A(n19498), .Z(n25958) );
  BUF_X1 U20283 ( .A(n19497), .Z(n25961) );
  BUF_X1 U20284 ( .A(n19496), .Z(n25964) );
  BUF_X1 U20285 ( .A(n19495), .Z(n25967) );
  BUF_X1 U20286 ( .A(n19494), .Z(n25970) );
  NAND2_X1 U20287 ( .A1(n23946), .A2(n23930), .ZN(n22789) );
  NAND2_X1 U20288 ( .A1(n22749), .A2(n22733), .ZN(n21592) );
  NAND2_X1 U20289 ( .A1(n23929), .A2(n23934), .ZN(n22769) );
  NAND2_X1 U20290 ( .A1(n22732), .A2(n22737), .ZN(n21572) );
  NAND2_X1 U20291 ( .A1(n23929), .A2(n23931), .ZN(n22759) );
  NAND2_X1 U20292 ( .A1(n23935), .A2(n23931), .ZN(n22764) );
  NAND2_X1 U20293 ( .A1(n22732), .A2(n22734), .ZN(n21562) );
  NAND2_X1 U20294 ( .A1(n22738), .A2(n22734), .ZN(n21567) );
  OAI21_X1 U20295 ( .B1(n21480), .B2(n21484), .A(n25973), .ZN(n21482) );
  OAI21_X1 U20296 ( .B1(n21480), .B2(n21490), .A(n25973), .ZN(n21488) );
  BUF_X1 U20297 ( .A(n19557), .Z(n25783) );
  BUF_X1 U20298 ( .A(n19556), .Z(n25786) );
  BUF_X1 U20299 ( .A(n19555), .Z(n25789) );
  BUF_X1 U20300 ( .A(n19554), .Z(n25792) );
  BUF_X1 U20301 ( .A(n19553), .Z(n25795) );
  BUF_X1 U20302 ( .A(n19552), .Z(n25798) );
  BUF_X1 U20303 ( .A(n19551), .Z(n25801) );
  BUF_X1 U20304 ( .A(n19550), .Z(n25804) );
  BUF_X1 U20305 ( .A(n19549), .Z(n25807) );
  BUF_X1 U20306 ( .A(n19548), .Z(n25810) );
  BUF_X1 U20307 ( .A(n19547), .Z(n25813) );
  BUF_X1 U20308 ( .A(n19546), .Z(n25816) );
  BUF_X1 U20309 ( .A(n19545), .Z(n25819) );
  BUF_X1 U20310 ( .A(n19544), .Z(n25822) );
  BUF_X1 U20311 ( .A(n19543), .Z(n25825) );
  BUF_X1 U20312 ( .A(n19542), .Z(n25828) );
  BUF_X1 U20313 ( .A(n19541), .Z(n25831) );
  BUF_X1 U20314 ( .A(n19540), .Z(n25834) );
  BUF_X1 U20315 ( .A(n19539), .Z(n25837) );
  BUF_X1 U20316 ( .A(n19538), .Z(n25840) );
  BUF_X1 U20317 ( .A(n19537), .Z(n25843) );
  BUF_X1 U20318 ( .A(n19536), .Z(n25846) );
  BUF_X1 U20319 ( .A(n19535), .Z(n25849) );
  BUF_X1 U20320 ( .A(n19534), .Z(n25852) );
  BUF_X1 U20321 ( .A(n19533), .Z(n25855) );
  BUF_X1 U20322 ( .A(n19532), .Z(n25858) );
  BUF_X1 U20323 ( .A(n19531), .Z(n25861) );
  BUF_X1 U20324 ( .A(n19530), .Z(n25864) );
  BUF_X1 U20325 ( .A(n19529), .Z(n25867) );
  BUF_X1 U20326 ( .A(n19528), .Z(n25870) );
  BUF_X1 U20327 ( .A(n19527), .Z(n25873) );
  BUF_X1 U20328 ( .A(n19526), .Z(n25876) );
  BUF_X1 U20329 ( .A(n19525), .Z(n25879) );
  BUF_X1 U20330 ( .A(n19524), .Z(n25882) );
  BUF_X1 U20331 ( .A(n19523), .Z(n25885) );
  BUF_X1 U20332 ( .A(n19522), .Z(n25888) );
  BUF_X1 U20333 ( .A(n19521), .Z(n25891) );
  BUF_X1 U20334 ( .A(n19520), .Z(n25894) );
  BUF_X1 U20335 ( .A(n19519), .Z(n25897) );
  BUF_X1 U20336 ( .A(n19518), .Z(n25900) );
  BUF_X1 U20337 ( .A(n19517), .Z(n25903) );
  BUF_X1 U20338 ( .A(n19516), .Z(n25906) );
  BUF_X1 U20339 ( .A(n19515), .Z(n25909) );
  BUF_X1 U20340 ( .A(n19514), .Z(n25912) );
  BUF_X1 U20341 ( .A(n19513), .Z(n25915) );
  BUF_X1 U20342 ( .A(n19512), .Z(n25918) );
  BUF_X1 U20343 ( .A(n19511), .Z(n25921) );
  BUF_X1 U20344 ( .A(n19510), .Z(n25924) );
  BUF_X1 U20345 ( .A(n19509), .Z(n25927) );
  BUF_X1 U20346 ( .A(n19508), .Z(n25930) );
  BUF_X1 U20347 ( .A(n19507), .Z(n25933) );
  BUF_X1 U20348 ( .A(n19506), .Z(n25936) );
  BUF_X1 U20349 ( .A(n19505), .Z(n25939) );
  BUF_X1 U20350 ( .A(n19504), .Z(n25942) );
  BUF_X1 U20351 ( .A(n19503), .Z(n25945) );
  BUF_X1 U20352 ( .A(n19502), .Z(n25948) );
  BUF_X1 U20353 ( .A(n19501), .Z(n25951) );
  BUF_X1 U20354 ( .A(n19500), .Z(n25954) );
  BUF_X1 U20355 ( .A(n19499), .Z(n25957) );
  BUF_X1 U20356 ( .A(n19498), .Z(n25960) );
  BUF_X1 U20357 ( .A(n19497), .Z(n25963) );
  BUF_X1 U20358 ( .A(n19496), .Z(n25966) );
  BUF_X1 U20359 ( .A(n19495), .Z(n25969) );
  BUF_X1 U20360 ( .A(n19494), .Z(n25972) );
  OAI21_X1 U20361 ( .B1(n21484), .B2(n21521), .A(n25974), .ZN(n21522) );
  OAI21_X1 U20362 ( .B1(n21490), .B2(n21503), .A(n25973), .ZN(n21508) );
  OAI21_X1 U20363 ( .B1(n21484), .B2(n21549), .A(n25974), .ZN(n21550) );
  OAI21_X1 U20364 ( .B1(n21490), .B2(n21549), .A(n25974), .ZN(n21554) );
  OAI21_X1 U20365 ( .B1(n21490), .B2(n21521), .A(n25974), .ZN(n21526) );
  OAI21_X1 U20366 ( .B1(n21481), .B2(n21494), .A(n25973), .ZN(n21492) );
  OAI21_X1 U20367 ( .B1(n21487), .B2(n21503), .A(n25973), .ZN(n21506) );
  OAI21_X1 U20368 ( .B1(n21487), .B2(n21521), .A(n25974), .ZN(n21524) );
  OAI21_X1 U20369 ( .B1(n21481), .B2(n21549), .A(n25975), .ZN(n21547) );
  OAI21_X1 U20370 ( .B1(n21487), .B2(n21549), .A(n25975), .ZN(n21552) );
  OAI21_X1 U20371 ( .B1(n21487), .B2(n21512), .A(n25974), .ZN(n21515) );
  OAI21_X1 U20372 ( .B1(n21481), .B2(n21503), .A(n25973), .ZN(n21501) );
  OAI21_X1 U20373 ( .B1(n21487), .B2(n21494), .A(n25973), .ZN(n21497) );
  OAI21_X1 U20374 ( .B1(n21484), .B2(n21494), .A(n25973), .ZN(n21495) );
  OAI21_X1 U20375 ( .B1(n21481), .B2(n21540), .A(n25975), .ZN(n21538) );
  OAI21_X1 U20376 ( .B1(n21487), .B2(n21540), .A(n25975), .ZN(n21543) );
  OAI21_X1 U20377 ( .B1(n21490), .B2(n21531), .A(n25975), .ZN(n21536) );
  OAI21_X1 U20378 ( .B1(n21484), .B2(n21540), .A(n25975), .ZN(n21541) );
  OAI21_X1 U20379 ( .B1(n21481), .B2(n21512), .A(n25974), .ZN(n21510) );
  OAI21_X1 U20380 ( .B1(n21481), .B2(n21531), .A(n25974), .ZN(n21529) );
  OAI21_X1 U20381 ( .B1(n21490), .B2(n21540), .A(n25975), .ZN(n21545) );
  OAI21_X1 U20382 ( .B1(n21487), .B2(n21531), .A(n25975), .ZN(n21534) );
  OAI21_X1 U20383 ( .B1(n21484), .B2(n21512), .A(n25974), .ZN(n21513) );
  OAI21_X1 U20384 ( .B1(n21484), .B2(n21503), .A(n25973), .ZN(n21504) );
  AND2_X1 U20385 ( .A1(n23930), .A2(n23939), .ZN(n22787) );
  AND2_X1 U20386 ( .A1(n22733), .A2(n22742), .ZN(n21590) );
  AND2_X1 U20387 ( .A1(n23934), .A2(n23937), .ZN(n22777) );
  AND2_X1 U20388 ( .A1(n22737), .A2(n22740), .ZN(n21580) );
  AND2_X1 U20389 ( .A1(n23935), .A2(n23934), .ZN(n22773) );
  AND2_X1 U20390 ( .A1(n23927), .A2(n23934), .ZN(n22767) );
  AND2_X1 U20391 ( .A1(n22738), .A2(n22737), .ZN(n21576) );
  AND2_X1 U20392 ( .A1(n22730), .A2(n22737), .ZN(n21570) );
  AND2_X1 U20393 ( .A1(n23939), .A2(n23931), .ZN(n22779) );
  AND2_X1 U20394 ( .A1(n23933), .A2(n23931), .ZN(n22768) );
  AND2_X1 U20395 ( .A1(n23946), .A2(n23931), .ZN(n22793) );
  AND2_X1 U20396 ( .A1(n23927), .A2(n23931), .ZN(n22803) );
  AND2_X1 U20397 ( .A1(n22742), .A2(n22734), .ZN(n21582) );
  AND2_X1 U20398 ( .A1(n22736), .A2(n22734), .ZN(n21571) );
  AND2_X1 U20399 ( .A1(n22749), .A2(n22734), .ZN(n21596) );
  AND2_X1 U20400 ( .A1(n22730), .A2(n22734), .ZN(n21606) );
  AND2_X1 U20401 ( .A1(n23928), .A2(n23940), .ZN(n22778) );
  AND2_X1 U20402 ( .A1(n22731), .A2(n22743), .ZN(n21581) );
  AND2_X1 U20403 ( .A1(n23929), .A2(n23928), .ZN(n22762) );
  AND2_X1 U20404 ( .A1(n23927), .A2(n23928), .ZN(n22763) );
  AND2_X1 U20405 ( .A1(n23935), .A2(n23928), .ZN(n22772) );
  AND2_X1 U20406 ( .A1(n23939), .A2(n23928), .ZN(n22792) );
  AND2_X1 U20407 ( .A1(n23933), .A2(n23928), .ZN(n22797) );
  AND2_X1 U20408 ( .A1(n23937), .A2(n23928), .ZN(n22802) );
  AND2_X1 U20409 ( .A1(n22732), .A2(n22731), .ZN(n21565) );
  AND2_X1 U20410 ( .A1(n22730), .A2(n22731), .ZN(n21566) );
  AND2_X1 U20411 ( .A1(n22738), .A2(n22731), .ZN(n21575) );
  AND2_X1 U20412 ( .A1(n22742), .A2(n22731), .ZN(n21595) );
  AND2_X1 U20413 ( .A1(n22736), .A2(n22731), .ZN(n21600) );
  AND2_X1 U20414 ( .A1(n22740), .A2(n22731), .ZN(n21605) );
  OAI221_X1 U20415 ( .B1(n19800), .B2(n25167), .C1(n19864), .C2(n25161), .A(
        n23710), .ZN(n23709) );
  AOI22_X1 U20416 ( .A1(n25155), .A2(n20120), .B1(n25149), .B2(n18220), .ZN(
        n23710) );
  OAI221_X1 U20417 ( .B1(n19799), .B2(n25167), .C1(n19863), .C2(n25161), .A(
        n23692), .ZN(n23691) );
  AOI22_X1 U20418 ( .A1(n25155), .A2(n20119), .B1(n25149), .B2(n18199), .ZN(
        n23692) );
  OAI221_X1 U20419 ( .B1(n19798), .B2(n25167), .C1(n19862), .C2(n25161), .A(
        n23674), .ZN(n23673) );
  AOI22_X1 U20420 ( .A1(n25155), .A2(n20118), .B1(n25149), .B2(n18178), .ZN(
        n23674) );
  OAI221_X1 U20421 ( .B1(n19797), .B2(n25167), .C1(n19861), .C2(n25161), .A(
        n23656), .ZN(n23655) );
  AOI22_X1 U20422 ( .A1(n25155), .A2(n20117), .B1(n25149), .B2(n18157), .ZN(
        n23656) );
  OAI221_X1 U20423 ( .B1(n19796), .B2(n25167), .C1(n19860), .C2(n25161), .A(
        n23638), .ZN(n23637) );
  AOI22_X1 U20424 ( .A1(n25155), .A2(n20116), .B1(n25149), .B2(n18136), .ZN(
        n23638) );
  OAI221_X1 U20425 ( .B1(n19795), .B2(n25167), .C1(n19859), .C2(n25161), .A(
        n23620), .ZN(n23619) );
  AOI22_X1 U20426 ( .A1(n25155), .A2(n20115), .B1(n25149), .B2(n18115), .ZN(
        n23620) );
  OAI221_X1 U20427 ( .B1(n19794), .B2(n25167), .C1(n19858), .C2(n25161), .A(
        n23602), .ZN(n23601) );
  AOI22_X1 U20428 ( .A1(n25155), .A2(n20114), .B1(n25149), .B2(n18094), .ZN(
        n23602) );
  OAI221_X1 U20429 ( .B1(n19793), .B2(n25167), .C1(n19857), .C2(n25161), .A(
        n23584), .ZN(n23583) );
  AOI22_X1 U20430 ( .A1(n25155), .A2(n20113), .B1(n25149), .B2(n18073), .ZN(
        n23584) );
  OAI221_X1 U20431 ( .B1(n19792), .B2(n25167), .C1(n19856), .C2(n25161), .A(
        n23566), .ZN(n23565) );
  AOI22_X1 U20432 ( .A1(n25155), .A2(n20112), .B1(n25149), .B2(n18052), .ZN(
        n23566) );
  OAI221_X1 U20433 ( .B1(n19791), .B2(n25167), .C1(n19855), .C2(n25161), .A(
        n23548), .ZN(n23547) );
  AOI22_X1 U20434 ( .A1(n25155), .A2(n20111), .B1(n25149), .B2(n18031), .ZN(
        n23548) );
  OAI221_X1 U20435 ( .B1(n19790), .B2(n25167), .C1(n19854), .C2(n25161), .A(
        n23530), .ZN(n23529) );
  AOI22_X1 U20436 ( .A1(n25155), .A2(n20110), .B1(n25149), .B2(n18010), .ZN(
        n23530) );
  OAI221_X1 U20437 ( .B1(n19789), .B2(n25167), .C1(n19853), .C2(n25161), .A(
        n23512), .ZN(n23511) );
  AOI22_X1 U20438 ( .A1(n25155), .A2(n20109), .B1(n25149), .B2(n17989), .ZN(
        n23512) );
  OAI221_X1 U20439 ( .B1(n19788), .B2(n25168), .C1(n19852), .C2(n25162), .A(
        n23494), .ZN(n23493) );
  AOI22_X1 U20440 ( .A1(n25156), .A2(n20108), .B1(n25150), .B2(n17968), .ZN(
        n23494) );
  OAI221_X1 U20441 ( .B1(n19787), .B2(n25168), .C1(n19851), .C2(n25162), .A(
        n23476), .ZN(n23475) );
  AOI22_X1 U20442 ( .A1(n25156), .A2(n20107), .B1(n25150), .B2(n17947), .ZN(
        n23476) );
  OAI221_X1 U20443 ( .B1(n19786), .B2(n25168), .C1(n19850), .C2(n25162), .A(
        n23458), .ZN(n23457) );
  AOI22_X1 U20444 ( .A1(n25156), .A2(n20106), .B1(n25150), .B2(n17926), .ZN(
        n23458) );
  OAI221_X1 U20445 ( .B1(n19785), .B2(n25168), .C1(n19849), .C2(n25162), .A(
        n23440), .ZN(n23439) );
  AOI22_X1 U20446 ( .A1(n25156), .A2(n20105), .B1(n25150), .B2(n17905), .ZN(
        n23440) );
  OAI221_X1 U20447 ( .B1(n19784), .B2(n25168), .C1(n19848), .C2(n25162), .A(
        n23422), .ZN(n23421) );
  AOI22_X1 U20448 ( .A1(n25156), .A2(n20104), .B1(n25150), .B2(n17884), .ZN(
        n23422) );
  OAI221_X1 U20449 ( .B1(n19783), .B2(n25168), .C1(n19847), .C2(n25162), .A(
        n23404), .ZN(n23403) );
  AOI22_X1 U20450 ( .A1(n25156), .A2(n20103), .B1(n25150), .B2(n17863), .ZN(
        n23404) );
  OAI221_X1 U20451 ( .B1(n19782), .B2(n25168), .C1(n19846), .C2(n25162), .A(
        n23386), .ZN(n23385) );
  AOI22_X1 U20452 ( .A1(n25156), .A2(n20102), .B1(n25150), .B2(n17842), .ZN(
        n23386) );
  OAI221_X1 U20453 ( .B1(n19781), .B2(n25168), .C1(n19845), .C2(n25162), .A(
        n23368), .ZN(n23367) );
  AOI22_X1 U20454 ( .A1(n25156), .A2(n20101), .B1(n25150), .B2(n17821), .ZN(
        n23368) );
  OAI221_X1 U20455 ( .B1(n19780), .B2(n25168), .C1(n19844), .C2(n25162), .A(
        n23350), .ZN(n23349) );
  AOI22_X1 U20456 ( .A1(n25156), .A2(n20100), .B1(n25150), .B2(n17800), .ZN(
        n23350) );
  OAI221_X1 U20457 ( .B1(n19779), .B2(n25168), .C1(n19843), .C2(n25162), .A(
        n23332), .ZN(n23331) );
  AOI22_X1 U20458 ( .A1(n25156), .A2(n20099), .B1(n25150), .B2(n17779), .ZN(
        n23332) );
  OAI221_X1 U20459 ( .B1(n19778), .B2(n25168), .C1(n19842), .C2(n25162), .A(
        n23314), .ZN(n23313) );
  AOI22_X1 U20460 ( .A1(n25156), .A2(n20098), .B1(n25150), .B2(n17758), .ZN(
        n23314) );
  OAI221_X1 U20461 ( .B1(n19777), .B2(n25168), .C1(n19841), .C2(n25162), .A(
        n23296), .ZN(n23295) );
  AOI22_X1 U20462 ( .A1(n25156), .A2(n20097), .B1(n25150), .B2(n17737), .ZN(
        n23296) );
  OAI221_X1 U20463 ( .B1(n19776), .B2(n25169), .C1(n19840), .C2(n25163), .A(
        n23278), .ZN(n23277) );
  AOI22_X1 U20464 ( .A1(n25157), .A2(n20096), .B1(n25151), .B2(n17716), .ZN(
        n23278) );
  OAI221_X1 U20465 ( .B1(n19775), .B2(n25169), .C1(n19839), .C2(n25163), .A(
        n23260), .ZN(n23259) );
  AOI22_X1 U20466 ( .A1(n25157), .A2(n20095), .B1(n25151), .B2(n17695), .ZN(
        n23260) );
  OAI221_X1 U20467 ( .B1(n19774), .B2(n25169), .C1(n19838), .C2(n25163), .A(
        n23242), .ZN(n23241) );
  AOI22_X1 U20468 ( .A1(n25157), .A2(n20094), .B1(n25151), .B2(n17674), .ZN(
        n23242) );
  OAI221_X1 U20469 ( .B1(n19773), .B2(n25169), .C1(n19837), .C2(n25163), .A(
        n23224), .ZN(n23223) );
  AOI22_X1 U20470 ( .A1(n25157), .A2(n20093), .B1(n25151), .B2(n17653), .ZN(
        n23224) );
  OAI221_X1 U20471 ( .B1(n19772), .B2(n25169), .C1(n19836), .C2(n25163), .A(
        n23206), .ZN(n23205) );
  AOI22_X1 U20472 ( .A1(n25157), .A2(n20092), .B1(n25151), .B2(n17632), .ZN(
        n23206) );
  OAI221_X1 U20473 ( .B1(n19771), .B2(n25169), .C1(n19835), .C2(n25163), .A(
        n23188), .ZN(n23187) );
  AOI22_X1 U20474 ( .A1(n25157), .A2(n20091), .B1(n25151), .B2(n17611), .ZN(
        n23188) );
  OAI221_X1 U20475 ( .B1(n19770), .B2(n25169), .C1(n19834), .C2(n25163), .A(
        n23170), .ZN(n23169) );
  AOI22_X1 U20476 ( .A1(n25157), .A2(n20090), .B1(n25151), .B2(n17590), .ZN(
        n23170) );
  OAI221_X1 U20477 ( .B1(n19769), .B2(n25169), .C1(n19833), .C2(n25163), .A(
        n23152), .ZN(n23151) );
  AOI22_X1 U20478 ( .A1(n25157), .A2(n20089), .B1(n25151), .B2(n17569), .ZN(
        n23152) );
  OAI221_X1 U20479 ( .B1(n19768), .B2(n25169), .C1(n19832), .C2(n25163), .A(
        n23134), .ZN(n23133) );
  AOI22_X1 U20480 ( .A1(n25157), .A2(n20088), .B1(n25151), .B2(n17548), .ZN(
        n23134) );
  OAI221_X1 U20481 ( .B1(n19767), .B2(n25169), .C1(n19831), .C2(n25163), .A(
        n23116), .ZN(n23115) );
  AOI22_X1 U20482 ( .A1(n25157), .A2(n20087), .B1(n25151), .B2(n17527), .ZN(
        n23116) );
  OAI221_X1 U20483 ( .B1(n19766), .B2(n25169), .C1(n19830), .C2(n25163), .A(
        n23098), .ZN(n23097) );
  AOI22_X1 U20484 ( .A1(n25157), .A2(n20086), .B1(n25151), .B2(n17506), .ZN(
        n23098) );
  OAI221_X1 U20485 ( .B1(n19765), .B2(n25169), .C1(n19829), .C2(n25163), .A(
        n23080), .ZN(n23079) );
  AOI22_X1 U20486 ( .A1(n25157), .A2(n20085), .B1(n25151), .B2(n17485), .ZN(
        n23080) );
  OAI221_X1 U20487 ( .B1(n19764), .B2(n25170), .C1(n19828), .C2(n25164), .A(
        n23062), .ZN(n23061) );
  AOI22_X1 U20488 ( .A1(n25158), .A2(n20084), .B1(n25152), .B2(n17464), .ZN(
        n23062) );
  OAI221_X1 U20489 ( .B1(n19763), .B2(n25170), .C1(n19827), .C2(n25164), .A(
        n23044), .ZN(n23043) );
  AOI22_X1 U20490 ( .A1(n25158), .A2(n20083), .B1(n25152), .B2(n17443), .ZN(
        n23044) );
  OAI221_X1 U20491 ( .B1(n19762), .B2(n25170), .C1(n19826), .C2(n25164), .A(
        n23026), .ZN(n23025) );
  AOI22_X1 U20492 ( .A1(n25158), .A2(n20082), .B1(n25152), .B2(n17422), .ZN(
        n23026) );
  OAI221_X1 U20493 ( .B1(n19761), .B2(n25170), .C1(n19825), .C2(n25164), .A(
        n23008), .ZN(n23007) );
  AOI22_X1 U20494 ( .A1(n25158), .A2(n20081), .B1(n25152), .B2(n17401), .ZN(
        n23008) );
  OAI221_X1 U20495 ( .B1(n19760), .B2(n25170), .C1(n19824), .C2(n25164), .A(
        n22990), .ZN(n22989) );
  AOI22_X1 U20496 ( .A1(n25158), .A2(n20080), .B1(n25152), .B2(n17380), .ZN(
        n22990) );
  OAI221_X1 U20497 ( .B1(n19759), .B2(n25170), .C1(n19823), .C2(n25164), .A(
        n22972), .ZN(n22971) );
  AOI22_X1 U20498 ( .A1(n25158), .A2(n20079), .B1(n25152), .B2(n17359), .ZN(
        n22972) );
  OAI221_X1 U20499 ( .B1(n19758), .B2(n25170), .C1(n19822), .C2(n25164), .A(
        n22954), .ZN(n22953) );
  AOI22_X1 U20500 ( .A1(n25158), .A2(n20078), .B1(n25152), .B2(n17338), .ZN(
        n22954) );
  OAI221_X1 U20501 ( .B1(n19757), .B2(n25170), .C1(n19821), .C2(n25164), .A(
        n22936), .ZN(n22935) );
  AOI22_X1 U20502 ( .A1(n25158), .A2(n20077), .B1(n25152), .B2(n17317), .ZN(
        n22936) );
  OAI221_X1 U20503 ( .B1(n19756), .B2(n25170), .C1(n19820), .C2(n25164), .A(
        n22918), .ZN(n22917) );
  AOI22_X1 U20504 ( .A1(n25158), .A2(n20076), .B1(n25152), .B2(n17296), .ZN(
        n22918) );
  OAI221_X1 U20505 ( .B1(n19755), .B2(n25170), .C1(n19819), .C2(n25164), .A(
        n22900), .ZN(n22899) );
  AOI22_X1 U20506 ( .A1(n25158), .A2(n20075), .B1(n25152), .B2(n17275), .ZN(
        n22900) );
  OAI221_X1 U20507 ( .B1(n19754), .B2(n25170), .C1(n19818), .C2(n25164), .A(
        n22882), .ZN(n22881) );
  AOI22_X1 U20508 ( .A1(n25158), .A2(n20074), .B1(n25152), .B2(n17254), .ZN(
        n22882) );
  OAI221_X1 U20509 ( .B1(n19753), .B2(n25170), .C1(n19817), .C2(n25164), .A(
        n22864), .ZN(n22863) );
  AOI22_X1 U20510 ( .A1(n25158), .A2(n20073), .B1(n25152), .B2(n17233), .ZN(
        n22864) );
  OAI221_X1 U20511 ( .B1(n19800), .B2(n25365), .C1(n19864), .C2(n25359), .A(
        n22513), .ZN(n22512) );
  AOI22_X1 U20512 ( .A1(n25353), .A2(n20120), .B1(n25347), .B2(n18220), .ZN(
        n22513) );
  OAI221_X1 U20513 ( .B1(n19799), .B2(n25365), .C1(n19863), .C2(n25359), .A(
        n22495), .ZN(n22494) );
  AOI22_X1 U20514 ( .A1(n25353), .A2(n20119), .B1(n25347), .B2(n18199), .ZN(
        n22495) );
  OAI221_X1 U20515 ( .B1(n19798), .B2(n25365), .C1(n19862), .C2(n25359), .A(
        n22477), .ZN(n22476) );
  AOI22_X1 U20516 ( .A1(n25353), .A2(n20118), .B1(n25347), .B2(n18178), .ZN(
        n22477) );
  OAI221_X1 U20517 ( .B1(n19797), .B2(n25365), .C1(n19861), .C2(n25359), .A(
        n22459), .ZN(n22458) );
  AOI22_X1 U20518 ( .A1(n25353), .A2(n20117), .B1(n25347), .B2(n18157), .ZN(
        n22459) );
  OAI221_X1 U20519 ( .B1(n19796), .B2(n25365), .C1(n19860), .C2(n25359), .A(
        n22441), .ZN(n22440) );
  AOI22_X1 U20520 ( .A1(n25353), .A2(n20116), .B1(n25347), .B2(n18136), .ZN(
        n22441) );
  OAI221_X1 U20521 ( .B1(n19795), .B2(n25365), .C1(n19859), .C2(n25359), .A(
        n22423), .ZN(n22422) );
  AOI22_X1 U20522 ( .A1(n25353), .A2(n20115), .B1(n25347), .B2(n18115), .ZN(
        n22423) );
  OAI221_X1 U20523 ( .B1(n19794), .B2(n25365), .C1(n19858), .C2(n25359), .A(
        n22405), .ZN(n22404) );
  AOI22_X1 U20524 ( .A1(n25353), .A2(n20114), .B1(n25347), .B2(n18094), .ZN(
        n22405) );
  OAI221_X1 U20525 ( .B1(n19793), .B2(n25365), .C1(n19857), .C2(n25359), .A(
        n22387), .ZN(n22386) );
  AOI22_X1 U20526 ( .A1(n25353), .A2(n20113), .B1(n25347), .B2(n18073), .ZN(
        n22387) );
  OAI221_X1 U20527 ( .B1(n19792), .B2(n25365), .C1(n19856), .C2(n25359), .A(
        n22369), .ZN(n22368) );
  AOI22_X1 U20528 ( .A1(n25353), .A2(n20112), .B1(n25347), .B2(n18052), .ZN(
        n22369) );
  OAI221_X1 U20529 ( .B1(n19791), .B2(n25365), .C1(n19855), .C2(n25359), .A(
        n22351), .ZN(n22350) );
  AOI22_X1 U20530 ( .A1(n25353), .A2(n20111), .B1(n25347), .B2(n18031), .ZN(
        n22351) );
  OAI221_X1 U20531 ( .B1(n19790), .B2(n25365), .C1(n19854), .C2(n25359), .A(
        n22333), .ZN(n22332) );
  AOI22_X1 U20532 ( .A1(n25353), .A2(n20110), .B1(n25347), .B2(n18010), .ZN(
        n22333) );
  OAI221_X1 U20533 ( .B1(n19789), .B2(n25365), .C1(n19853), .C2(n25359), .A(
        n22315), .ZN(n22314) );
  AOI22_X1 U20534 ( .A1(n25353), .A2(n20109), .B1(n25347), .B2(n17989), .ZN(
        n22315) );
  OAI221_X1 U20535 ( .B1(n19788), .B2(n25366), .C1(n19852), .C2(n25360), .A(
        n22297), .ZN(n22296) );
  AOI22_X1 U20536 ( .A1(n25354), .A2(n20108), .B1(n25348), .B2(n17968), .ZN(
        n22297) );
  OAI221_X1 U20537 ( .B1(n19787), .B2(n25366), .C1(n19851), .C2(n25360), .A(
        n22279), .ZN(n22278) );
  AOI22_X1 U20538 ( .A1(n25354), .A2(n20107), .B1(n25348), .B2(n17947), .ZN(
        n22279) );
  OAI221_X1 U20539 ( .B1(n19786), .B2(n25366), .C1(n19850), .C2(n25360), .A(
        n22261), .ZN(n22260) );
  AOI22_X1 U20540 ( .A1(n25354), .A2(n20106), .B1(n25348), .B2(n17926), .ZN(
        n22261) );
  OAI221_X1 U20541 ( .B1(n19785), .B2(n25366), .C1(n19849), .C2(n25360), .A(
        n22243), .ZN(n22242) );
  AOI22_X1 U20542 ( .A1(n25354), .A2(n20105), .B1(n25348), .B2(n17905), .ZN(
        n22243) );
  OAI221_X1 U20543 ( .B1(n19784), .B2(n25366), .C1(n19848), .C2(n25360), .A(
        n22225), .ZN(n22224) );
  AOI22_X1 U20544 ( .A1(n25354), .A2(n20104), .B1(n25348), .B2(n17884), .ZN(
        n22225) );
  OAI221_X1 U20545 ( .B1(n19783), .B2(n25366), .C1(n19847), .C2(n25360), .A(
        n22207), .ZN(n22206) );
  AOI22_X1 U20546 ( .A1(n25354), .A2(n20103), .B1(n25348), .B2(n17863), .ZN(
        n22207) );
  OAI221_X1 U20547 ( .B1(n19782), .B2(n25366), .C1(n19846), .C2(n25360), .A(
        n22189), .ZN(n22188) );
  AOI22_X1 U20548 ( .A1(n25354), .A2(n20102), .B1(n25348), .B2(n17842), .ZN(
        n22189) );
  OAI221_X1 U20549 ( .B1(n19781), .B2(n25366), .C1(n19845), .C2(n25360), .A(
        n22171), .ZN(n22170) );
  AOI22_X1 U20550 ( .A1(n25354), .A2(n20101), .B1(n25348), .B2(n17821), .ZN(
        n22171) );
  OAI221_X1 U20551 ( .B1(n19780), .B2(n25366), .C1(n19844), .C2(n25360), .A(
        n22153), .ZN(n22152) );
  AOI22_X1 U20552 ( .A1(n25354), .A2(n20100), .B1(n25348), .B2(n17800), .ZN(
        n22153) );
  OAI221_X1 U20553 ( .B1(n19779), .B2(n25366), .C1(n19843), .C2(n25360), .A(
        n22135), .ZN(n22134) );
  AOI22_X1 U20554 ( .A1(n25354), .A2(n20099), .B1(n25348), .B2(n17779), .ZN(
        n22135) );
  OAI221_X1 U20555 ( .B1(n19778), .B2(n25366), .C1(n19842), .C2(n25360), .A(
        n22117), .ZN(n22116) );
  AOI22_X1 U20556 ( .A1(n25354), .A2(n20098), .B1(n25348), .B2(n17758), .ZN(
        n22117) );
  OAI221_X1 U20557 ( .B1(n19777), .B2(n25366), .C1(n19841), .C2(n25360), .A(
        n22099), .ZN(n22098) );
  AOI22_X1 U20558 ( .A1(n25354), .A2(n20097), .B1(n25348), .B2(n17737), .ZN(
        n22099) );
  OAI221_X1 U20559 ( .B1(n19776), .B2(n25367), .C1(n19840), .C2(n25361), .A(
        n22081), .ZN(n22080) );
  AOI22_X1 U20560 ( .A1(n25355), .A2(n20096), .B1(n25349), .B2(n17716), .ZN(
        n22081) );
  OAI221_X1 U20561 ( .B1(n19775), .B2(n25367), .C1(n19839), .C2(n25361), .A(
        n22063), .ZN(n22062) );
  AOI22_X1 U20562 ( .A1(n25355), .A2(n20095), .B1(n25349), .B2(n17695), .ZN(
        n22063) );
  OAI221_X1 U20563 ( .B1(n19774), .B2(n25367), .C1(n19838), .C2(n25361), .A(
        n22045), .ZN(n22044) );
  AOI22_X1 U20564 ( .A1(n25355), .A2(n20094), .B1(n25349), .B2(n17674), .ZN(
        n22045) );
  OAI221_X1 U20565 ( .B1(n19773), .B2(n25367), .C1(n19837), .C2(n25361), .A(
        n22027), .ZN(n22026) );
  AOI22_X1 U20566 ( .A1(n25355), .A2(n20093), .B1(n25349), .B2(n17653), .ZN(
        n22027) );
  OAI221_X1 U20567 ( .B1(n19772), .B2(n25367), .C1(n19836), .C2(n25361), .A(
        n22009), .ZN(n22008) );
  AOI22_X1 U20568 ( .A1(n25355), .A2(n20092), .B1(n25349), .B2(n17632), .ZN(
        n22009) );
  OAI221_X1 U20569 ( .B1(n19771), .B2(n25367), .C1(n19835), .C2(n25361), .A(
        n21991), .ZN(n21990) );
  AOI22_X1 U20570 ( .A1(n25355), .A2(n20091), .B1(n25349), .B2(n17611), .ZN(
        n21991) );
  OAI221_X1 U20571 ( .B1(n19770), .B2(n25367), .C1(n19834), .C2(n25361), .A(
        n21973), .ZN(n21972) );
  AOI22_X1 U20572 ( .A1(n25355), .A2(n20090), .B1(n25349), .B2(n17590), .ZN(
        n21973) );
  OAI221_X1 U20573 ( .B1(n19769), .B2(n25367), .C1(n19833), .C2(n25361), .A(
        n21955), .ZN(n21954) );
  AOI22_X1 U20574 ( .A1(n25355), .A2(n20089), .B1(n25349), .B2(n17569), .ZN(
        n21955) );
  OAI221_X1 U20575 ( .B1(n19768), .B2(n25367), .C1(n19832), .C2(n25361), .A(
        n21937), .ZN(n21936) );
  AOI22_X1 U20576 ( .A1(n25355), .A2(n20088), .B1(n25349), .B2(n17548), .ZN(
        n21937) );
  OAI221_X1 U20577 ( .B1(n19767), .B2(n25367), .C1(n19831), .C2(n25361), .A(
        n21919), .ZN(n21918) );
  AOI22_X1 U20578 ( .A1(n25355), .A2(n20087), .B1(n25349), .B2(n17527), .ZN(
        n21919) );
  OAI221_X1 U20579 ( .B1(n19766), .B2(n25367), .C1(n19830), .C2(n25361), .A(
        n21901), .ZN(n21900) );
  AOI22_X1 U20580 ( .A1(n25355), .A2(n20086), .B1(n25349), .B2(n17506), .ZN(
        n21901) );
  OAI221_X1 U20581 ( .B1(n19765), .B2(n25367), .C1(n19829), .C2(n25361), .A(
        n21883), .ZN(n21882) );
  AOI22_X1 U20582 ( .A1(n25355), .A2(n20085), .B1(n25349), .B2(n17485), .ZN(
        n21883) );
  OAI221_X1 U20583 ( .B1(n19764), .B2(n25368), .C1(n19828), .C2(n25362), .A(
        n21865), .ZN(n21864) );
  AOI22_X1 U20584 ( .A1(n25356), .A2(n20084), .B1(n25350), .B2(n17464), .ZN(
        n21865) );
  OAI221_X1 U20585 ( .B1(n19763), .B2(n25368), .C1(n19827), .C2(n25362), .A(
        n21847), .ZN(n21846) );
  AOI22_X1 U20586 ( .A1(n25356), .A2(n20083), .B1(n25350), .B2(n17443), .ZN(
        n21847) );
  OAI221_X1 U20587 ( .B1(n19762), .B2(n25368), .C1(n19826), .C2(n25362), .A(
        n21829), .ZN(n21828) );
  AOI22_X1 U20588 ( .A1(n25356), .A2(n20082), .B1(n25350), .B2(n17422), .ZN(
        n21829) );
  OAI221_X1 U20589 ( .B1(n19761), .B2(n25368), .C1(n19825), .C2(n25362), .A(
        n21811), .ZN(n21810) );
  AOI22_X1 U20590 ( .A1(n25356), .A2(n20081), .B1(n25350), .B2(n17401), .ZN(
        n21811) );
  OAI221_X1 U20591 ( .B1(n19760), .B2(n25368), .C1(n19824), .C2(n25362), .A(
        n21793), .ZN(n21792) );
  AOI22_X1 U20592 ( .A1(n25356), .A2(n20080), .B1(n25350), .B2(n17380), .ZN(
        n21793) );
  OAI221_X1 U20593 ( .B1(n19759), .B2(n25368), .C1(n19823), .C2(n25362), .A(
        n21775), .ZN(n21774) );
  AOI22_X1 U20594 ( .A1(n25356), .A2(n20079), .B1(n25350), .B2(n17359), .ZN(
        n21775) );
  OAI221_X1 U20595 ( .B1(n19758), .B2(n25368), .C1(n19822), .C2(n25362), .A(
        n21757), .ZN(n21756) );
  AOI22_X1 U20596 ( .A1(n25356), .A2(n20078), .B1(n25350), .B2(n17338), .ZN(
        n21757) );
  OAI221_X1 U20597 ( .B1(n19757), .B2(n25368), .C1(n19821), .C2(n25362), .A(
        n21739), .ZN(n21738) );
  AOI22_X1 U20598 ( .A1(n25356), .A2(n20077), .B1(n25350), .B2(n17317), .ZN(
        n21739) );
  OAI221_X1 U20599 ( .B1(n19756), .B2(n25368), .C1(n19820), .C2(n25362), .A(
        n21721), .ZN(n21720) );
  AOI22_X1 U20600 ( .A1(n25356), .A2(n20076), .B1(n25350), .B2(n17296), .ZN(
        n21721) );
  OAI221_X1 U20601 ( .B1(n19755), .B2(n25368), .C1(n19819), .C2(n25362), .A(
        n21703), .ZN(n21702) );
  AOI22_X1 U20602 ( .A1(n25356), .A2(n20075), .B1(n25350), .B2(n17275), .ZN(
        n21703) );
  OAI221_X1 U20603 ( .B1(n19754), .B2(n25368), .C1(n19818), .C2(n25362), .A(
        n21685), .ZN(n21684) );
  AOI22_X1 U20604 ( .A1(n25356), .A2(n20074), .B1(n25350), .B2(n17254), .ZN(
        n21685) );
  OAI221_X1 U20605 ( .B1(n19753), .B2(n25368), .C1(n19817), .C2(n25362), .A(
        n21667), .ZN(n21666) );
  AOI22_X1 U20606 ( .A1(n25356), .A2(n20073), .B1(n25350), .B2(n17233), .ZN(
        n21667) );
  OAI221_X1 U20607 ( .B1(n20133), .B2(n25171), .C1(n19813), .C2(n25165), .A(
        n22761), .ZN(n22758) );
  AOI22_X1 U20608 ( .A1(n25159), .A2(n20069), .B1(n25153), .B2(n17149), .ZN(
        n22761) );
  OAI221_X1 U20609 ( .B1(n21098), .B2(n25069), .C1(n20134), .C2(n25063), .A(
        n22786), .ZN(n22783) );
  AOI22_X1 U20610 ( .A1(n25057), .A2(n24085), .B1(n25048), .B2(OUT2[63]), .ZN(
        n22786) );
  OAI221_X1 U20611 ( .B1(n19752), .B2(n25171), .C1(n19816), .C2(n25165), .A(
        n22846), .ZN(n22845) );
  AOI22_X1 U20612 ( .A1(n25159), .A2(n20072), .B1(n25153), .B2(n17212), .ZN(
        n22846) );
  OAI221_X1 U20613 ( .B1(n21101), .B2(n25069), .C1(n20137), .C2(n25063), .A(
        n22854), .ZN(n22853) );
  AOI22_X1 U20614 ( .A1(n25057), .A2(n24079), .B1(n25046), .B2(OUT2[60]), .ZN(
        n22854) );
  OAI221_X1 U20615 ( .B1(n19751), .B2(n25171), .C1(n19815), .C2(n25165), .A(
        n22828), .ZN(n22827) );
  AOI22_X1 U20616 ( .A1(n25159), .A2(n20071), .B1(n25153), .B2(n17191), .ZN(
        n22828) );
  OAI221_X1 U20617 ( .B1(n21100), .B2(n25069), .C1(n20136), .C2(n25063), .A(
        n22836), .ZN(n22835) );
  AOI22_X1 U20618 ( .A1(n25057), .A2(n24081), .B1(n25046), .B2(OUT2[61]), .ZN(
        n22836) );
  OAI221_X1 U20619 ( .B1(n19750), .B2(n25171), .C1(n19814), .C2(n25165), .A(
        n22810), .ZN(n22809) );
  AOI22_X1 U20620 ( .A1(n25159), .A2(n20070), .B1(n25153), .B2(n17170), .ZN(
        n22810) );
  OAI221_X1 U20621 ( .B1(n21099), .B2(n25069), .C1(n20135), .C2(n25063), .A(
        n22818), .ZN(n22817) );
  AOI22_X1 U20622 ( .A1(n25057), .A2(n24083), .B1(n25046), .B2(OUT2[62]), .ZN(
        n22818) );
  OAI221_X1 U20623 ( .B1(n19752), .B2(n25369), .C1(n19816), .C2(n25363), .A(
        n21649), .ZN(n21648) );
  AOI22_X1 U20624 ( .A1(n25357), .A2(n20072), .B1(n25351), .B2(n17212), .ZN(
        n21649) );
  OAI221_X1 U20625 ( .B1(n21101), .B2(n25267), .C1(n20137), .C2(n25261), .A(
        n21657), .ZN(n21656) );
  AOI22_X1 U20626 ( .A1(n25255), .A2(n24079), .B1(n25244), .B2(OUT1[60]), .ZN(
        n21657) );
  OAI221_X1 U20627 ( .B1(n19751), .B2(n25369), .C1(n19815), .C2(n25363), .A(
        n21631), .ZN(n21630) );
  AOI22_X1 U20628 ( .A1(n25357), .A2(n20071), .B1(n25351), .B2(n17191), .ZN(
        n21631) );
  OAI221_X1 U20629 ( .B1(n21100), .B2(n25267), .C1(n20136), .C2(n25261), .A(
        n21639), .ZN(n21638) );
  AOI22_X1 U20630 ( .A1(n25255), .A2(n24081), .B1(n25244), .B2(OUT1[61]), .ZN(
        n21639) );
  OAI221_X1 U20631 ( .B1(n19750), .B2(n25369), .C1(n19814), .C2(n25363), .A(
        n21613), .ZN(n21612) );
  AOI22_X1 U20632 ( .A1(n25357), .A2(n20070), .B1(n25351), .B2(n17170), .ZN(
        n21613) );
  OAI221_X1 U20633 ( .B1(n21099), .B2(n25267), .C1(n20135), .C2(n25261), .A(
        n21621), .ZN(n21620) );
  AOI22_X1 U20634 ( .A1(n25255), .A2(n24083), .B1(n25244), .B2(OUT1[62]), .ZN(
        n21621) );
  OAI221_X1 U20635 ( .B1(n20133), .B2(n25369), .C1(n19813), .C2(n25363), .A(
        n21564), .ZN(n21561) );
  AOI22_X1 U20636 ( .A1(n25357), .A2(n20069), .B1(n25351), .B2(n17149), .ZN(
        n21564) );
  OAI221_X1 U20637 ( .B1(n21098), .B2(n25267), .C1(n20134), .C2(n25261), .A(
        n21589), .ZN(n21586) );
  AOI22_X1 U20638 ( .A1(n25255), .A2(n24085), .B1(n25246), .B2(OUT1[63]), .ZN(
        n21589) );
  OAI221_X1 U20639 ( .B1(n19812), .B2(n25166), .C1(n19876), .C2(n25160), .A(
        n23926), .ZN(n23925) );
  AOI22_X1 U20640 ( .A1(n25154), .A2(n20132), .B1(n25148), .B2(n18472), .ZN(
        n23926) );
  OAI221_X1 U20641 ( .B1(n19811), .B2(n25166), .C1(n19875), .C2(n25160), .A(
        n23908), .ZN(n23907) );
  AOI22_X1 U20642 ( .A1(n25154), .A2(n20131), .B1(n25148), .B2(n18451), .ZN(
        n23908) );
  OAI221_X1 U20643 ( .B1(n19810), .B2(n25166), .C1(n19874), .C2(n25160), .A(
        n23890), .ZN(n23889) );
  AOI22_X1 U20644 ( .A1(n25154), .A2(n20130), .B1(n25148), .B2(n18430), .ZN(
        n23890) );
  OAI221_X1 U20645 ( .B1(n19809), .B2(n25166), .C1(n19873), .C2(n25160), .A(
        n23872), .ZN(n23871) );
  AOI22_X1 U20646 ( .A1(n25154), .A2(n20129), .B1(n25148), .B2(n18409), .ZN(
        n23872) );
  OAI221_X1 U20647 ( .B1(n19808), .B2(n25166), .C1(n19872), .C2(n25160), .A(
        n23854), .ZN(n23853) );
  AOI22_X1 U20648 ( .A1(n25154), .A2(n20128), .B1(n25148), .B2(n18388), .ZN(
        n23854) );
  OAI221_X1 U20649 ( .B1(n19807), .B2(n25166), .C1(n19871), .C2(n25160), .A(
        n23836), .ZN(n23835) );
  AOI22_X1 U20650 ( .A1(n25154), .A2(n20127), .B1(n25148), .B2(n18367), .ZN(
        n23836) );
  OAI221_X1 U20651 ( .B1(n19806), .B2(n25166), .C1(n19870), .C2(n25160), .A(
        n23818), .ZN(n23817) );
  AOI22_X1 U20652 ( .A1(n25154), .A2(n20126), .B1(n25148), .B2(n18346), .ZN(
        n23818) );
  OAI221_X1 U20653 ( .B1(n19805), .B2(n25166), .C1(n19869), .C2(n25160), .A(
        n23800), .ZN(n23799) );
  AOI22_X1 U20654 ( .A1(n25154), .A2(n20125), .B1(n25148), .B2(n18325), .ZN(
        n23800) );
  OAI221_X1 U20655 ( .B1(n19804), .B2(n25166), .C1(n19868), .C2(n25160), .A(
        n23782), .ZN(n23781) );
  AOI22_X1 U20656 ( .A1(n25154), .A2(n20124), .B1(n25148), .B2(n18304), .ZN(
        n23782) );
  OAI221_X1 U20657 ( .B1(n19803), .B2(n25166), .C1(n19867), .C2(n25160), .A(
        n23764), .ZN(n23763) );
  AOI22_X1 U20658 ( .A1(n25154), .A2(n20123), .B1(n25148), .B2(n18283), .ZN(
        n23764) );
  OAI221_X1 U20659 ( .B1(n19802), .B2(n25166), .C1(n19866), .C2(n25160), .A(
        n23746), .ZN(n23745) );
  AOI22_X1 U20660 ( .A1(n25154), .A2(n20122), .B1(n25148), .B2(n18262), .ZN(
        n23746) );
  OAI221_X1 U20661 ( .B1(n19801), .B2(n25166), .C1(n19865), .C2(n25160), .A(
        n23728), .ZN(n23727) );
  AOI22_X1 U20662 ( .A1(n25154), .A2(n20121), .B1(n25148), .B2(n18241), .ZN(
        n23728) );
  OAI221_X1 U20663 ( .B1(n19812), .B2(n25364), .C1(n19876), .C2(n25358), .A(
        n22729), .ZN(n22728) );
  AOI22_X1 U20664 ( .A1(n25352), .A2(n20132), .B1(n25346), .B2(n18472), .ZN(
        n22729) );
  OAI221_X1 U20665 ( .B1(n19811), .B2(n25364), .C1(n19875), .C2(n25358), .A(
        n22711), .ZN(n22710) );
  AOI22_X1 U20666 ( .A1(n25352), .A2(n20131), .B1(n25346), .B2(n18451), .ZN(
        n22711) );
  OAI221_X1 U20667 ( .B1(n19810), .B2(n25364), .C1(n19874), .C2(n25358), .A(
        n22693), .ZN(n22692) );
  AOI22_X1 U20668 ( .A1(n25352), .A2(n20130), .B1(n25346), .B2(n18430), .ZN(
        n22693) );
  OAI221_X1 U20669 ( .B1(n19809), .B2(n25364), .C1(n19873), .C2(n25358), .A(
        n22675), .ZN(n22674) );
  AOI22_X1 U20670 ( .A1(n25352), .A2(n20129), .B1(n25346), .B2(n18409), .ZN(
        n22675) );
  OAI221_X1 U20671 ( .B1(n19808), .B2(n25364), .C1(n19872), .C2(n25358), .A(
        n22657), .ZN(n22656) );
  AOI22_X1 U20672 ( .A1(n25352), .A2(n20128), .B1(n25346), .B2(n18388), .ZN(
        n22657) );
  OAI221_X1 U20673 ( .B1(n19807), .B2(n25364), .C1(n19871), .C2(n25358), .A(
        n22639), .ZN(n22638) );
  AOI22_X1 U20674 ( .A1(n25352), .A2(n20127), .B1(n25346), .B2(n18367), .ZN(
        n22639) );
  OAI221_X1 U20675 ( .B1(n19806), .B2(n25364), .C1(n19870), .C2(n25358), .A(
        n22621), .ZN(n22620) );
  AOI22_X1 U20676 ( .A1(n25352), .A2(n20126), .B1(n25346), .B2(n18346), .ZN(
        n22621) );
  OAI221_X1 U20677 ( .B1(n19805), .B2(n25364), .C1(n19869), .C2(n25358), .A(
        n22603), .ZN(n22602) );
  AOI22_X1 U20678 ( .A1(n25352), .A2(n20125), .B1(n25346), .B2(n18325), .ZN(
        n22603) );
  OAI221_X1 U20679 ( .B1(n19804), .B2(n25364), .C1(n19868), .C2(n25358), .A(
        n22585), .ZN(n22584) );
  AOI22_X1 U20680 ( .A1(n25352), .A2(n20124), .B1(n25346), .B2(n18304), .ZN(
        n22585) );
  OAI221_X1 U20681 ( .B1(n19803), .B2(n25364), .C1(n19867), .C2(n25358), .A(
        n22567), .ZN(n22566) );
  AOI22_X1 U20682 ( .A1(n25352), .A2(n20123), .B1(n25346), .B2(n18283), .ZN(
        n22567) );
  OAI221_X1 U20683 ( .B1(n19802), .B2(n25364), .C1(n19866), .C2(n25358), .A(
        n22549), .ZN(n22548) );
  AOI22_X1 U20684 ( .A1(n25352), .A2(n20122), .B1(n25346), .B2(n18262), .ZN(
        n22549) );
  OAI221_X1 U20685 ( .B1(n19801), .B2(n25364), .C1(n19865), .C2(n25358), .A(
        n22531), .ZN(n22530) );
  AOI22_X1 U20686 ( .A1(n25352), .A2(n20121), .B1(n25346), .B2(n18241), .ZN(
        n22531) );
  OAI221_X1 U20687 ( .B1(n9466), .B2(n25143), .C1(n20449), .C2(n25137), .A(
        n23711), .ZN(n23708) );
  AOI22_X1 U20688 ( .A1(n25131), .A2(n24030), .B1(n25125), .B2(n18219), .ZN(
        n23711) );
  OAI221_X1 U20689 ( .B1(n21149), .B2(n25041), .C1(n20385), .C2(n25035), .A(
        n23719), .ZN(n23716) );
  AOI22_X1 U20690 ( .A1(n25029), .A2(n24339), .B1(n25023), .B2(n18232), .ZN(
        n23719) );
  OAI221_X1 U20691 ( .B1(n9465), .B2(n25143), .C1(n20448), .C2(n25137), .A(
        n23693), .ZN(n23690) );
  AOI22_X1 U20692 ( .A1(n25131), .A2(n24031), .B1(n25125), .B2(n18198), .ZN(
        n23693) );
  OAI221_X1 U20693 ( .B1(n21148), .B2(n25041), .C1(n20384), .C2(n25035), .A(
        n23701), .ZN(n23698) );
  AOI22_X1 U20694 ( .A1(n25029), .A2(n24341), .B1(n25023), .B2(n18211), .ZN(
        n23701) );
  OAI221_X1 U20695 ( .B1(n9464), .B2(n25143), .C1(n20447), .C2(n25137), .A(
        n23675), .ZN(n23672) );
  AOI22_X1 U20696 ( .A1(n25131), .A2(n24032), .B1(n25125), .B2(n18177), .ZN(
        n23675) );
  OAI221_X1 U20697 ( .B1(n21147), .B2(n25041), .C1(n20383), .C2(n25035), .A(
        n23683), .ZN(n23680) );
  AOI22_X1 U20698 ( .A1(n25029), .A2(n24343), .B1(n25023), .B2(n18190), .ZN(
        n23683) );
  OAI221_X1 U20699 ( .B1(n9463), .B2(n25143), .C1(n20446), .C2(n25137), .A(
        n23657), .ZN(n23654) );
  AOI22_X1 U20700 ( .A1(n25131), .A2(n24033), .B1(n25125), .B2(n18156), .ZN(
        n23657) );
  OAI221_X1 U20701 ( .B1(n21146), .B2(n25041), .C1(n20382), .C2(n25035), .A(
        n23665), .ZN(n23662) );
  AOI22_X1 U20702 ( .A1(n25029), .A2(n24345), .B1(n25023), .B2(n18169), .ZN(
        n23665) );
  OAI221_X1 U20703 ( .B1(n9462), .B2(n25143), .C1(n20445), .C2(n25137), .A(
        n23639), .ZN(n23636) );
  AOI22_X1 U20704 ( .A1(n25131), .A2(n24034), .B1(n25125), .B2(n18135), .ZN(
        n23639) );
  OAI221_X1 U20705 ( .B1(n21145), .B2(n25041), .C1(n20381), .C2(n25035), .A(
        n23647), .ZN(n23644) );
  AOI22_X1 U20706 ( .A1(n25029), .A2(n24347), .B1(n25023), .B2(n18148), .ZN(
        n23647) );
  OAI221_X1 U20707 ( .B1(n9461), .B2(n25143), .C1(n20444), .C2(n25137), .A(
        n23621), .ZN(n23618) );
  AOI22_X1 U20708 ( .A1(n25131), .A2(n24035), .B1(n25125), .B2(n18114), .ZN(
        n23621) );
  OAI221_X1 U20709 ( .B1(n21144), .B2(n25041), .C1(n20380), .C2(n25035), .A(
        n23629), .ZN(n23626) );
  AOI22_X1 U20710 ( .A1(n25029), .A2(n24349), .B1(n25023), .B2(n18127), .ZN(
        n23629) );
  OAI221_X1 U20711 ( .B1(n9460), .B2(n25143), .C1(n20443), .C2(n25137), .A(
        n23603), .ZN(n23600) );
  AOI22_X1 U20712 ( .A1(n25131), .A2(n24036), .B1(n25125), .B2(n18093), .ZN(
        n23603) );
  OAI221_X1 U20713 ( .B1(n21143), .B2(n25041), .C1(n20379), .C2(n25035), .A(
        n23611), .ZN(n23608) );
  AOI22_X1 U20714 ( .A1(n25029), .A2(n24351), .B1(n25023), .B2(n18106), .ZN(
        n23611) );
  OAI221_X1 U20715 ( .B1(n9459), .B2(n25143), .C1(n20442), .C2(n25137), .A(
        n23585), .ZN(n23582) );
  AOI22_X1 U20716 ( .A1(n25131), .A2(n24037), .B1(n25125), .B2(n18072), .ZN(
        n23585) );
  OAI221_X1 U20717 ( .B1(n21142), .B2(n25041), .C1(n20378), .C2(n25035), .A(
        n23593), .ZN(n23590) );
  AOI22_X1 U20718 ( .A1(n25029), .A2(n24353), .B1(n25023), .B2(n18085), .ZN(
        n23593) );
  OAI221_X1 U20719 ( .B1(n9458), .B2(n25143), .C1(n20441), .C2(n25137), .A(
        n23567), .ZN(n23564) );
  AOI22_X1 U20720 ( .A1(n25131), .A2(n24038), .B1(n25125), .B2(n18051), .ZN(
        n23567) );
  OAI221_X1 U20721 ( .B1(n21141), .B2(n25041), .C1(n20377), .C2(n25035), .A(
        n23575), .ZN(n23572) );
  AOI22_X1 U20722 ( .A1(n25029), .A2(n24355), .B1(n25023), .B2(n18064), .ZN(
        n23575) );
  OAI221_X1 U20723 ( .B1(n9457), .B2(n25143), .C1(n20440), .C2(n25137), .A(
        n23549), .ZN(n23546) );
  AOI22_X1 U20724 ( .A1(n25131), .A2(n24039), .B1(n25125), .B2(n18030), .ZN(
        n23549) );
  OAI221_X1 U20725 ( .B1(n21140), .B2(n25041), .C1(n20376), .C2(n25035), .A(
        n23557), .ZN(n23554) );
  AOI22_X1 U20726 ( .A1(n25029), .A2(n24357), .B1(n25023), .B2(n18043), .ZN(
        n23557) );
  OAI221_X1 U20727 ( .B1(n9456), .B2(n25143), .C1(n20439), .C2(n25137), .A(
        n23531), .ZN(n23528) );
  AOI22_X1 U20728 ( .A1(n25131), .A2(n24040), .B1(n25125), .B2(n18009), .ZN(
        n23531) );
  OAI221_X1 U20729 ( .B1(n21139), .B2(n25041), .C1(n20375), .C2(n25035), .A(
        n23539), .ZN(n23536) );
  AOI22_X1 U20730 ( .A1(n25029), .A2(n24359), .B1(n25023), .B2(n18022), .ZN(
        n23539) );
  OAI221_X1 U20731 ( .B1(n9455), .B2(n25143), .C1(n20438), .C2(n25137), .A(
        n23513), .ZN(n23510) );
  AOI22_X1 U20732 ( .A1(n25131), .A2(n24041), .B1(n25125), .B2(n17988), .ZN(
        n23513) );
  OAI221_X1 U20733 ( .B1(n21138), .B2(n25041), .C1(n20374), .C2(n25035), .A(
        n23521), .ZN(n23518) );
  AOI22_X1 U20734 ( .A1(n25029), .A2(n24361), .B1(n25023), .B2(n18001), .ZN(
        n23521) );
  OAI221_X1 U20735 ( .B1(n9454), .B2(n25144), .C1(n20437), .C2(n25138), .A(
        n23495), .ZN(n23492) );
  AOI22_X1 U20736 ( .A1(n25132), .A2(n24042), .B1(n25126), .B2(n17967), .ZN(
        n23495) );
  OAI221_X1 U20737 ( .B1(n21137), .B2(n25042), .C1(n20373), .C2(n25036), .A(
        n23503), .ZN(n23500) );
  AOI22_X1 U20738 ( .A1(n25030), .A2(n24363), .B1(n25024), .B2(n17980), .ZN(
        n23503) );
  OAI221_X1 U20739 ( .B1(n9453), .B2(n25144), .C1(n20436), .C2(n25138), .A(
        n23477), .ZN(n23474) );
  AOI22_X1 U20740 ( .A1(n25132), .A2(n24043), .B1(n25126), .B2(n17946), .ZN(
        n23477) );
  OAI221_X1 U20741 ( .B1(n21136), .B2(n25042), .C1(n20372), .C2(n25036), .A(
        n23485), .ZN(n23482) );
  AOI22_X1 U20742 ( .A1(n25030), .A2(n24365), .B1(n25024), .B2(n17959), .ZN(
        n23485) );
  OAI221_X1 U20743 ( .B1(n9452), .B2(n25144), .C1(n20435), .C2(n25138), .A(
        n23459), .ZN(n23456) );
  AOI22_X1 U20744 ( .A1(n25132), .A2(n24044), .B1(n25126), .B2(n17925), .ZN(
        n23459) );
  OAI221_X1 U20745 ( .B1(n21135), .B2(n25042), .C1(n20371), .C2(n25036), .A(
        n23467), .ZN(n23464) );
  AOI22_X1 U20746 ( .A1(n25030), .A2(n24367), .B1(n25024), .B2(n17938), .ZN(
        n23467) );
  OAI221_X1 U20747 ( .B1(n9451), .B2(n25144), .C1(n20434), .C2(n25138), .A(
        n23441), .ZN(n23438) );
  AOI22_X1 U20748 ( .A1(n25132), .A2(n24045), .B1(n25126), .B2(n17904), .ZN(
        n23441) );
  OAI221_X1 U20749 ( .B1(n21134), .B2(n25042), .C1(n20370), .C2(n25036), .A(
        n23449), .ZN(n23446) );
  AOI22_X1 U20750 ( .A1(n25030), .A2(n24369), .B1(n25024), .B2(n17917), .ZN(
        n23449) );
  OAI221_X1 U20751 ( .B1(n9450), .B2(n25144), .C1(n20433), .C2(n25138), .A(
        n23423), .ZN(n23420) );
  AOI22_X1 U20752 ( .A1(n25132), .A2(n24046), .B1(n25126), .B2(n17883), .ZN(
        n23423) );
  OAI221_X1 U20753 ( .B1(n21133), .B2(n25042), .C1(n20369), .C2(n25036), .A(
        n23431), .ZN(n23428) );
  AOI22_X1 U20754 ( .A1(n25030), .A2(n24371), .B1(n25024), .B2(n17896), .ZN(
        n23431) );
  OAI221_X1 U20755 ( .B1(n9449), .B2(n25144), .C1(n20432), .C2(n25138), .A(
        n23405), .ZN(n23402) );
  AOI22_X1 U20756 ( .A1(n25132), .A2(n24047), .B1(n25126), .B2(n17862), .ZN(
        n23405) );
  OAI221_X1 U20757 ( .B1(n21132), .B2(n25042), .C1(n20368), .C2(n25036), .A(
        n23413), .ZN(n23410) );
  AOI22_X1 U20758 ( .A1(n25030), .A2(n24373), .B1(n25024), .B2(n17875), .ZN(
        n23413) );
  OAI221_X1 U20759 ( .B1(n9448), .B2(n25144), .C1(n20431), .C2(n25138), .A(
        n23387), .ZN(n23384) );
  AOI22_X1 U20760 ( .A1(n25132), .A2(n24048), .B1(n25126), .B2(n17841), .ZN(
        n23387) );
  OAI221_X1 U20761 ( .B1(n21131), .B2(n25042), .C1(n20367), .C2(n25036), .A(
        n23395), .ZN(n23392) );
  AOI22_X1 U20762 ( .A1(n25030), .A2(n24375), .B1(n25024), .B2(n17854), .ZN(
        n23395) );
  OAI221_X1 U20763 ( .B1(n9447), .B2(n25144), .C1(n20430), .C2(n25138), .A(
        n23369), .ZN(n23366) );
  AOI22_X1 U20764 ( .A1(n25132), .A2(n24049), .B1(n25126), .B2(n17820), .ZN(
        n23369) );
  OAI221_X1 U20765 ( .B1(n21130), .B2(n25042), .C1(n20366), .C2(n25036), .A(
        n23377), .ZN(n23374) );
  AOI22_X1 U20766 ( .A1(n25030), .A2(n24377), .B1(n25024), .B2(n17833), .ZN(
        n23377) );
  OAI221_X1 U20767 ( .B1(n9446), .B2(n25144), .C1(n20429), .C2(n25138), .A(
        n23351), .ZN(n23348) );
  AOI22_X1 U20768 ( .A1(n25132), .A2(n24050), .B1(n25126), .B2(n17799), .ZN(
        n23351) );
  OAI221_X1 U20769 ( .B1(n21129), .B2(n25042), .C1(n20365), .C2(n25036), .A(
        n23359), .ZN(n23356) );
  AOI22_X1 U20770 ( .A1(n25030), .A2(n24379), .B1(n25024), .B2(n17812), .ZN(
        n23359) );
  OAI221_X1 U20771 ( .B1(n9445), .B2(n25144), .C1(n20428), .C2(n25138), .A(
        n23333), .ZN(n23330) );
  AOI22_X1 U20772 ( .A1(n25132), .A2(n24051), .B1(n25126), .B2(n17778), .ZN(
        n23333) );
  OAI221_X1 U20773 ( .B1(n21128), .B2(n25042), .C1(n20364), .C2(n25036), .A(
        n23341), .ZN(n23338) );
  AOI22_X1 U20774 ( .A1(n25030), .A2(n24381), .B1(n25024), .B2(n17791), .ZN(
        n23341) );
  OAI221_X1 U20775 ( .B1(n9444), .B2(n25144), .C1(n20427), .C2(n25138), .A(
        n23315), .ZN(n23312) );
  AOI22_X1 U20776 ( .A1(n25132), .A2(n24052), .B1(n25126), .B2(n17757), .ZN(
        n23315) );
  OAI221_X1 U20777 ( .B1(n21127), .B2(n25042), .C1(n20363), .C2(n25036), .A(
        n23323), .ZN(n23320) );
  AOI22_X1 U20778 ( .A1(n25030), .A2(n24383), .B1(n25024), .B2(n17770), .ZN(
        n23323) );
  OAI221_X1 U20779 ( .B1(n9443), .B2(n25144), .C1(n20426), .C2(n25138), .A(
        n23297), .ZN(n23294) );
  AOI22_X1 U20780 ( .A1(n25132), .A2(n24053), .B1(n25126), .B2(n17736), .ZN(
        n23297) );
  OAI221_X1 U20781 ( .B1(n21126), .B2(n25042), .C1(n20362), .C2(n25036), .A(
        n23305), .ZN(n23302) );
  AOI22_X1 U20782 ( .A1(n25030), .A2(n24385), .B1(n25024), .B2(n17749), .ZN(
        n23305) );
  OAI221_X1 U20783 ( .B1(n9442), .B2(n25145), .C1(n20425), .C2(n25139), .A(
        n23279), .ZN(n23276) );
  AOI22_X1 U20784 ( .A1(n25133), .A2(n24054), .B1(n25127), .B2(n17715), .ZN(
        n23279) );
  OAI221_X1 U20785 ( .B1(n21125), .B2(n25043), .C1(n20361), .C2(n25037), .A(
        n23287), .ZN(n23284) );
  AOI22_X1 U20786 ( .A1(n25031), .A2(n24387), .B1(n25025), .B2(n17728), .ZN(
        n23287) );
  OAI221_X1 U20787 ( .B1(n9441), .B2(n25145), .C1(n20424), .C2(n25139), .A(
        n23261), .ZN(n23258) );
  AOI22_X1 U20788 ( .A1(n25133), .A2(n24055), .B1(n25127), .B2(n17694), .ZN(
        n23261) );
  OAI221_X1 U20789 ( .B1(n21124), .B2(n25043), .C1(n20360), .C2(n25037), .A(
        n23269), .ZN(n23266) );
  AOI22_X1 U20790 ( .A1(n25031), .A2(n24389), .B1(n25025), .B2(n17707), .ZN(
        n23269) );
  OAI221_X1 U20791 ( .B1(n9440), .B2(n25145), .C1(n20423), .C2(n25139), .A(
        n23243), .ZN(n23240) );
  AOI22_X1 U20792 ( .A1(n25133), .A2(n24056), .B1(n25127), .B2(n17673), .ZN(
        n23243) );
  OAI221_X1 U20793 ( .B1(n21123), .B2(n25043), .C1(n20359), .C2(n25037), .A(
        n23251), .ZN(n23248) );
  AOI22_X1 U20794 ( .A1(n25031), .A2(n24391), .B1(n25025), .B2(n17686), .ZN(
        n23251) );
  OAI221_X1 U20795 ( .B1(n9439), .B2(n25145), .C1(n20422), .C2(n25139), .A(
        n23225), .ZN(n23222) );
  AOI22_X1 U20796 ( .A1(n25133), .A2(n24057), .B1(n25127), .B2(n17652), .ZN(
        n23225) );
  OAI221_X1 U20797 ( .B1(n21122), .B2(n25043), .C1(n20358), .C2(n25037), .A(
        n23233), .ZN(n23230) );
  AOI22_X1 U20798 ( .A1(n25031), .A2(n24393), .B1(n25025), .B2(n17665), .ZN(
        n23233) );
  OAI221_X1 U20799 ( .B1(n9438), .B2(n25145), .C1(n20421), .C2(n25139), .A(
        n23207), .ZN(n23204) );
  AOI22_X1 U20800 ( .A1(n25133), .A2(n24058), .B1(n25127), .B2(n17631), .ZN(
        n23207) );
  OAI221_X1 U20801 ( .B1(n21121), .B2(n25043), .C1(n20357), .C2(n25037), .A(
        n23215), .ZN(n23212) );
  AOI22_X1 U20802 ( .A1(n25031), .A2(n24395), .B1(n25025), .B2(n17644), .ZN(
        n23215) );
  OAI221_X1 U20803 ( .B1(n9437), .B2(n25145), .C1(n20420), .C2(n25139), .A(
        n23189), .ZN(n23186) );
  AOI22_X1 U20804 ( .A1(n25133), .A2(n24059), .B1(n25127), .B2(n17610), .ZN(
        n23189) );
  OAI221_X1 U20805 ( .B1(n21120), .B2(n25043), .C1(n20356), .C2(n25037), .A(
        n23197), .ZN(n23194) );
  AOI22_X1 U20806 ( .A1(n25031), .A2(n24397), .B1(n25025), .B2(n17623), .ZN(
        n23197) );
  OAI221_X1 U20807 ( .B1(n9436), .B2(n25145), .C1(n20419), .C2(n25139), .A(
        n23171), .ZN(n23168) );
  AOI22_X1 U20808 ( .A1(n25133), .A2(n24060), .B1(n25127), .B2(n17589), .ZN(
        n23171) );
  OAI221_X1 U20809 ( .B1(n21119), .B2(n25043), .C1(n20355), .C2(n25037), .A(
        n23179), .ZN(n23176) );
  AOI22_X1 U20810 ( .A1(n25031), .A2(n24399), .B1(n25025), .B2(n17602), .ZN(
        n23179) );
  OAI221_X1 U20811 ( .B1(n9435), .B2(n25145), .C1(n20418), .C2(n25139), .A(
        n23153), .ZN(n23150) );
  AOI22_X1 U20812 ( .A1(n25133), .A2(n24061), .B1(n25127), .B2(n17568), .ZN(
        n23153) );
  OAI221_X1 U20813 ( .B1(n21118), .B2(n25043), .C1(n20354), .C2(n25037), .A(
        n23161), .ZN(n23158) );
  AOI22_X1 U20814 ( .A1(n25031), .A2(n24401), .B1(n25025), .B2(n17581), .ZN(
        n23161) );
  OAI221_X1 U20815 ( .B1(n9434), .B2(n25145), .C1(n20417), .C2(n25139), .A(
        n23135), .ZN(n23132) );
  AOI22_X1 U20816 ( .A1(n25133), .A2(n24062), .B1(n25127), .B2(n17547), .ZN(
        n23135) );
  OAI221_X1 U20817 ( .B1(n21117), .B2(n25043), .C1(n20353), .C2(n25037), .A(
        n23143), .ZN(n23140) );
  AOI22_X1 U20818 ( .A1(n25031), .A2(n24403), .B1(n25025), .B2(n17560), .ZN(
        n23143) );
  OAI221_X1 U20819 ( .B1(n9433), .B2(n25145), .C1(n20416), .C2(n25139), .A(
        n23117), .ZN(n23114) );
  AOI22_X1 U20820 ( .A1(n25133), .A2(n24063), .B1(n25127), .B2(n17526), .ZN(
        n23117) );
  OAI221_X1 U20821 ( .B1(n21116), .B2(n25043), .C1(n20352), .C2(n25037), .A(
        n23125), .ZN(n23122) );
  AOI22_X1 U20822 ( .A1(n25031), .A2(n24405), .B1(n25025), .B2(n17539), .ZN(
        n23125) );
  OAI221_X1 U20823 ( .B1(n9432), .B2(n25145), .C1(n20415), .C2(n25139), .A(
        n23099), .ZN(n23096) );
  AOI22_X1 U20824 ( .A1(n25133), .A2(n24064), .B1(n25127), .B2(n17505), .ZN(
        n23099) );
  OAI221_X1 U20825 ( .B1(n21115), .B2(n25043), .C1(n20351), .C2(n25037), .A(
        n23107), .ZN(n23104) );
  AOI22_X1 U20826 ( .A1(n25031), .A2(n24407), .B1(n25025), .B2(n17518), .ZN(
        n23107) );
  OAI221_X1 U20827 ( .B1(n9431), .B2(n25145), .C1(n20414), .C2(n25139), .A(
        n23081), .ZN(n23078) );
  AOI22_X1 U20828 ( .A1(n25133), .A2(n24065), .B1(n25127), .B2(n17484), .ZN(
        n23081) );
  OAI221_X1 U20829 ( .B1(n21114), .B2(n25043), .C1(n20350), .C2(n25037), .A(
        n23089), .ZN(n23086) );
  AOI22_X1 U20830 ( .A1(n25031), .A2(n24409), .B1(n25025), .B2(n17497), .ZN(
        n23089) );
  OAI221_X1 U20831 ( .B1(n9430), .B2(n25146), .C1(n20413), .C2(n25140), .A(
        n23063), .ZN(n23060) );
  AOI22_X1 U20832 ( .A1(n25134), .A2(n24066), .B1(n25128), .B2(n17463), .ZN(
        n23063) );
  OAI221_X1 U20833 ( .B1(n21113), .B2(n25044), .C1(n20349), .C2(n25038), .A(
        n23071), .ZN(n23068) );
  AOI22_X1 U20834 ( .A1(n25032), .A2(n24411), .B1(n25026), .B2(n17476), .ZN(
        n23071) );
  OAI221_X1 U20835 ( .B1(n9429), .B2(n25146), .C1(n20412), .C2(n25140), .A(
        n23045), .ZN(n23042) );
  AOI22_X1 U20836 ( .A1(n25134), .A2(n24067), .B1(n25128), .B2(n17442), .ZN(
        n23045) );
  OAI221_X1 U20837 ( .B1(n21112), .B2(n25044), .C1(n20348), .C2(n25038), .A(
        n23053), .ZN(n23050) );
  AOI22_X1 U20838 ( .A1(n25032), .A2(n24413), .B1(n25026), .B2(n17455), .ZN(
        n23053) );
  OAI221_X1 U20839 ( .B1(n9428), .B2(n25146), .C1(n20411), .C2(n25140), .A(
        n23027), .ZN(n23024) );
  AOI22_X1 U20840 ( .A1(n25134), .A2(n24068), .B1(n25128), .B2(n17421), .ZN(
        n23027) );
  OAI221_X1 U20841 ( .B1(n21111), .B2(n25044), .C1(n20347), .C2(n25038), .A(
        n23035), .ZN(n23032) );
  AOI22_X1 U20842 ( .A1(n25032), .A2(n24415), .B1(n25026), .B2(n17434), .ZN(
        n23035) );
  OAI221_X1 U20843 ( .B1(n9427), .B2(n25146), .C1(n20410), .C2(n25140), .A(
        n23009), .ZN(n23006) );
  AOI22_X1 U20844 ( .A1(n25134), .A2(n24069), .B1(n25128), .B2(n17400), .ZN(
        n23009) );
  OAI221_X1 U20845 ( .B1(n21110), .B2(n25044), .C1(n20346), .C2(n25038), .A(
        n23017), .ZN(n23014) );
  AOI22_X1 U20846 ( .A1(n25032), .A2(n24417), .B1(n25026), .B2(n17413), .ZN(
        n23017) );
  OAI221_X1 U20847 ( .B1(n9426), .B2(n25146), .C1(n20409), .C2(n25140), .A(
        n22991), .ZN(n22988) );
  AOI22_X1 U20848 ( .A1(n25134), .A2(n24070), .B1(n25128), .B2(n17379), .ZN(
        n22991) );
  OAI221_X1 U20849 ( .B1(n21109), .B2(n25044), .C1(n20345), .C2(n25038), .A(
        n22999), .ZN(n22996) );
  AOI22_X1 U20850 ( .A1(n25032), .A2(n24419), .B1(n25026), .B2(n17392), .ZN(
        n22999) );
  OAI221_X1 U20851 ( .B1(n9425), .B2(n25146), .C1(n20408), .C2(n25140), .A(
        n22973), .ZN(n22970) );
  AOI22_X1 U20852 ( .A1(n25134), .A2(n24071), .B1(n25128), .B2(n17358), .ZN(
        n22973) );
  OAI221_X1 U20853 ( .B1(n21108), .B2(n25044), .C1(n20344), .C2(n25038), .A(
        n22981), .ZN(n22978) );
  AOI22_X1 U20854 ( .A1(n25032), .A2(n24421), .B1(n25026), .B2(n17371), .ZN(
        n22981) );
  OAI221_X1 U20855 ( .B1(n9424), .B2(n25146), .C1(n20407), .C2(n25140), .A(
        n22955), .ZN(n22952) );
  AOI22_X1 U20856 ( .A1(n25134), .A2(n24072), .B1(n25128), .B2(n17337), .ZN(
        n22955) );
  OAI221_X1 U20857 ( .B1(n21107), .B2(n25044), .C1(n20343), .C2(n25038), .A(
        n22963), .ZN(n22960) );
  AOI22_X1 U20858 ( .A1(n25032), .A2(n24423), .B1(n25026), .B2(n17350), .ZN(
        n22963) );
  OAI221_X1 U20859 ( .B1(n9423), .B2(n25146), .C1(n20406), .C2(n25140), .A(
        n22937), .ZN(n22934) );
  AOI22_X1 U20860 ( .A1(n25134), .A2(n24073), .B1(n25128), .B2(n17316), .ZN(
        n22937) );
  OAI221_X1 U20861 ( .B1(n21106), .B2(n25044), .C1(n20342), .C2(n25038), .A(
        n22945), .ZN(n22942) );
  AOI22_X1 U20862 ( .A1(n25032), .A2(n24425), .B1(n25026), .B2(n17329), .ZN(
        n22945) );
  OAI221_X1 U20863 ( .B1(n9422), .B2(n25146), .C1(n20405), .C2(n25140), .A(
        n22919), .ZN(n22916) );
  AOI22_X1 U20864 ( .A1(n25134), .A2(n24074), .B1(n25128), .B2(n17295), .ZN(
        n22919) );
  OAI221_X1 U20865 ( .B1(n21105), .B2(n25044), .C1(n20341), .C2(n25038), .A(
        n22927), .ZN(n22924) );
  AOI22_X1 U20866 ( .A1(n25032), .A2(n24427), .B1(n25026), .B2(n17308), .ZN(
        n22927) );
  OAI221_X1 U20867 ( .B1(n9421), .B2(n25146), .C1(n20404), .C2(n25140), .A(
        n22901), .ZN(n22898) );
  AOI22_X1 U20868 ( .A1(n25134), .A2(n24075), .B1(n25128), .B2(n17274), .ZN(
        n22901) );
  OAI221_X1 U20869 ( .B1(n21104), .B2(n25044), .C1(n20340), .C2(n25038), .A(
        n22909), .ZN(n22906) );
  AOI22_X1 U20870 ( .A1(n25032), .A2(n24429), .B1(n25026), .B2(n17287), .ZN(
        n22909) );
  OAI221_X1 U20871 ( .B1(n9420), .B2(n25146), .C1(n20403), .C2(n25140), .A(
        n22883), .ZN(n22880) );
  AOI22_X1 U20872 ( .A1(n25134), .A2(n24076), .B1(n25128), .B2(n17253), .ZN(
        n22883) );
  OAI221_X1 U20873 ( .B1(n21103), .B2(n25044), .C1(n20339), .C2(n25038), .A(
        n22891), .ZN(n22888) );
  AOI22_X1 U20874 ( .A1(n25032), .A2(n24431), .B1(n25026), .B2(n17266), .ZN(
        n22891) );
  OAI221_X1 U20875 ( .B1(n9419), .B2(n25146), .C1(n20402), .C2(n25140), .A(
        n22865), .ZN(n22862) );
  AOI22_X1 U20876 ( .A1(n25134), .A2(n24077), .B1(n25128), .B2(n17232), .ZN(
        n22865) );
  OAI221_X1 U20877 ( .B1(n21102), .B2(n25044), .C1(n20338), .C2(n25038), .A(
        n22873), .ZN(n22870) );
  AOI22_X1 U20878 ( .A1(n25032), .A2(n24433), .B1(n25026), .B2(n17245), .ZN(
        n22873) );
  OAI221_X1 U20879 ( .B1(n9466), .B2(n25341), .C1(n20449), .C2(n25335), .A(
        n22514), .ZN(n22511) );
  AOI22_X1 U20880 ( .A1(n25329), .A2(n24030), .B1(n25323), .B2(n18219), .ZN(
        n22514) );
  OAI221_X1 U20881 ( .B1(n21149), .B2(n25239), .C1(n20385), .C2(n25233), .A(
        n22522), .ZN(n22519) );
  AOI22_X1 U20882 ( .A1(n25227), .A2(n24339), .B1(n25221), .B2(n18232), .ZN(
        n22522) );
  OAI221_X1 U20883 ( .B1(n9465), .B2(n25341), .C1(n20448), .C2(n25335), .A(
        n22496), .ZN(n22493) );
  AOI22_X1 U20884 ( .A1(n25329), .A2(n24031), .B1(n25323), .B2(n18198), .ZN(
        n22496) );
  OAI221_X1 U20885 ( .B1(n21148), .B2(n25239), .C1(n20384), .C2(n25233), .A(
        n22504), .ZN(n22501) );
  AOI22_X1 U20886 ( .A1(n25227), .A2(n24341), .B1(n25221), .B2(n18211), .ZN(
        n22504) );
  OAI221_X1 U20887 ( .B1(n9464), .B2(n25341), .C1(n20447), .C2(n25335), .A(
        n22478), .ZN(n22475) );
  AOI22_X1 U20888 ( .A1(n25329), .A2(n24032), .B1(n25323), .B2(n18177), .ZN(
        n22478) );
  OAI221_X1 U20889 ( .B1(n21147), .B2(n25239), .C1(n20383), .C2(n25233), .A(
        n22486), .ZN(n22483) );
  AOI22_X1 U20890 ( .A1(n25227), .A2(n24343), .B1(n25221), .B2(n18190), .ZN(
        n22486) );
  OAI221_X1 U20891 ( .B1(n9463), .B2(n25341), .C1(n20446), .C2(n25335), .A(
        n22460), .ZN(n22457) );
  AOI22_X1 U20892 ( .A1(n25329), .A2(n24033), .B1(n25323), .B2(n18156), .ZN(
        n22460) );
  OAI221_X1 U20893 ( .B1(n21146), .B2(n25239), .C1(n20382), .C2(n25233), .A(
        n22468), .ZN(n22465) );
  AOI22_X1 U20894 ( .A1(n25227), .A2(n24345), .B1(n25221), .B2(n18169), .ZN(
        n22468) );
  OAI221_X1 U20895 ( .B1(n9462), .B2(n25341), .C1(n20445), .C2(n25335), .A(
        n22442), .ZN(n22439) );
  AOI22_X1 U20896 ( .A1(n25329), .A2(n24034), .B1(n25323), .B2(n18135), .ZN(
        n22442) );
  OAI221_X1 U20897 ( .B1(n21145), .B2(n25239), .C1(n20381), .C2(n25233), .A(
        n22450), .ZN(n22447) );
  AOI22_X1 U20898 ( .A1(n25227), .A2(n24347), .B1(n25221), .B2(n18148), .ZN(
        n22450) );
  OAI221_X1 U20899 ( .B1(n9461), .B2(n25341), .C1(n20444), .C2(n25335), .A(
        n22424), .ZN(n22421) );
  AOI22_X1 U20900 ( .A1(n25329), .A2(n24035), .B1(n25323), .B2(n18114), .ZN(
        n22424) );
  OAI221_X1 U20901 ( .B1(n21144), .B2(n25239), .C1(n20380), .C2(n25233), .A(
        n22432), .ZN(n22429) );
  AOI22_X1 U20902 ( .A1(n25227), .A2(n24349), .B1(n25221), .B2(n18127), .ZN(
        n22432) );
  OAI221_X1 U20903 ( .B1(n9460), .B2(n25341), .C1(n20443), .C2(n25335), .A(
        n22406), .ZN(n22403) );
  AOI22_X1 U20904 ( .A1(n25329), .A2(n24036), .B1(n25323), .B2(n18093), .ZN(
        n22406) );
  OAI221_X1 U20905 ( .B1(n21143), .B2(n25239), .C1(n20379), .C2(n25233), .A(
        n22414), .ZN(n22411) );
  AOI22_X1 U20906 ( .A1(n25227), .A2(n24351), .B1(n25221), .B2(n18106), .ZN(
        n22414) );
  OAI221_X1 U20907 ( .B1(n9459), .B2(n25341), .C1(n20442), .C2(n25335), .A(
        n22388), .ZN(n22385) );
  AOI22_X1 U20908 ( .A1(n25329), .A2(n24037), .B1(n25323), .B2(n18072), .ZN(
        n22388) );
  OAI221_X1 U20909 ( .B1(n21142), .B2(n25239), .C1(n20378), .C2(n25233), .A(
        n22396), .ZN(n22393) );
  AOI22_X1 U20910 ( .A1(n25227), .A2(n24353), .B1(n25221), .B2(n18085), .ZN(
        n22396) );
  OAI221_X1 U20911 ( .B1(n9458), .B2(n25341), .C1(n20441), .C2(n25335), .A(
        n22370), .ZN(n22367) );
  AOI22_X1 U20912 ( .A1(n25329), .A2(n24038), .B1(n25323), .B2(n18051), .ZN(
        n22370) );
  OAI221_X1 U20913 ( .B1(n21141), .B2(n25239), .C1(n20377), .C2(n25233), .A(
        n22378), .ZN(n22375) );
  AOI22_X1 U20914 ( .A1(n25227), .A2(n24355), .B1(n25221), .B2(n18064), .ZN(
        n22378) );
  OAI221_X1 U20915 ( .B1(n9457), .B2(n25341), .C1(n20440), .C2(n25335), .A(
        n22352), .ZN(n22349) );
  AOI22_X1 U20916 ( .A1(n25329), .A2(n24039), .B1(n25323), .B2(n18030), .ZN(
        n22352) );
  OAI221_X1 U20917 ( .B1(n21140), .B2(n25239), .C1(n20376), .C2(n25233), .A(
        n22360), .ZN(n22357) );
  AOI22_X1 U20918 ( .A1(n25227), .A2(n24357), .B1(n25221), .B2(n18043), .ZN(
        n22360) );
  OAI221_X1 U20919 ( .B1(n9456), .B2(n25341), .C1(n20439), .C2(n25335), .A(
        n22334), .ZN(n22331) );
  AOI22_X1 U20920 ( .A1(n25329), .A2(n24040), .B1(n25323), .B2(n18009), .ZN(
        n22334) );
  OAI221_X1 U20921 ( .B1(n21139), .B2(n25239), .C1(n20375), .C2(n25233), .A(
        n22342), .ZN(n22339) );
  AOI22_X1 U20922 ( .A1(n25227), .A2(n24359), .B1(n25221), .B2(n18022), .ZN(
        n22342) );
  OAI221_X1 U20923 ( .B1(n9455), .B2(n25341), .C1(n20438), .C2(n25335), .A(
        n22316), .ZN(n22313) );
  AOI22_X1 U20924 ( .A1(n25329), .A2(n24041), .B1(n25323), .B2(n17988), .ZN(
        n22316) );
  OAI221_X1 U20925 ( .B1(n21138), .B2(n25239), .C1(n20374), .C2(n25233), .A(
        n22324), .ZN(n22321) );
  AOI22_X1 U20926 ( .A1(n25227), .A2(n24361), .B1(n25221), .B2(n18001), .ZN(
        n22324) );
  OAI221_X1 U20927 ( .B1(n9454), .B2(n25342), .C1(n20437), .C2(n25336), .A(
        n22298), .ZN(n22295) );
  AOI22_X1 U20928 ( .A1(n25330), .A2(n24042), .B1(n25324), .B2(n17967), .ZN(
        n22298) );
  OAI221_X1 U20929 ( .B1(n21137), .B2(n25240), .C1(n20373), .C2(n25234), .A(
        n22306), .ZN(n22303) );
  AOI22_X1 U20930 ( .A1(n25228), .A2(n24363), .B1(n25222), .B2(n17980), .ZN(
        n22306) );
  OAI221_X1 U20931 ( .B1(n9453), .B2(n25342), .C1(n20436), .C2(n25336), .A(
        n22280), .ZN(n22277) );
  AOI22_X1 U20932 ( .A1(n25330), .A2(n24043), .B1(n25324), .B2(n17946), .ZN(
        n22280) );
  OAI221_X1 U20933 ( .B1(n21136), .B2(n25240), .C1(n20372), .C2(n25234), .A(
        n22288), .ZN(n22285) );
  AOI22_X1 U20934 ( .A1(n25228), .A2(n24365), .B1(n25222), .B2(n17959), .ZN(
        n22288) );
  OAI221_X1 U20935 ( .B1(n9452), .B2(n25342), .C1(n20435), .C2(n25336), .A(
        n22262), .ZN(n22259) );
  AOI22_X1 U20936 ( .A1(n25330), .A2(n24044), .B1(n25324), .B2(n17925), .ZN(
        n22262) );
  OAI221_X1 U20937 ( .B1(n21135), .B2(n25240), .C1(n20371), .C2(n25234), .A(
        n22270), .ZN(n22267) );
  AOI22_X1 U20938 ( .A1(n25228), .A2(n24367), .B1(n25222), .B2(n17938), .ZN(
        n22270) );
  OAI221_X1 U20939 ( .B1(n9451), .B2(n25342), .C1(n20434), .C2(n25336), .A(
        n22244), .ZN(n22241) );
  AOI22_X1 U20940 ( .A1(n25330), .A2(n24045), .B1(n25324), .B2(n17904), .ZN(
        n22244) );
  OAI221_X1 U20941 ( .B1(n21134), .B2(n25240), .C1(n20370), .C2(n25234), .A(
        n22252), .ZN(n22249) );
  AOI22_X1 U20942 ( .A1(n25228), .A2(n24369), .B1(n25222), .B2(n17917), .ZN(
        n22252) );
  OAI221_X1 U20943 ( .B1(n9450), .B2(n25342), .C1(n20433), .C2(n25336), .A(
        n22226), .ZN(n22223) );
  AOI22_X1 U20944 ( .A1(n25330), .A2(n24046), .B1(n25324), .B2(n17883), .ZN(
        n22226) );
  OAI221_X1 U20945 ( .B1(n21133), .B2(n25240), .C1(n20369), .C2(n25234), .A(
        n22234), .ZN(n22231) );
  AOI22_X1 U20946 ( .A1(n25228), .A2(n24371), .B1(n25222), .B2(n17896), .ZN(
        n22234) );
  OAI221_X1 U20947 ( .B1(n9449), .B2(n25342), .C1(n20432), .C2(n25336), .A(
        n22208), .ZN(n22205) );
  AOI22_X1 U20948 ( .A1(n25330), .A2(n24047), .B1(n25324), .B2(n17862), .ZN(
        n22208) );
  OAI221_X1 U20949 ( .B1(n21132), .B2(n25240), .C1(n20368), .C2(n25234), .A(
        n22216), .ZN(n22213) );
  AOI22_X1 U20950 ( .A1(n25228), .A2(n24373), .B1(n25222), .B2(n17875), .ZN(
        n22216) );
  OAI221_X1 U20951 ( .B1(n9448), .B2(n25342), .C1(n20431), .C2(n25336), .A(
        n22190), .ZN(n22187) );
  AOI22_X1 U20952 ( .A1(n25330), .A2(n24048), .B1(n25324), .B2(n17841), .ZN(
        n22190) );
  OAI221_X1 U20953 ( .B1(n21131), .B2(n25240), .C1(n20367), .C2(n25234), .A(
        n22198), .ZN(n22195) );
  AOI22_X1 U20954 ( .A1(n25228), .A2(n24375), .B1(n25222), .B2(n17854), .ZN(
        n22198) );
  OAI221_X1 U20955 ( .B1(n9447), .B2(n25342), .C1(n20430), .C2(n25336), .A(
        n22172), .ZN(n22169) );
  AOI22_X1 U20956 ( .A1(n25330), .A2(n24049), .B1(n25324), .B2(n17820), .ZN(
        n22172) );
  OAI221_X1 U20957 ( .B1(n21130), .B2(n25240), .C1(n20366), .C2(n25234), .A(
        n22180), .ZN(n22177) );
  AOI22_X1 U20958 ( .A1(n25228), .A2(n24377), .B1(n25222), .B2(n17833), .ZN(
        n22180) );
  OAI221_X1 U20959 ( .B1(n9446), .B2(n25342), .C1(n20429), .C2(n25336), .A(
        n22154), .ZN(n22151) );
  AOI22_X1 U20960 ( .A1(n25330), .A2(n24050), .B1(n25324), .B2(n17799), .ZN(
        n22154) );
  OAI221_X1 U20961 ( .B1(n21129), .B2(n25240), .C1(n20365), .C2(n25234), .A(
        n22162), .ZN(n22159) );
  AOI22_X1 U20962 ( .A1(n25228), .A2(n24379), .B1(n25222), .B2(n17812), .ZN(
        n22162) );
  OAI221_X1 U20963 ( .B1(n9445), .B2(n25342), .C1(n20428), .C2(n25336), .A(
        n22136), .ZN(n22133) );
  AOI22_X1 U20964 ( .A1(n25330), .A2(n24051), .B1(n25324), .B2(n17778), .ZN(
        n22136) );
  OAI221_X1 U20965 ( .B1(n21128), .B2(n25240), .C1(n20364), .C2(n25234), .A(
        n22144), .ZN(n22141) );
  AOI22_X1 U20966 ( .A1(n25228), .A2(n24381), .B1(n25222), .B2(n17791), .ZN(
        n22144) );
  OAI221_X1 U20967 ( .B1(n9444), .B2(n25342), .C1(n20427), .C2(n25336), .A(
        n22118), .ZN(n22115) );
  AOI22_X1 U20968 ( .A1(n25330), .A2(n24052), .B1(n25324), .B2(n17757), .ZN(
        n22118) );
  OAI221_X1 U20969 ( .B1(n21127), .B2(n25240), .C1(n20363), .C2(n25234), .A(
        n22126), .ZN(n22123) );
  AOI22_X1 U20970 ( .A1(n25228), .A2(n24383), .B1(n25222), .B2(n17770), .ZN(
        n22126) );
  OAI221_X1 U20971 ( .B1(n9443), .B2(n25342), .C1(n20426), .C2(n25336), .A(
        n22100), .ZN(n22097) );
  AOI22_X1 U20972 ( .A1(n25330), .A2(n24053), .B1(n25324), .B2(n17736), .ZN(
        n22100) );
  OAI221_X1 U20973 ( .B1(n21126), .B2(n25240), .C1(n20362), .C2(n25234), .A(
        n22108), .ZN(n22105) );
  AOI22_X1 U20974 ( .A1(n25228), .A2(n24385), .B1(n25222), .B2(n17749), .ZN(
        n22108) );
  OAI221_X1 U20975 ( .B1(n9442), .B2(n25343), .C1(n20425), .C2(n25337), .A(
        n22082), .ZN(n22079) );
  AOI22_X1 U20976 ( .A1(n25331), .A2(n24054), .B1(n25325), .B2(n17715), .ZN(
        n22082) );
  OAI221_X1 U20977 ( .B1(n21125), .B2(n25241), .C1(n20361), .C2(n25235), .A(
        n22090), .ZN(n22087) );
  AOI22_X1 U20978 ( .A1(n25229), .A2(n24387), .B1(n25223), .B2(n17728), .ZN(
        n22090) );
  OAI221_X1 U20979 ( .B1(n9441), .B2(n25343), .C1(n20424), .C2(n25337), .A(
        n22064), .ZN(n22061) );
  AOI22_X1 U20980 ( .A1(n25331), .A2(n24055), .B1(n25325), .B2(n17694), .ZN(
        n22064) );
  OAI221_X1 U20981 ( .B1(n21124), .B2(n25241), .C1(n20360), .C2(n25235), .A(
        n22072), .ZN(n22069) );
  AOI22_X1 U20982 ( .A1(n25229), .A2(n24389), .B1(n25223), .B2(n17707), .ZN(
        n22072) );
  OAI221_X1 U20983 ( .B1(n9440), .B2(n25343), .C1(n20423), .C2(n25337), .A(
        n22046), .ZN(n22043) );
  AOI22_X1 U20984 ( .A1(n25331), .A2(n24056), .B1(n25325), .B2(n17673), .ZN(
        n22046) );
  OAI221_X1 U20985 ( .B1(n21123), .B2(n25241), .C1(n20359), .C2(n25235), .A(
        n22054), .ZN(n22051) );
  AOI22_X1 U20986 ( .A1(n25229), .A2(n24391), .B1(n25223), .B2(n17686), .ZN(
        n22054) );
  OAI221_X1 U20987 ( .B1(n9439), .B2(n25343), .C1(n20422), .C2(n25337), .A(
        n22028), .ZN(n22025) );
  AOI22_X1 U20988 ( .A1(n25331), .A2(n24057), .B1(n25325), .B2(n17652), .ZN(
        n22028) );
  OAI221_X1 U20989 ( .B1(n21122), .B2(n25241), .C1(n20358), .C2(n25235), .A(
        n22036), .ZN(n22033) );
  AOI22_X1 U20990 ( .A1(n25229), .A2(n24393), .B1(n25223), .B2(n17665), .ZN(
        n22036) );
  OAI221_X1 U20991 ( .B1(n9438), .B2(n25343), .C1(n20421), .C2(n25337), .A(
        n22010), .ZN(n22007) );
  AOI22_X1 U20992 ( .A1(n25331), .A2(n24058), .B1(n25325), .B2(n17631), .ZN(
        n22010) );
  OAI221_X1 U20993 ( .B1(n21121), .B2(n25241), .C1(n20357), .C2(n25235), .A(
        n22018), .ZN(n22015) );
  AOI22_X1 U20994 ( .A1(n25229), .A2(n24395), .B1(n25223), .B2(n17644), .ZN(
        n22018) );
  OAI221_X1 U20995 ( .B1(n9437), .B2(n25343), .C1(n20420), .C2(n25337), .A(
        n21992), .ZN(n21989) );
  AOI22_X1 U20996 ( .A1(n25331), .A2(n24059), .B1(n25325), .B2(n17610), .ZN(
        n21992) );
  OAI221_X1 U20997 ( .B1(n21120), .B2(n25241), .C1(n20356), .C2(n25235), .A(
        n22000), .ZN(n21997) );
  AOI22_X1 U20998 ( .A1(n25229), .A2(n24397), .B1(n25223), .B2(n17623), .ZN(
        n22000) );
  OAI221_X1 U20999 ( .B1(n9436), .B2(n25343), .C1(n20419), .C2(n25337), .A(
        n21974), .ZN(n21971) );
  AOI22_X1 U21000 ( .A1(n25331), .A2(n24060), .B1(n25325), .B2(n17589), .ZN(
        n21974) );
  OAI221_X1 U21001 ( .B1(n21119), .B2(n25241), .C1(n20355), .C2(n25235), .A(
        n21982), .ZN(n21979) );
  AOI22_X1 U21002 ( .A1(n25229), .A2(n24399), .B1(n25223), .B2(n17602), .ZN(
        n21982) );
  OAI221_X1 U21003 ( .B1(n9435), .B2(n25343), .C1(n20418), .C2(n25337), .A(
        n21956), .ZN(n21953) );
  AOI22_X1 U21004 ( .A1(n25331), .A2(n24061), .B1(n25325), .B2(n17568), .ZN(
        n21956) );
  OAI221_X1 U21005 ( .B1(n21118), .B2(n25241), .C1(n20354), .C2(n25235), .A(
        n21964), .ZN(n21961) );
  AOI22_X1 U21006 ( .A1(n25229), .A2(n24401), .B1(n25223), .B2(n17581), .ZN(
        n21964) );
  OAI221_X1 U21007 ( .B1(n9434), .B2(n25343), .C1(n20417), .C2(n25337), .A(
        n21938), .ZN(n21935) );
  AOI22_X1 U21008 ( .A1(n25331), .A2(n24062), .B1(n25325), .B2(n17547), .ZN(
        n21938) );
  OAI221_X1 U21009 ( .B1(n21117), .B2(n25241), .C1(n20353), .C2(n25235), .A(
        n21946), .ZN(n21943) );
  AOI22_X1 U21010 ( .A1(n25229), .A2(n24403), .B1(n25223), .B2(n17560), .ZN(
        n21946) );
  OAI221_X1 U21011 ( .B1(n9433), .B2(n25343), .C1(n20416), .C2(n25337), .A(
        n21920), .ZN(n21917) );
  AOI22_X1 U21012 ( .A1(n25331), .A2(n24063), .B1(n25325), .B2(n17526), .ZN(
        n21920) );
  OAI221_X1 U21013 ( .B1(n21116), .B2(n25241), .C1(n20352), .C2(n25235), .A(
        n21928), .ZN(n21925) );
  AOI22_X1 U21014 ( .A1(n25229), .A2(n24405), .B1(n25223), .B2(n17539), .ZN(
        n21928) );
  OAI221_X1 U21015 ( .B1(n9432), .B2(n25343), .C1(n20415), .C2(n25337), .A(
        n21902), .ZN(n21899) );
  AOI22_X1 U21016 ( .A1(n25331), .A2(n24064), .B1(n25325), .B2(n17505), .ZN(
        n21902) );
  OAI221_X1 U21017 ( .B1(n21115), .B2(n25241), .C1(n20351), .C2(n25235), .A(
        n21910), .ZN(n21907) );
  AOI22_X1 U21018 ( .A1(n25229), .A2(n24407), .B1(n25223), .B2(n17518), .ZN(
        n21910) );
  OAI221_X1 U21019 ( .B1(n9431), .B2(n25343), .C1(n20414), .C2(n25337), .A(
        n21884), .ZN(n21881) );
  AOI22_X1 U21020 ( .A1(n25331), .A2(n24065), .B1(n25325), .B2(n17484), .ZN(
        n21884) );
  OAI221_X1 U21021 ( .B1(n21114), .B2(n25241), .C1(n20350), .C2(n25235), .A(
        n21892), .ZN(n21889) );
  AOI22_X1 U21022 ( .A1(n25229), .A2(n24409), .B1(n25223), .B2(n17497), .ZN(
        n21892) );
  OAI221_X1 U21023 ( .B1(n9430), .B2(n25344), .C1(n20413), .C2(n25338), .A(
        n21866), .ZN(n21863) );
  AOI22_X1 U21024 ( .A1(n25332), .A2(n24066), .B1(n25326), .B2(n17463), .ZN(
        n21866) );
  OAI221_X1 U21025 ( .B1(n21113), .B2(n25242), .C1(n20349), .C2(n25236), .A(
        n21874), .ZN(n21871) );
  AOI22_X1 U21026 ( .A1(n25230), .A2(n24411), .B1(n25224), .B2(n17476), .ZN(
        n21874) );
  OAI221_X1 U21027 ( .B1(n9429), .B2(n25344), .C1(n20412), .C2(n25338), .A(
        n21848), .ZN(n21845) );
  AOI22_X1 U21028 ( .A1(n25332), .A2(n24067), .B1(n25326), .B2(n17442), .ZN(
        n21848) );
  OAI221_X1 U21029 ( .B1(n21112), .B2(n25242), .C1(n20348), .C2(n25236), .A(
        n21856), .ZN(n21853) );
  AOI22_X1 U21030 ( .A1(n25230), .A2(n24413), .B1(n25224), .B2(n17455), .ZN(
        n21856) );
  OAI221_X1 U21031 ( .B1(n9428), .B2(n25344), .C1(n20411), .C2(n25338), .A(
        n21830), .ZN(n21827) );
  AOI22_X1 U21032 ( .A1(n25332), .A2(n24068), .B1(n25326), .B2(n17421), .ZN(
        n21830) );
  OAI221_X1 U21033 ( .B1(n21111), .B2(n25242), .C1(n20347), .C2(n25236), .A(
        n21838), .ZN(n21835) );
  AOI22_X1 U21034 ( .A1(n25230), .A2(n24415), .B1(n25224), .B2(n17434), .ZN(
        n21838) );
  OAI221_X1 U21035 ( .B1(n9427), .B2(n25344), .C1(n20410), .C2(n25338), .A(
        n21812), .ZN(n21809) );
  AOI22_X1 U21036 ( .A1(n25332), .A2(n24069), .B1(n25326), .B2(n17400), .ZN(
        n21812) );
  OAI221_X1 U21037 ( .B1(n21110), .B2(n25242), .C1(n20346), .C2(n25236), .A(
        n21820), .ZN(n21817) );
  AOI22_X1 U21038 ( .A1(n25230), .A2(n24417), .B1(n25224), .B2(n17413), .ZN(
        n21820) );
  OAI221_X1 U21039 ( .B1(n9426), .B2(n25344), .C1(n20409), .C2(n25338), .A(
        n21794), .ZN(n21791) );
  AOI22_X1 U21040 ( .A1(n25332), .A2(n24070), .B1(n25326), .B2(n17379), .ZN(
        n21794) );
  OAI221_X1 U21041 ( .B1(n21109), .B2(n25242), .C1(n20345), .C2(n25236), .A(
        n21802), .ZN(n21799) );
  AOI22_X1 U21042 ( .A1(n25230), .A2(n24419), .B1(n25224), .B2(n17392), .ZN(
        n21802) );
  OAI221_X1 U21043 ( .B1(n9425), .B2(n25344), .C1(n20408), .C2(n25338), .A(
        n21776), .ZN(n21773) );
  AOI22_X1 U21044 ( .A1(n25332), .A2(n24071), .B1(n25326), .B2(n17358), .ZN(
        n21776) );
  OAI221_X1 U21045 ( .B1(n21108), .B2(n25242), .C1(n20344), .C2(n25236), .A(
        n21784), .ZN(n21781) );
  AOI22_X1 U21046 ( .A1(n25230), .A2(n24421), .B1(n25224), .B2(n17371), .ZN(
        n21784) );
  OAI221_X1 U21047 ( .B1(n9424), .B2(n25344), .C1(n20407), .C2(n25338), .A(
        n21758), .ZN(n21755) );
  AOI22_X1 U21048 ( .A1(n25332), .A2(n24072), .B1(n25326), .B2(n17337), .ZN(
        n21758) );
  OAI221_X1 U21049 ( .B1(n21107), .B2(n25242), .C1(n20343), .C2(n25236), .A(
        n21766), .ZN(n21763) );
  AOI22_X1 U21050 ( .A1(n25230), .A2(n24423), .B1(n25224), .B2(n17350), .ZN(
        n21766) );
  OAI221_X1 U21051 ( .B1(n9423), .B2(n25344), .C1(n20406), .C2(n25338), .A(
        n21740), .ZN(n21737) );
  AOI22_X1 U21052 ( .A1(n25332), .A2(n24073), .B1(n25326), .B2(n17316), .ZN(
        n21740) );
  OAI221_X1 U21053 ( .B1(n21106), .B2(n25242), .C1(n20342), .C2(n25236), .A(
        n21748), .ZN(n21745) );
  AOI22_X1 U21054 ( .A1(n25230), .A2(n24425), .B1(n25224), .B2(n17329), .ZN(
        n21748) );
  OAI221_X1 U21055 ( .B1(n9422), .B2(n25344), .C1(n20405), .C2(n25338), .A(
        n21722), .ZN(n21719) );
  AOI22_X1 U21056 ( .A1(n25332), .A2(n24074), .B1(n25326), .B2(n17295), .ZN(
        n21722) );
  OAI221_X1 U21057 ( .B1(n21105), .B2(n25242), .C1(n20341), .C2(n25236), .A(
        n21730), .ZN(n21727) );
  AOI22_X1 U21058 ( .A1(n25230), .A2(n24427), .B1(n25224), .B2(n17308), .ZN(
        n21730) );
  OAI221_X1 U21059 ( .B1(n9421), .B2(n25344), .C1(n20404), .C2(n25338), .A(
        n21704), .ZN(n21701) );
  AOI22_X1 U21060 ( .A1(n25332), .A2(n24075), .B1(n25326), .B2(n17274), .ZN(
        n21704) );
  OAI221_X1 U21061 ( .B1(n21104), .B2(n25242), .C1(n20340), .C2(n25236), .A(
        n21712), .ZN(n21709) );
  AOI22_X1 U21062 ( .A1(n25230), .A2(n24429), .B1(n25224), .B2(n17287), .ZN(
        n21712) );
  OAI221_X1 U21063 ( .B1(n9420), .B2(n25344), .C1(n20403), .C2(n25338), .A(
        n21686), .ZN(n21683) );
  AOI22_X1 U21064 ( .A1(n25332), .A2(n24076), .B1(n25326), .B2(n17253), .ZN(
        n21686) );
  OAI221_X1 U21065 ( .B1(n21103), .B2(n25242), .C1(n20339), .C2(n25236), .A(
        n21694), .ZN(n21691) );
  AOI22_X1 U21066 ( .A1(n25230), .A2(n24431), .B1(n25224), .B2(n17266), .ZN(
        n21694) );
  OAI221_X1 U21067 ( .B1(n9419), .B2(n25344), .C1(n20402), .C2(n25338), .A(
        n21668), .ZN(n21665) );
  AOI22_X1 U21068 ( .A1(n25332), .A2(n24077), .B1(n25326), .B2(n17232), .ZN(
        n21668) );
  OAI221_X1 U21069 ( .B1(n21102), .B2(n25242), .C1(n20338), .C2(n25236), .A(
        n21676), .ZN(n21673) );
  AOI22_X1 U21070 ( .A1(n25230), .A2(n24433), .B1(n25224), .B2(n17245), .ZN(
        n21676) );
  OAI221_X1 U21071 ( .B1(n9415), .B2(n25147), .C1(n20398), .C2(n25141), .A(
        n22766), .ZN(n22757) );
  AOI22_X1 U21072 ( .A1(n25135), .A2(n23957), .B1(n25129), .B2(n17148), .ZN(
        n22766) );
  OAI221_X1 U21073 ( .B1(n21094), .B2(n25045), .C1(n20334), .C2(n25039), .A(
        n22791), .ZN(n22782) );
  AOI22_X1 U21074 ( .A1(n25033), .A2(n24441), .B1(n25027), .B2(n17161), .ZN(
        n22791) );
  OAI221_X1 U21075 ( .B1(n9418), .B2(n25147), .C1(n20401), .C2(n25141), .A(
        n22847), .ZN(n22844) );
  AOI22_X1 U21076 ( .A1(n25135), .A2(n23954), .B1(n25129), .B2(n17211), .ZN(
        n22847) );
  OAI221_X1 U21077 ( .B1(n21097), .B2(n25045), .C1(n20337), .C2(n25039), .A(
        n22855), .ZN(n22852) );
  AOI22_X1 U21078 ( .A1(n25033), .A2(n24435), .B1(n25027), .B2(n17224), .ZN(
        n22855) );
  OAI221_X1 U21079 ( .B1(n9417), .B2(n25147), .C1(n20400), .C2(n25141), .A(
        n22829), .ZN(n22826) );
  AOI22_X1 U21080 ( .A1(n25135), .A2(n23955), .B1(n25129), .B2(n17190), .ZN(
        n22829) );
  OAI221_X1 U21081 ( .B1(n21096), .B2(n25045), .C1(n20336), .C2(n25039), .A(
        n22837), .ZN(n22834) );
  AOI22_X1 U21082 ( .A1(n25033), .A2(n24437), .B1(n25027), .B2(n17203), .ZN(
        n22837) );
  OAI221_X1 U21083 ( .B1(n9416), .B2(n25147), .C1(n20399), .C2(n25141), .A(
        n22811), .ZN(n22808) );
  AOI22_X1 U21084 ( .A1(n25135), .A2(n23956), .B1(n25129), .B2(n17169), .ZN(
        n22811) );
  OAI221_X1 U21085 ( .B1(n21095), .B2(n25045), .C1(n20335), .C2(n25039), .A(
        n22819), .ZN(n22816) );
  AOI22_X1 U21086 ( .A1(n25033), .A2(n24439), .B1(n25027), .B2(n17182), .ZN(
        n22819) );
  OAI221_X1 U21087 ( .B1(n9418), .B2(n25345), .C1(n20401), .C2(n25339), .A(
        n21650), .ZN(n21647) );
  AOI22_X1 U21088 ( .A1(n25333), .A2(n23954), .B1(n25327), .B2(n17211), .ZN(
        n21650) );
  OAI221_X1 U21089 ( .B1(n21097), .B2(n25243), .C1(n20337), .C2(n25237), .A(
        n21658), .ZN(n21655) );
  AOI22_X1 U21090 ( .A1(n25231), .A2(n24435), .B1(n25225), .B2(n17224), .ZN(
        n21658) );
  OAI221_X1 U21091 ( .B1(n9417), .B2(n25345), .C1(n20400), .C2(n25339), .A(
        n21632), .ZN(n21629) );
  AOI22_X1 U21092 ( .A1(n25333), .A2(n23955), .B1(n25327), .B2(n17190), .ZN(
        n21632) );
  OAI221_X1 U21093 ( .B1(n21096), .B2(n25243), .C1(n20336), .C2(n25237), .A(
        n21640), .ZN(n21637) );
  AOI22_X1 U21094 ( .A1(n25231), .A2(n24437), .B1(n25225), .B2(n17203), .ZN(
        n21640) );
  OAI221_X1 U21095 ( .B1(n9416), .B2(n25345), .C1(n20399), .C2(n25339), .A(
        n21614), .ZN(n21611) );
  AOI22_X1 U21096 ( .A1(n25333), .A2(n23956), .B1(n25327), .B2(n17169), .ZN(
        n21614) );
  OAI221_X1 U21097 ( .B1(n21095), .B2(n25243), .C1(n20335), .C2(n25237), .A(
        n21622), .ZN(n21619) );
  AOI22_X1 U21098 ( .A1(n25231), .A2(n24439), .B1(n25225), .B2(n17182), .ZN(
        n21622) );
  OAI221_X1 U21099 ( .B1(n9415), .B2(n25345), .C1(n20398), .C2(n25339), .A(
        n21569), .ZN(n21560) );
  AOI22_X1 U21100 ( .A1(n25333), .A2(n23957), .B1(n25327), .B2(n17148), .ZN(
        n21569) );
  OAI221_X1 U21101 ( .B1(n21094), .B2(n25243), .C1(n20334), .C2(n25237), .A(
        n21594), .ZN(n21585) );
  AOI22_X1 U21102 ( .A1(n25231), .A2(n24441), .B1(n25225), .B2(n17161), .ZN(
        n21594) );
  OAI221_X1 U21103 ( .B1(n9478), .B2(n25142), .C1(n20461), .C2(n25136), .A(
        n23932), .ZN(n23924) );
  AOI22_X1 U21104 ( .A1(n25130), .A2(n24018), .B1(n25124), .B2(n18471), .ZN(
        n23932) );
  OAI221_X1 U21105 ( .B1(n9477), .B2(n25142), .C1(n20460), .C2(n25136), .A(
        n23909), .ZN(n23906) );
  AOI22_X1 U21106 ( .A1(n25130), .A2(n24019), .B1(n25124), .B2(n18450), .ZN(
        n23909) );
  OAI221_X1 U21107 ( .B1(n9476), .B2(n25142), .C1(n20459), .C2(n25136), .A(
        n23891), .ZN(n23888) );
  AOI22_X1 U21108 ( .A1(n25130), .A2(n24020), .B1(n25124), .B2(n18429), .ZN(
        n23891) );
  OAI221_X1 U21109 ( .B1(n9475), .B2(n25142), .C1(n20458), .C2(n25136), .A(
        n23873), .ZN(n23870) );
  AOI22_X1 U21110 ( .A1(n25130), .A2(n24021), .B1(n25124), .B2(n18408), .ZN(
        n23873) );
  OAI221_X1 U21111 ( .B1(n9474), .B2(n25142), .C1(n20457), .C2(n25136), .A(
        n23855), .ZN(n23852) );
  AOI22_X1 U21112 ( .A1(n25130), .A2(n24022), .B1(n25124), .B2(n18387), .ZN(
        n23855) );
  OAI221_X1 U21113 ( .B1(n9473), .B2(n25142), .C1(n20456), .C2(n25136), .A(
        n23837), .ZN(n23834) );
  AOI22_X1 U21114 ( .A1(n25130), .A2(n24023), .B1(n25124), .B2(n18366), .ZN(
        n23837) );
  OAI221_X1 U21115 ( .B1(n9472), .B2(n25142), .C1(n20455), .C2(n25136), .A(
        n23819), .ZN(n23816) );
  AOI22_X1 U21116 ( .A1(n25130), .A2(n24024), .B1(n25124), .B2(n18345), .ZN(
        n23819) );
  OAI221_X1 U21117 ( .B1(n9471), .B2(n25142), .C1(n20454), .C2(n25136), .A(
        n23801), .ZN(n23798) );
  AOI22_X1 U21118 ( .A1(n25130), .A2(n24025), .B1(n25124), .B2(n18324), .ZN(
        n23801) );
  OAI221_X1 U21119 ( .B1(n9470), .B2(n25142), .C1(n20453), .C2(n25136), .A(
        n23783), .ZN(n23780) );
  AOI22_X1 U21120 ( .A1(n25130), .A2(n24026), .B1(n25124), .B2(n18303), .ZN(
        n23783) );
  OAI221_X1 U21121 ( .B1(n9469), .B2(n25142), .C1(n20452), .C2(n25136), .A(
        n23765), .ZN(n23762) );
  AOI22_X1 U21122 ( .A1(n25130), .A2(n24027), .B1(n25124), .B2(n18282), .ZN(
        n23765) );
  OAI221_X1 U21123 ( .B1(n9468), .B2(n25142), .C1(n20451), .C2(n25136), .A(
        n23747), .ZN(n23744) );
  AOI22_X1 U21124 ( .A1(n25130), .A2(n24028), .B1(n25124), .B2(n18261), .ZN(
        n23747) );
  OAI221_X1 U21125 ( .B1(n9467), .B2(n25142), .C1(n20450), .C2(n25136), .A(
        n23729), .ZN(n23726) );
  AOI22_X1 U21126 ( .A1(n25130), .A2(n24029), .B1(n25124), .B2(n18240), .ZN(
        n23729) );
  OAI221_X1 U21127 ( .B1(n9478), .B2(n25340), .C1(n20461), .C2(n25334), .A(
        n22735), .ZN(n22727) );
  AOI22_X1 U21128 ( .A1(n25328), .A2(n24018), .B1(n25322), .B2(n18471), .ZN(
        n22735) );
  OAI221_X1 U21129 ( .B1(n9477), .B2(n25340), .C1(n20460), .C2(n25334), .A(
        n22712), .ZN(n22709) );
  AOI22_X1 U21130 ( .A1(n25328), .A2(n24019), .B1(n25322), .B2(n18450), .ZN(
        n22712) );
  OAI221_X1 U21131 ( .B1(n9476), .B2(n25340), .C1(n20459), .C2(n25334), .A(
        n22694), .ZN(n22691) );
  AOI22_X1 U21132 ( .A1(n25328), .A2(n24020), .B1(n25322), .B2(n18429), .ZN(
        n22694) );
  OAI221_X1 U21133 ( .B1(n9475), .B2(n25340), .C1(n20458), .C2(n25334), .A(
        n22676), .ZN(n22673) );
  AOI22_X1 U21134 ( .A1(n25328), .A2(n24021), .B1(n25322), .B2(n18408), .ZN(
        n22676) );
  OAI221_X1 U21135 ( .B1(n9474), .B2(n25340), .C1(n20457), .C2(n25334), .A(
        n22658), .ZN(n22655) );
  AOI22_X1 U21136 ( .A1(n25328), .A2(n24022), .B1(n25322), .B2(n18387), .ZN(
        n22658) );
  OAI221_X1 U21137 ( .B1(n9473), .B2(n25340), .C1(n20456), .C2(n25334), .A(
        n22640), .ZN(n22637) );
  AOI22_X1 U21138 ( .A1(n25328), .A2(n24023), .B1(n25322), .B2(n18366), .ZN(
        n22640) );
  OAI221_X1 U21139 ( .B1(n9472), .B2(n25340), .C1(n20455), .C2(n25334), .A(
        n22622), .ZN(n22619) );
  AOI22_X1 U21140 ( .A1(n25328), .A2(n24024), .B1(n25322), .B2(n18345), .ZN(
        n22622) );
  OAI221_X1 U21141 ( .B1(n9471), .B2(n25340), .C1(n20454), .C2(n25334), .A(
        n22604), .ZN(n22601) );
  AOI22_X1 U21142 ( .A1(n25328), .A2(n24025), .B1(n25322), .B2(n18324), .ZN(
        n22604) );
  OAI221_X1 U21143 ( .B1(n9470), .B2(n25340), .C1(n20453), .C2(n25334), .A(
        n22586), .ZN(n22583) );
  AOI22_X1 U21144 ( .A1(n25328), .A2(n24026), .B1(n25322), .B2(n18303), .ZN(
        n22586) );
  OAI221_X1 U21145 ( .B1(n9469), .B2(n25340), .C1(n20452), .C2(n25334), .A(
        n22568), .ZN(n22565) );
  AOI22_X1 U21146 ( .A1(n25328), .A2(n24027), .B1(n25322), .B2(n18282), .ZN(
        n22568) );
  OAI221_X1 U21147 ( .B1(n9468), .B2(n25340), .C1(n20451), .C2(n25334), .A(
        n22550), .ZN(n22547) );
  AOI22_X1 U21148 ( .A1(n25328), .A2(n24028), .B1(n25322), .B2(n18261), .ZN(
        n22550) );
  OAI221_X1 U21149 ( .B1(n9467), .B2(n25340), .C1(n20450), .C2(n25334), .A(
        n22532), .ZN(n22529) );
  AOI22_X1 U21150 ( .A1(n25328), .A2(n24029), .B1(n25322), .B2(n18240), .ZN(
        n22532) );
  OAI221_X1 U21151 ( .B1(n21161), .B2(n25040), .C1(n20397), .C2(n25034), .A(
        n23947), .ZN(n23943) );
  AOI22_X1 U21152 ( .A1(n25028), .A2(n24443), .B1(n25022), .B2(n18484), .ZN(
        n23947) );
  OAI221_X1 U21153 ( .B1(n21160), .B2(n25040), .C1(n20396), .C2(n25034), .A(
        n23917), .ZN(n23914) );
  AOI22_X1 U21154 ( .A1(n25028), .A2(n24445), .B1(n25022), .B2(n18463), .ZN(
        n23917) );
  OAI221_X1 U21155 ( .B1(n21159), .B2(n25040), .C1(n20395), .C2(n25034), .A(
        n23899), .ZN(n23896) );
  AOI22_X1 U21156 ( .A1(n25028), .A2(n24447), .B1(n25022), .B2(n18442), .ZN(
        n23899) );
  OAI221_X1 U21157 ( .B1(n21158), .B2(n25040), .C1(n20394), .C2(n25034), .A(
        n23881), .ZN(n23878) );
  AOI22_X1 U21158 ( .A1(n25028), .A2(n24449), .B1(n25022), .B2(n18421), .ZN(
        n23881) );
  OAI221_X1 U21159 ( .B1(n21157), .B2(n25040), .C1(n20393), .C2(n25034), .A(
        n23863), .ZN(n23860) );
  AOI22_X1 U21160 ( .A1(n25028), .A2(n24451), .B1(n25022), .B2(n18400), .ZN(
        n23863) );
  OAI221_X1 U21161 ( .B1(n21156), .B2(n25040), .C1(n20392), .C2(n25034), .A(
        n23845), .ZN(n23842) );
  AOI22_X1 U21162 ( .A1(n25028), .A2(n24453), .B1(n25022), .B2(n18379), .ZN(
        n23845) );
  OAI221_X1 U21163 ( .B1(n21155), .B2(n25040), .C1(n20391), .C2(n25034), .A(
        n23827), .ZN(n23824) );
  AOI22_X1 U21164 ( .A1(n25028), .A2(n24455), .B1(n25022), .B2(n18358), .ZN(
        n23827) );
  OAI221_X1 U21165 ( .B1(n21154), .B2(n25040), .C1(n20390), .C2(n25034), .A(
        n23809), .ZN(n23806) );
  AOI22_X1 U21166 ( .A1(n25028), .A2(n24457), .B1(n25022), .B2(n18337), .ZN(
        n23809) );
  OAI221_X1 U21167 ( .B1(n21153), .B2(n25040), .C1(n20389), .C2(n25034), .A(
        n23791), .ZN(n23788) );
  AOI22_X1 U21168 ( .A1(n25028), .A2(n24459), .B1(n25022), .B2(n18316), .ZN(
        n23791) );
  OAI221_X1 U21169 ( .B1(n21152), .B2(n25040), .C1(n20388), .C2(n25034), .A(
        n23773), .ZN(n23770) );
  AOI22_X1 U21170 ( .A1(n25028), .A2(n24461), .B1(n25022), .B2(n18295), .ZN(
        n23773) );
  OAI221_X1 U21171 ( .B1(n21151), .B2(n25040), .C1(n20387), .C2(n25034), .A(
        n23755), .ZN(n23752) );
  AOI22_X1 U21172 ( .A1(n25028), .A2(n24463), .B1(n25022), .B2(n18274), .ZN(
        n23755) );
  OAI221_X1 U21173 ( .B1(n21150), .B2(n25040), .C1(n20386), .C2(n25034), .A(
        n23737), .ZN(n23734) );
  AOI22_X1 U21174 ( .A1(n25028), .A2(n24465), .B1(n25022), .B2(n18253), .ZN(
        n23737) );
  OAI221_X1 U21175 ( .B1(n21161), .B2(n25238), .C1(n20397), .C2(n25232), .A(
        n22750), .ZN(n22746) );
  AOI22_X1 U21176 ( .A1(n25226), .A2(n24443), .B1(n25220), .B2(n18484), .ZN(
        n22750) );
  OAI221_X1 U21177 ( .B1(n21160), .B2(n25238), .C1(n20396), .C2(n25232), .A(
        n22720), .ZN(n22717) );
  AOI22_X1 U21178 ( .A1(n25226), .A2(n24445), .B1(n25220), .B2(n18463), .ZN(
        n22720) );
  OAI221_X1 U21179 ( .B1(n21159), .B2(n25238), .C1(n20395), .C2(n25232), .A(
        n22702), .ZN(n22699) );
  AOI22_X1 U21180 ( .A1(n25226), .A2(n24447), .B1(n25220), .B2(n18442), .ZN(
        n22702) );
  OAI221_X1 U21181 ( .B1(n21158), .B2(n25238), .C1(n20394), .C2(n25232), .A(
        n22684), .ZN(n22681) );
  AOI22_X1 U21182 ( .A1(n25226), .A2(n24449), .B1(n25220), .B2(n18421), .ZN(
        n22684) );
  OAI221_X1 U21183 ( .B1(n21157), .B2(n25238), .C1(n20393), .C2(n25232), .A(
        n22666), .ZN(n22663) );
  AOI22_X1 U21184 ( .A1(n25226), .A2(n24451), .B1(n25220), .B2(n18400), .ZN(
        n22666) );
  OAI221_X1 U21185 ( .B1(n21156), .B2(n25238), .C1(n20392), .C2(n25232), .A(
        n22648), .ZN(n22645) );
  AOI22_X1 U21186 ( .A1(n25226), .A2(n24453), .B1(n25220), .B2(n18379), .ZN(
        n22648) );
  OAI221_X1 U21187 ( .B1(n21155), .B2(n25238), .C1(n20391), .C2(n25232), .A(
        n22630), .ZN(n22627) );
  AOI22_X1 U21188 ( .A1(n25226), .A2(n24455), .B1(n25220), .B2(n18358), .ZN(
        n22630) );
  OAI221_X1 U21189 ( .B1(n21154), .B2(n25238), .C1(n20390), .C2(n25232), .A(
        n22612), .ZN(n22609) );
  AOI22_X1 U21190 ( .A1(n25226), .A2(n24457), .B1(n25220), .B2(n18337), .ZN(
        n22612) );
  OAI221_X1 U21191 ( .B1(n21153), .B2(n25238), .C1(n20389), .C2(n25232), .A(
        n22594), .ZN(n22591) );
  AOI22_X1 U21192 ( .A1(n25226), .A2(n24459), .B1(n25220), .B2(n18316), .ZN(
        n22594) );
  OAI221_X1 U21193 ( .B1(n21152), .B2(n25238), .C1(n20388), .C2(n25232), .A(
        n22576), .ZN(n22573) );
  AOI22_X1 U21194 ( .A1(n25226), .A2(n24461), .B1(n25220), .B2(n18295), .ZN(
        n22576) );
  OAI221_X1 U21195 ( .B1(n21151), .B2(n25238), .C1(n20387), .C2(n25232), .A(
        n22558), .ZN(n22555) );
  AOI22_X1 U21196 ( .A1(n25226), .A2(n24463), .B1(n25220), .B2(n18274), .ZN(
        n22558) );
  OAI221_X1 U21197 ( .B1(n21150), .B2(n25238), .C1(n20386), .C2(n25232), .A(
        n22540), .ZN(n22537) );
  AOI22_X1 U21198 ( .A1(n25226), .A2(n24465), .B1(n25220), .B2(n18253), .ZN(
        n22540) );
  OAI221_X1 U21199 ( .B1(n21401), .B2(n25017), .C1(n20321), .C2(n25011), .A(
        n23720), .ZN(n23715) );
  AOI22_X1 U21200 ( .A1(n25005), .A2(n24626), .B1(n24999), .B2(n18234), .ZN(
        n23720) );
  OAI221_X1 U21201 ( .B1(n21400), .B2(n25017), .C1(n20320), .C2(n25011), .A(
        n23702), .ZN(n23697) );
  AOI22_X1 U21202 ( .A1(n25005), .A2(n24627), .B1(n24999), .B2(n18213), .ZN(
        n23702) );
  OAI221_X1 U21203 ( .B1(n21399), .B2(n25017), .C1(n20319), .C2(n25011), .A(
        n23684), .ZN(n23679) );
  AOI22_X1 U21204 ( .A1(n25005), .A2(n24628), .B1(n24999), .B2(n18192), .ZN(
        n23684) );
  OAI221_X1 U21205 ( .B1(n21398), .B2(n25017), .C1(n20318), .C2(n25011), .A(
        n23666), .ZN(n23661) );
  AOI22_X1 U21206 ( .A1(n25005), .A2(n24629), .B1(n24999), .B2(n18171), .ZN(
        n23666) );
  OAI221_X1 U21207 ( .B1(n21397), .B2(n25017), .C1(n20317), .C2(n25011), .A(
        n23648), .ZN(n23643) );
  AOI22_X1 U21208 ( .A1(n25005), .A2(n24630), .B1(n24999), .B2(n18150), .ZN(
        n23648) );
  OAI221_X1 U21209 ( .B1(n21396), .B2(n25017), .C1(n20316), .C2(n25011), .A(
        n23630), .ZN(n23625) );
  AOI22_X1 U21210 ( .A1(n25005), .A2(n24631), .B1(n24999), .B2(n18129), .ZN(
        n23630) );
  OAI221_X1 U21211 ( .B1(n21395), .B2(n25017), .C1(n20315), .C2(n25011), .A(
        n23612), .ZN(n23607) );
  AOI22_X1 U21212 ( .A1(n25005), .A2(n24632), .B1(n24999), .B2(n18108), .ZN(
        n23612) );
  OAI221_X1 U21213 ( .B1(n21394), .B2(n25017), .C1(n20314), .C2(n25011), .A(
        n23594), .ZN(n23589) );
  AOI22_X1 U21214 ( .A1(n25005), .A2(n24633), .B1(n24999), .B2(n18087), .ZN(
        n23594) );
  OAI221_X1 U21215 ( .B1(n21393), .B2(n25017), .C1(n20313), .C2(n25011), .A(
        n23576), .ZN(n23571) );
  AOI22_X1 U21216 ( .A1(n25005), .A2(n24634), .B1(n24999), .B2(n18066), .ZN(
        n23576) );
  OAI221_X1 U21217 ( .B1(n21392), .B2(n25017), .C1(n20312), .C2(n25011), .A(
        n23558), .ZN(n23553) );
  AOI22_X1 U21218 ( .A1(n25005), .A2(n24635), .B1(n24999), .B2(n18045), .ZN(
        n23558) );
  OAI221_X1 U21219 ( .B1(n21391), .B2(n25017), .C1(n20311), .C2(n25011), .A(
        n23540), .ZN(n23535) );
  AOI22_X1 U21220 ( .A1(n25005), .A2(n24636), .B1(n24999), .B2(n18024), .ZN(
        n23540) );
  OAI221_X1 U21221 ( .B1(n21390), .B2(n25017), .C1(n20310), .C2(n25011), .A(
        n23522), .ZN(n23517) );
  AOI22_X1 U21222 ( .A1(n25005), .A2(n24637), .B1(n24999), .B2(n18003), .ZN(
        n23522) );
  OAI221_X1 U21223 ( .B1(n21389), .B2(n25018), .C1(n20309), .C2(n25012), .A(
        n23504), .ZN(n23499) );
  AOI22_X1 U21224 ( .A1(n25006), .A2(n24638), .B1(n25000), .B2(n17982), .ZN(
        n23504) );
  OAI221_X1 U21225 ( .B1(n21388), .B2(n25018), .C1(n20308), .C2(n25012), .A(
        n23486), .ZN(n23481) );
  AOI22_X1 U21226 ( .A1(n25006), .A2(n24639), .B1(n25000), .B2(n17961), .ZN(
        n23486) );
  OAI221_X1 U21227 ( .B1(n21387), .B2(n25018), .C1(n20307), .C2(n25012), .A(
        n23468), .ZN(n23463) );
  AOI22_X1 U21228 ( .A1(n25006), .A2(n24640), .B1(n25000), .B2(n17940), .ZN(
        n23468) );
  OAI221_X1 U21229 ( .B1(n21386), .B2(n25018), .C1(n20306), .C2(n25012), .A(
        n23450), .ZN(n23445) );
  AOI22_X1 U21230 ( .A1(n25006), .A2(n24641), .B1(n25000), .B2(n17919), .ZN(
        n23450) );
  OAI221_X1 U21231 ( .B1(n21385), .B2(n25018), .C1(n20305), .C2(n25012), .A(
        n23432), .ZN(n23427) );
  AOI22_X1 U21232 ( .A1(n25006), .A2(n24642), .B1(n25000), .B2(n17898), .ZN(
        n23432) );
  OAI221_X1 U21233 ( .B1(n21384), .B2(n25018), .C1(n20304), .C2(n25012), .A(
        n23414), .ZN(n23409) );
  AOI22_X1 U21234 ( .A1(n25006), .A2(n24643), .B1(n25000), .B2(n17877), .ZN(
        n23414) );
  OAI221_X1 U21235 ( .B1(n21383), .B2(n25018), .C1(n20303), .C2(n25012), .A(
        n23396), .ZN(n23391) );
  AOI22_X1 U21236 ( .A1(n25006), .A2(n24644), .B1(n25000), .B2(n17856), .ZN(
        n23396) );
  OAI221_X1 U21237 ( .B1(n21382), .B2(n25018), .C1(n20302), .C2(n25012), .A(
        n23378), .ZN(n23373) );
  AOI22_X1 U21238 ( .A1(n25006), .A2(n24645), .B1(n25000), .B2(n17835), .ZN(
        n23378) );
  OAI221_X1 U21239 ( .B1(n21381), .B2(n25018), .C1(n20301), .C2(n25012), .A(
        n23360), .ZN(n23355) );
  AOI22_X1 U21240 ( .A1(n25006), .A2(n24646), .B1(n25000), .B2(n17814), .ZN(
        n23360) );
  OAI221_X1 U21241 ( .B1(n21380), .B2(n25018), .C1(n20300), .C2(n25012), .A(
        n23342), .ZN(n23337) );
  AOI22_X1 U21242 ( .A1(n25006), .A2(n24647), .B1(n25000), .B2(n17793), .ZN(
        n23342) );
  OAI221_X1 U21243 ( .B1(n21379), .B2(n25018), .C1(n20299), .C2(n25012), .A(
        n23324), .ZN(n23319) );
  AOI22_X1 U21244 ( .A1(n25006), .A2(n24648), .B1(n25000), .B2(n17772), .ZN(
        n23324) );
  OAI221_X1 U21245 ( .B1(n21378), .B2(n25018), .C1(n20298), .C2(n25012), .A(
        n23306), .ZN(n23301) );
  AOI22_X1 U21246 ( .A1(n25006), .A2(n24649), .B1(n25000), .B2(n17751), .ZN(
        n23306) );
  OAI221_X1 U21247 ( .B1(n21377), .B2(n25019), .C1(n20297), .C2(n25013), .A(
        n23288), .ZN(n23283) );
  AOI22_X1 U21248 ( .A1(n25007), .A2(n24650), .B1(n25001), .B2(n17730), .ZN(
        n23288) );
  OAI221_X1 U21249 ( .B1(n21376), .B2(n25019), .C1(n20296), .C2(n25013), .A(
        n23270), .ZN(n23265) );
  AOI22_X1 U21250 ( .A1(n25007), .A2(n24651), .B1(n25001), .B2(n17709), .ZN(
        n23270) );
  OAI221_X1 U21251 ( .B1(n21375), .B2(n25019), .C1(n20295), .C2(n25013), .A(
        n23252), .ZN(n23247) );
  AOI22_X1 U21252 ( .A1(n25007), .A2(n24652), .B1(n25001), .B2(n17688), .ZN(
        n23252) );
  OAI221_X1 U21253 ( .B1(n21374), .B2(n25019), .C1(n20294), .C2(n25013), .A(
        n23234), .ZN(n23229) );
  AOI22_X1 U21254 ( .A1(n25007), .A2(n24653), .B1(n25001), .B2(n17667), .ZN(
        n23234) );
  OAI221_X1 U21255 ( .B1(n21373), .B2(n25019), .C1(n20293), .C2(n25013), .A(
        n23216), .ZN(n23211) );
  AOI22_X1 U21256 ( .A1(n25007), .A2(n24654), .B1(n25001), .B2(n17646), .ZN(
        n23216) );
  OAI221_X1 U21257 ( .B1(n21372), .B2(n25019), .C1(n20292), .C2(n25013), .A(
        n23198), .ZN(n23193) );
  AOI22_X1 U21258 ( .A1(n25007), .A2(n24655), .B1(n25001), .B2(n17625), .ZN(
        n23198) );
  OAI221_X1 U21259 ( .B1(n21371), .B2(n25019), .C1(n20291), .C2(n25013), .A(
        n23180), .ZN(n23175) );
  AOI22_X1 U21260 ( .A1(n25007), .A2(n24656), .B1(n25001), .B2(n17604), .ZN(
        n23180) );
  OAI221_X1 U21261 ( .B1(n21370), .B2(n25019), .C1(n20290), .C2(n25013), .A(
        n23162), .ZN(n23157) );
  AOI22_X1 U21262 ( .A1(n25007), .A2(n24657), .B1(n25001), .B2(n17583), .ZN(
        n23162) );
  OAI221_X1 U21263 ( .B1(n21369), .B2(n25019), .C1(n20289), .C2(n25013), .A(
        n23144), .ZN(n23139) );
  AOI22_X1 U21264 ( .A1(n25007), .A2(n24658), .B1(n25001), .B2(n17562), .ZN(
        n23144) );
  OAI221_X1 U21265 ( .B1(n21368), .B2(n25019), .C1(n20288), .C2(n25013), .A(
        n23126), .ZN(n23121) );
  AOI22_X1 U21266 ( .A1(n25007), .A2(n24659), .B1(n25001), .B2(n17541), .ZN(
        n23126) );
  OAI221_X1 U21267 ( .B1(n21367), .B2(n25019), .C1(n20287), .C2(n25013), .A(
        n23108), .ZN(n23103) );
  AOI22_X1 U21268 ( .A1(n25007), .A2(n24660), .B1(n25001), .B2(n17520), .ZN(
        n23108) );
  OAI221_X1 U21269 ( .B1(n21366), .B2(n25019), .C1(n20286), .C2(n25013), .A(
        n23090), .ZN(n23085) );
  AOI22_X1 U21270 ( .A1(n25007), .A2(n24661), .B1(n25001), .B2(n17499), .ZN(
        n23090) );
  OAI221_X1 U21271 ( .B1(n21365), .B2(n25020), .C1(n20285), .C2(n25014), .A(
        n23072), .ZN(n23067) );
  AOI22_X1 U21272 ( .A1(n25008), .A2(n24662), .B1(n25002), .B2(n17478), .ZN(
        n23072) );
  OAI221_X1 U21273 ( .B1(n21364), .B2(n25020), .C1(n20284), .C2(n25014), .A(
        n23054), .ZN(n23049) );
  AOI22_X1 U21274 ( .A1(n25008), .A2(n24663), .B1(n25002), .B2(n17457), .ZN(
        n23054) );
  OAI221_X1 U21275 ( .B1(n21363), .B2(n25020), .C1(n20283), .C2(n25014), .A(
        n23036), .ZN(n23031) );
  AOI22_X1 U21276 ( .A1(n25008), .A2(n24664), .B1(n25002), .B2(n17436), .ZN(
        n23036) );
  OAI221_X1 U21277 ( .B1(n21362), .B2(n25020), .C1(n20282), .C2(n25014), .A(
        n23018), .ZN(n23013) );
  AOI22_X1 U21278 ( .A1(n25008), .A2(n24665), .B1(n25002), .B2(n17415), .ZN(
        n23018) );
  OAI221_X1 U21279 ( .B1(n21361), .B2(n25020), .C1(n20281), .C2(n25014), .A(
        n23000), .ZN(n22995) );
  AOI22_X1 U21280 ( .A1(n25008), .A2(n24666), .B1(n25002), .B2(n17394), .ZN(
        n23000) );
  OAI221_X1 U21281 ( .B1(n21360), .B2(n25020), .C1(n20280), .C2(n25014), .A(
        n22982), .ZN(n22977) );
  AOI22_X1 U21282 ( .A1(n25008), .A2(n24667), .B1(n25002), .B2(n17373), .ZN(
        n22982) );
  OAI221_X1 U21283 ( .B1(n21359), .B2(n25020), .C1(n20279), .C2(n25014), .A(
        n22964), .ZN(n22959) );
  AOI22_X1 U21284 ( .A1(n25008), .A2(n24668), .B1(n25002), .B2(n17352), .ZN(
        n22964) );
  OAI221_X1 U21285 ( .B1(n21358), .B2(n25020), .C1(n20278), .C2(n25014), .A(
        n22946), .ZN(n22941) );
  AOI22_X1 U21286 ( .A1(n25008), .A2(n24669), .B1(n25002), .B2(n17331), .ZN(
        n22946) );
  OAI221_X1 U21287 ( .B1(n21357), .B2(n25020), .C1(n20277), .C2(n25014), .A(
        n22928), .ZN(n22923) );
  AOI22_X1 U21288 ( .A1(n25008), .A2(n24670), .B1(n25002), .B2(n17310), .ZN(
        n22928) );
  OAI221_X1 U21289 ( .B1(n21356), .B2(n25020), .C1(n20276), .C2(n25014), .A(
        n22910), .ZN(n22905) );
  AOI22_X1 U21290 ( .A1(n25008), .A2(n24671), .B1(n25002), .B2(n17289), .ZN(
        n22910) );
  OAI221_X1 U21291 ( .B1(n21355), .B2(n25020), .C1(n20275), .C2(n25014), .A(
        n22892), .ZN(n22887) );
  AOI22_X1 U21292 ( .A1(n25008), .A2(n24672), .B1(n25002), .B2(n17268), .ZN(
        n22892) );
  OAI221_X1 U21293 ( .B1(n21354), .B2(n25020), .C1(n20274), .C2(n25014), .A(
        n22874), .ZN(n22869) );
  AOI22_X1 U21294 ( .A1(n25008), .A2(n24673), .B1(n25002), .B2(n17247), .ZN(
        n22874) );
  OAI221_X1 U21295 ( .B1(n21401), .B2(n25215), .C1(n20321), .C2(n25209), .A(
        n22523), .ZN(n22518) );
  AOI22_X1 U21296 ( .A1(n25203), .A2(n24626), .B1(n25197), .B2(n18234), .ZN(
        n22523) );
  OAI221_X1 U21297 ( .B1(n21400), .B2(n25215), .C1(n20320), .C2(n25209), .A(
        n22505), .ZN(n22500) );
  AOI22_X1 U21298 ( .A1(n25203), .A2(n24627), .B1(n25197), .B2(n18213), .ZN(
        n22505) );
  OAI221_X1 U21299 ( .B1(n21399), .B2(n25215), .C1(n20319), .C2(n25209), .A(
        n22487), .ZN(n22482) );
  AOI22_X1 U21300 ( .A1(n25203), .A2(n24628), .B1(n25197), .B2(n18192), .ZN(
        n22487) );
  OAI221_X1 U21301 ( .B1(n21398), .B2(n25215), .C1(n20318), .C2(n25209), .A(
        n22469), .ZN(n22464) );
  AOI22_X1 U21302 ( .A1(n25203), .A2(n24629), .B1(n25197), .B2(n18171), .ZN(
        n22469) );
  OAI221_X1 U21303 ( .B1(n21397), .B2(n25215), .C1(n20317), .C2(n25209), .A(
        n22451), .ZN(n22446) );
  AOI22_X1 U21304 ( .A1(n25203), .A2(n24630), .B1(n25197), .B2(n18150), .ZN(
        n22451) );
  OAI221_X1 U21305 ( .B1(n21396), .B2(n25215), .C1(n20316), .C2(n25209), .A(
        n22433), .ZN(n22428) );
  AOI22_X1 U21306 ( .A1(n25203), .A2(n24631), .B1(n25197), .B2(n18129), .ZN(
        n22433) );
  OAI221_X1 U21307 ( .B1(n21395), .B2(n25215), .C1(n20315), .C2(n25209), .A(
        n22415), .ZN(n22410) );
  AOI22_X1 U21308 ( .A1(n25203), .A2(n24632), .B1(n25197), .B2(n18108), .ZN(
        n22415) );
  OAI221_X1 U21309 ( .B1(n21394), .B2(n25215), .C1(n20314), .C2(n25209), .A(
        n22397), .ZN(n22392) );
  AOI22_X1 U21310 ( .A1(n25203), .A2(n24633), .B1(n25197), .B2(n18087), .ZN(
        n22397) );
  OAI221_X1 U21311 ( .B1(n21393), .B2(n25215), .C1(n20313), .C2(n25209), .A(
        n22379), .ZN(n22374) );
  AOI22_X1 U21312 ( .A1(n25203), .A2(n24634), .B1(n25197), .B2(n18066), .ZN(
        n22379) );
  OAI221_X1 U21313 ( .B1(n21392), .B2(n25215), .C1(n20312), .C2(n25209), .A(
        n22361), .ZN(n22356) );
  AOI22_X1 U21314 ( .A1(n25203), .A2(n24635), .B1(n25197), .B2(n18045), .ZN(
        n22361) );
  OAI221_X1 U21315 ( .B1(n21391), .B2(n25215), .C1(n20311), .C2(n25209), .A(
        n22343), .ZN(n22338) );
  AOI22_X1 U21316 ( .A1(n25203), .A2(n24636), .B1(n25197), .B2(n18024), .ZN(
        n22343) );
  OAI221_X1 U21317 ( .B1(n21390), .B2(n25215), .C1(n20310), .C2(n25209), .A(
        n22325), .ZN(n22320) );
  AOI22_X1 U21318 ( .A1(n25203), .A2(n24637), .B1(n25197), .B2(n18003), .ZN(
        n22325) );
  OAI221_X1 U21319 ( .B1(n21389), .B2(n25216), .C1(n20309), .C2(n25210), .A(
        n22307), .ZN(n22302) );
  AOI22_X1 U21320 ( .A1(n25204), .A2(n24638), .B1(n25198), .B2(n17982), .ZN(
        n22307) );
  OAI221_X1 U21321 ( .B1(n21388), .B2(n25216), .C1(n20308), .C2(n25210), .A(
        n22289), .ZN(n22284) );
  AOI22_X1 U21322 ( .A1(n25204), .A2(n24639), .B1(n25198), .B2(n17961), .ZN(
        n22289) );
  OAI221_X1 U21323 ( .B1(n21387), .B2(n25216), .C1(n20307), .C2(n25210), .A(
        n22271), .ZN(n22266) );
  AOI22_X1 U21324 ( .A1(n25204), .A2(n24640), .B1(n25198), .B2(n17940), .ZN(
        n22271) );
  OAI221_X1 U21325 ( .B1(n21386), .B2(n25216), .C1(n20306), .C2(n25210), .A(
        n22253), .ZN(n22248) );
  AOI22_X1 U21326 ( .A1(n25204), .A2(n24641), .B1(n25198), .B2(n17919), .ZN(
        n22253) );
  OAI221_X1 U21327 ( .B1(n21385), .B2(n25216), .C1(n20305), .C2(n25210), .A(
        n22235), .ZN(n22230) );
  AOI22_X1 U21328 ( .A1(n25204), .A2(n24642), .B1(n25198), .B2(n17898), .ZN(
        n22235) );
  OAI221_X1 U21329 ( .B1(n21384), .B2(n25216), .C1(n20304), .C2(n25210), .A(
        n22217), .ZN(n22212) );
  AOI22_X1 U21330 ( .A1(n25204), .A2(n24643), .B1(n25198), .B2(n17877), .ZN(
        n22217) );
  OAI221_X1 U21331 ( .B1(n21383), .B2(n25216), .C1(n20303), .C2(n25210), .A(
        n22199), .ZN(n22194) );
  AOI22_X1 U21332 ( .A1(n25204), .A2(n24644), .B1(n25198), .B2(n17856), .ZN(
        n22199) );
  OAI221_X1 U21333 ( .B1(n21382), .B2(n25216), .C1(n20302), .C2(n25210), .A(
        n22181), .ZN(n22176) );
  AOI22_X1 U21334 ( .A1(n25204), .A2(n24645), .B1(n25198), .B2(n17835), .ZN(
        n22181) );
  OAI221_X1 U21335 ( .B1(n21381), .B2(n25216), .C1(n20301), .C2(n25210), .A(
        n22163), .ZN(n22158) );
  AOI22_X1 U21336 ( .A1(n25204), .A2(n24646), .B1(n25198), .B2(n17814), .ZN(
        n22163) );
  OAI221_X1 U21337 ( .B1(n21380), .B2(n25216), .C1(n20300), .C2(n25210), .A(
        n22145), .ZN(n22140) );
  AOI22_X1 U21338 ( .A1(n25204), .A2(n24647), .B1(n25198), .B2(n17793), .ZN(
        n22145) );
  OAI221_X1 U21339 ( .B1(n21379), .B2(n25216), .C1(n20299), .C2(n25210), .A(
        n22127), .ZN(n22122) );
  AOI22_X1 U21340 ( .A1(n25204), .A2(n24648), .B1(n25198), .B2(n17772), .ZN(
        n22127) );
  OAI221_X1 U21341 ( .B1(n21378), .B2(n25216), .C1(n20298), .C2(n25210), .A(
        n22109), .ZN(n22104) );
  AOI22_X1 U21342 ( .A1(n25204), .A2(n24649), .B1(n25198), .B2(n17751), .ZN(
        n22109) );
  OAI221_X1 U21343 ( .B1(n21377), .B2(n25217), .C1(n20297), .C2(n25211), .A(
        n22091), .ZN(n22086) );
  AOI22_X1 U21344 ( .A1(n25205), .A2(n24650), .B1(n25199), .B2(n17730), .ZN(
        n22091) );
  OAI221_X1 U21345 ( .B1(n21376), .B2(n25217), .C1(n20296), .C2(n25211), .A(
        n22073), .ZN(n22068) );
  AOI22_X1 U21346 ( .A1(n25205), .A2(n24651), .B1(n25199), .B2(n17709), .ZN(
        n22073) );
  OAI221_X1 U21347 ( .B1(n21375), .B2(n25217), .C1(n20295), .C2(n25211), .A(
        n22055), .ZN(n22050) );
  AOI22_X1 U21348 ( .A1(n25205), .A2(n24652), .B1(n25199), .B2(n17688), .ZN(
        n22055) );
  OAI221_X1 U21349 ( .B1(n21374), .B2(n25217), .C1(n20294), .C2(n25211), .A(
        n22037), .ZN(n22032) );
  AOI22_X1 U21350 ( .A1(n25205), .A2(n24653), .B1(n25199), .B2(n17667), .ZN(
        n22037) );
  OAI221_X1 U21351 ( .B1(n21373), .B2(n25217), .C1(n20293), .C2(n25211), .A(
        n22019), .ZN(n22014) );
  AOI22_X1 U21352 ( .A1(n25205), .A2(n24654), .B1(n25199), .B2(n17646), .ZN(
        n22019) );
  OAI221_X1 U21353 ( .B1(n21372), .B2(n25217), .C1(n20292), .C2(n25211), .A(
        n22001), .ZN(n21996) );
  AOI22_X1 U21354 ( .A1(n25205), .A2(n24655), .B1(n25199), .B2(n17625), .ZN(
        n22001) );
  OAI221_X1 U21355 ( .B1(n21371), .B2(n25217), .C1(n20291), .C2(n25211), .A(
        n21983), .ZN(n21978) );
  AOI22_X1 U21356 ( .A1(n25205), .A2(n24656), .B1(n25199), .B2(n17604), .ZN(
        n21983) );
  OAI221_X1 U21357 ( .B1(n21370), .B2(n25217), .C1(n20290), .C2(n25211), .A(
        n21965), .ZN(n21960) );
  AOI22_X1 U21358 ( .A1(n25205), .A2(n24657), .B1(n25199), .B2(n17583), .ZN(
        n21965) );
  OAI221_X1 U21359 ( .B1(n21369), .B2(n25217), .C1(n20289), .C2(n25211), .A(
        n21947), .ZN(n21942) );
  AOI22_X1 U21360 ( .A1(n25205), .A2(n24658), .B1(n25199), .B2(n17562), .ZN(
        n21947) );
  OAI221_X1 U21361 ( .B1(n21368), .B2(n25217), .C1(n20288), .C2(n25211), .A(
        n21929), .ZN(n21924) );
  AOI22_X1 U21362 ( .A1(n25205), .A2(n24659), .B1(n25199), .B2(n17541), .ZN(
        n21929) );
  OAI221_X1 U21363 ( .B1(n21367), .B2(n25217), .C1(n20287), .C2(n25211), .A(
        n21911), .ZN(n21906) );
  AOI22_X1 U21364 ( .A1(n25205), .A2(n24660), .B1(n25199), .B2(n17520), .ZN(
        n21911) );
  OAI221_X1 U21365 ( .B1(n21366), .B2(n25217), .C1(n20286), .C2(n25211), .A(
        n21893), .ZN(n21888) );
  AOI22_X1 U21366 ( .A1(n25205), .A2(n24661), .B1(n25199), .B2(n17499), .ZN(
        n21893) );
  OAI221_X1 U21367 ( .B1(n21365), .B2(n25218), .C1(n20285), .C2(n25212), .A(
        n21875), .ZN(n21870) );
  AOI22_X1 U21368 ( .A1(n25206), .A2(n24662), .B1(n25200), .B2(n17478), .ZN(
        n21875) );
  OAI221_X1 U21369 ( .B1(n21364), .B2(n25218), .C1(n20284), .C2(n25212), .A(
        n21857), .ZN(n21852) );
  AOI22_X1 U21370 ( .A1(n25206), .A2(n24663), .B1(n25200), .B2(n17457), .ZN(
        n21857) );
  OAI221_X1 U21371 ( .B1(n21363), .B2(n25218), .C1(n20283), .C2(n25212), .A(
        n21839), .ZN(n21834) );
  AOI22_X1 U21372 ( .A1(n25206), .A2(n24664), .B1(n25200), .B2(n17436), .ZN(
        n21839) );
  OAI221_X1 U21373 ( .B1(n21362), .B2(n25218), .C1(n20282), .C2(n25212), .A(
        n21821), .ZN(n21816) );
  AOI22_X1 U21374 ( .A1(n25206), .A2(n24665), .B1(n25200), .B2(n17415), .ZN(
        n21821) );
  OAI221_X1 U21375 ( .B1(n21361), .B2(n25218), .C1(n20281), .C2(n25212), .A(
        n21803), .ZN(n21798) );
  AOI22_X1 U21376 ( .A1(n25206), .A2(n24666), .B1(n25200), .B2(n17394), .ZN(
        n21803) );
  OAI221_X1 U21377 ( .B1(n21360), .B2(n25218), .C1(n20280), .C2(n25212), .A(
        n21785), .ZN(n21780) );
  AOI22_X1 U21378 ( .A1(n25206), .A2(n24667), .B1(n25200), .B2(n17373), .ZN(
        n21785) );
  OAI221_X1 U21379 ( .B1(n21359), .B2(n25218), .C1(n20279), .C2(n25212), .A(
        n21767), .ZN(n21762) );
  AOI22_X1 U21380 ( .A1(n25206), .A2(n24668), .B1(n25200), .B2(n17352), .ZN(
        n21767) );
  OAI221_X1 U21381 ( .B1(n21358), .B2(n25218), .C1(n20278), .C2(n25212), .A(
        n21749), .ZN(n21744) );
  AOI22_X1 U21382 ( .A1(n25206), .A2(n24669), .B1(n25200), .B2(n17331), .ZN(
        n21749) );
  OAI221_X1 U21383 ( .B1(n21357), .B2(n25218), .C1(n20277), .C2(n25212), .A(
        n21731), .ZN(n21726) );
  AOI22_X1 U21384 ( .A1(n25206), .A2(n24670), .B1(n25200), .B2(n17310), .ZN(
        n21731) );
  OAI221_X1 U21385 ( .B1(n21356), .B2(n25218), .C1(n20276), .C2(n25212), .A(
        n21713), .ZN(n21708) );
  AOI22_X1 U21386 ( .A1(n25206), .A2(n24671), .B1(n25200), .B2(n17289), .ZN(
        n21713) );
  OAI221_X1 U21387 ( .B1(n21355), .B2(n25218), .C1(n20275), .C2(n25212), .A(
        n21695), .ZN(n21690) );
  AOI22_X1 U21388 ( .A1(n25206), .A2(n24672), .B1(n25200), .B2(n17268), .ZN(
        n21695) );
  OAI221_X1 U21389 ( .B1(n21354), .B2(n25218), .C1(n20274), .C2(n25212), .A(
        n21677), .ZN(n21672) );
  AOI22_X1 U21390 ( .A1(n25206), .A2(n24673), .B1(n25200), .B2(n17247), .ZN(
        n21677) );
  OAI221_X1 U21391 ( .B1(n21222), .B2(n25123), .C1(n19558), .C2(n25117), .A(
        n22771), .ZN(n22756) );
  AOI22_X1 U21392 ( .A1(n25111), .A2(n24481), .B1(n25105), .B2(n20005), .ZN(
        n22771) );
  OAI221_X1 U21393 ( .B1(n21350), .B2(n25021), .C1(n20270), .C2(n25015), .A(
        n22796), .ZN(n22781) );
  AOI22_X1 U21394 ( .A1(n25009), .A2(n24613), .B1(n25003), .B2(n17163), .ZN(
        n22796) );
  OAI221_X1 U21395 ( .B1(n21225), .B2(n25123), .C1(n19561), .C2(n25117), .A(
        n22848), .ZN(n22843) );
  AOI22_X1 U21396 ( .A1(n25111), .A2(n24478), .B1(n25105), .B2(n20008), .ZN(
        n22848) );
  OAI221_X1 U21397 ( .B1(n21353), .B2(n25021), .C1(n20273), .C2(n25015), .A(
        n22856), .ZN(n22851) );
  AOI22_X1 U21398 ( .A1(n25009), .A2(n24607), .B1(n25003), .B2(n17226), .ZN(
        n22856) );
  OAI221_X1 U21399 ( .B1(n21224), .B2(n25123), .C1(n19560), .C2(n25117), .A(
        n22830), .ZN(n22825) );
  AOI22_X1 U21400 ( .A1(n25111), .A2(n24479), .B1(n25105), .B2(n20007), .ZN(
        n22830) );
  OAI221_X1 U21401 ( .B1(n21352), .B2(n25021), .C1(n20272), .C2(n25015), .A(
        n22838), .ZN(n22833) );
  AOI22_X1 U21402 ( .A1(n25009), .A2(n24609), .B1(n25003), .B2(n17205), .ZN(
        n22838) );
  OAI221_X1 U21403 ( .B1(n21223), .B2(n25123), .C1(n19559), .C2(n25117), .A(
        n22812), .ZN(n22807) );
  AOI22_X1 U21404 ( .A1(n25111), .A2(n24480), .B1(n25105), .B2(n20006), .ZN(
        n22812) );
  OAI221_X1 U21405 ( .B1(n21351), .B2(n25021), .C1(n20271), .C2(n25015), .A(
        n22820), .ZN(n22815) );
  AOI22_X1 U21406 ( .A1(n25009), .A2(n24611), .B1(n25003), .B2(n17184), .ZN(
        n22820) );
  OAI221_X1 U21407 ( .B1(n21225), .B2(n25321), .C1(n19561), .C2(n25315), .A(
        n21651), .ZN(n21646) );
  AOI22_X1 U21408 ( .A1(n25309), .A2(n24478), .B1(n25303), .B2(n20008), .ZN(
        n21651) );
  OAI221_X1 U21409 ( .B1(n21353), .B2(n25219), .C1(n20273), .C2(n25213), .A(
        n21659), .ZN(n21654) );
  AOI22_X1 U21410 ( .A1(n25207), .A2(n24607), .B1(n25201), .B2(n17226), .ZN(
        n21659) );
  OAI221_X1 U21411 ( .B1(n21224), .B2(n25321), .C1(n19560), .C2(n25315), .A(
        n21633), .ZN(n21628) );
  AOI22_X1 U21412 ( .A1(n25309), .A2(n24479), .B1(n25303), .B2(n20007), .ZN(
        n21633) );
  OAI221_X1 U21413 ( .B1(n21352), .B2(n25219), .C1(n20272), .C2(n25213), .A(
        n21641), .ZN(n21636) );
  AOI22_X1 U21414 ( .A1(n25207), .A2(n24609), .B1(n25201), .B2(n17205), .ZN(
        n21641) );
  OAI221_X1 U21415 ( .B1(n21223), .B2(n25321), .C1(n19559), .C2(n25315), .A(
        n21615), .ZN(n21610) );
  AOI22_X1 U21416 ( .A1(n25309), .A2(n24480), .B1(n25303), .B2(n20006), .ZN(
        n21615) );
  OAI221_X1 U21417 ( .B1(n21351), .B2(n25219), .C1(n20271), .C2(n25213), .A(
        n21623), .ZN(n21618) );
  AOI22_X1 U21418 ( .A1(n25207), .A2(n24611), .B1(n25201), .B2(n17184), .ZN(
        n21623) );
  OAI221_X1 U21419 ( .B1(n21222), .B2(n25321), .C1(n19558), .C2(n25315), .A(
        n21574), .ZN(n21559) );
  AOI22_X1 U21420 ( .A1(n25309), .A2(n24481), .B1(n25303), .B2(n20005), .ZN(
        n21574) );
  OAI221_X1 U21421 ( .B1(n21350), .B2(n25219), .C1(n20270), .C2(n25213), .A(
        n21599), .ZN(n21584) );
  AOI22_X1 U21422 ( .A1(n25207), .A2(n24613), .B1(n25201), .B2(n17163), .ZN(
        n21599) );
  OAI221_X1 U21423 ( .B1(n20697), .B2(n25095), .C1(n21017), .C2(n25089), .A(
        n23713), .ZN(n23706) );
  AOI222_X1 U21424 ( .A1(n25083), .A2(n24206), .B1(n25077), .B2(n18228), .C1(
        n25071), .C2(n18227), .ZN(n23713) );
  OAI221_X1 U21425 ( .B1(n20696), .B2(n25095), .C1(n21016), .C2(n25089), .A(
        n23695), .ZN(n23688) );
  AOI222_X1 U21426 ( .A1(n25083), .A2(n24208), .B1(n25077), .B2(n18207), .C1(
        n25071), .C2(n18206), .ZN(n23695) );
  OAI221_X1 U21427 ( .B1(n20695), .B2(n25095), .C1(n21015), .C2(n25089), .A(
        n23677), .ZN(n23670) );
  AOI222_X1 U21428 ( .A1(n25083), .A2(n24210), .B1(n25077), .B2(n18186), .C1(
        n25071), .C2(n18185), .ZN(n23677) );
  OAI221_X1 U21429 ( .B1(n20694), .B2(n25095), .C1(n21014), .C2(n25089), .A(
        n23659), .ZN(n23652) );
  AOI222_X1 U21430 ( .A1(n25083), .A2(n24212), .B1(n25077), .B2(n18165), .C1(
        n25071), .C2(n18164), .ZN(n23659) );
  OAI221_X1 U21431 ( .B1(n20693), .B2(n25095), .C1(n21013), .C2(n25089), .A(
        n23641), .ZN(n23634) );
  AOI222_X1 U21432 ( .A1(n25083), .A2(n24214), .B1(n25077), .B2(n18144), .C1(
        n25071), .C2(n18143), .ZN(n23641) );
  OAI221_X1 U21433 ( .B1(n20692), .B2(n25095), .C1(n21012), .C2(n25089), .A(
        n23623), .ZN(n23616) );
  AOI222_X1 U21434 ( .A1(n25083), .A2(n24216), .B1(n25077), .B2(n18123), .C1(
        n25071), .C2(n18122), .ZN(n23623) );
  OAI221_X1 U21435 ( .B1(n20691), .B2(n25095), .C1(n21011), .C2(n25089), .A(
        n23605), .ZN(n23598) );
  AOI222_X1 U21436 ( .A1(n25083), .A2(n24218), .B1(n25077), .B2(n18102), .C1(
        n25071), .C2(n18101), .ZN(n23605) );
  OAI221_X1 U21437 ( .B1(n20690), .B2(n25095), .C1(n21010), .C2(n25089), .A(
        n23587), .ZN(n23580) );
  AOI222_X1 U21438 ( .A1(n25083), .A2(n24220), .B1(n25077), .B2(n18081), .C1(
        n25071), .C2(n18080), .ZN(n23587) );
  OAI221_X1 U21439 ( .B1(n20689), .B2(n25095), .C1(n21009), .C2(n25089), .A(
        n23569), .ZN(n23562) );
  AOI222_X1 U21440 ( .A1(n25083), .A2(n24222), .B1(n25077), .B2(n18060), .C1(
        n25071), .C2(n18059), .ZN(n23569) );
  OAI221_X1 U21441 ( .B1(n20688), .B2(n25095), .C1(n21008), .C2(n25089), .A(
        n23551), .ZN(n23544) );
  AOI222_X1 U21442 ( .A1(n25083), .A2(n24224), .B1(n25077), .B2(n18039), .C1(
        n25071), .C2(n18038), .ZN(n23551) );
  OAI221_X1 U21443 ( .B1(n20687), .B2(n25095), .C1(n21007), .C2(n25089), .A(
        n23533), .ZN(n23526) );
  AOI222_X1 U21444 ( .A1(n25083), .A2(n24226), .B1(n25077), .B2(n18018), .C1(
        n25071), .C2(n18017), .ZN(n23533) );
  OAI221_X1 U21445 ( .B1(n20686), .B2(n25095), .C1(n21006), .C2(n25089), .A(
        n23515), .ZN(n23508) );
  AOI222_X1 U21446 ( .A1(n25083), .A2(n24228), .B1(n25077), .B2(n17997), .C1(
        n25071), .C2(n17996), .ZN(n23515) );
  OAI221_X1 U21447 ( .B1(n20685), .B2(n25096), .C1(n21005), .C2(n25090), .A(
        n23497), .ZN(n23490) );
  AOI222_X1 U21448 ( .A1(n25084), .A2(n24230), .B1(n25078), .B2(n17976), .C1(
        n25072), .C2(n17975), .ZN(n23497) );
  OAI221_X1 U21449 ( .B1(n20684), .B2(n25096), .C1(n21004), .C2(n25090), .A(
        n23479), .ZN(n23472) );
  AOI222_X1 U21450 ( .A1(n25084), .A2(n24232), .B1(n25078), .B2(n17955), .C1(
        n25072), .C2(n17954), .ZN(n23479) );
  OAI221_X1 U21451 ( .B1(n20683), .B2(n25096), .C1(n21003), .C2(n25090), .A(
        n23461), .ZN(n23454) );
  AOI222_X1 U21452 ( .A1(n25084), .A2(n24234), .B1(n25078), .B2(n17934), .C1(
        n25072), .C2(n17933), .ZN(n23461) );
  OAI221_X1 U21453 ( .B1(n20682), .B2(n25096), .C1(n21002), .C2(n25090), .A(
        n23443), .ZN(n23436) );
  AOI222_X1 U21454 ( .A1(n25084), .A2(n24236), .B1(n25078), .B2(n17913), .C1(
        n25072), .C2(n17912), .ZN(n23443) );
  OAI221_X1 U21455 ( .B1(n20681), .B2(n25096), .C1(n21001), .C2(n25090), .A(
        n23425), .ZN(n23418) );
  AOI222_X1 U21456 ( .A1(n25084), .A2(n24238), .B1(n25078), .B2(n17892), .C1(
        n25072), .C2(n17891), .ZN(n23425) );
  OAI221_X1 U21457 ( .B1(n20680), .B2(n25096), .C1(n21000), .C2(n25090), .A(
        n23407), .ZN(n23400) );
  AOI222_X1 U21458 ( .A1(n25084), .A2(n24240), .B1(n25078), .B2(n17871), .C1(
        n25072), .C2(n17870), .ZN(n23407) );
  OAI221_X1 U21459 ( .B1(n20679), .B2(n25096), .C1(n20999), .C2(n25090), .A(
        n23389), .ZN(n23382) );
  AOI222_X1 U21460 ( .A1(n25084), .A2(n24242), .B1(n25078), .B2(n17850), .C1(
        n25072), .C2(n17849), .ZN(n23389) );
  OAI221_X1 U21461 ( .B1(n20678), .B2(n25096), .C1(n20998), .C2(n25090), .A(
        n23371), .ZN(n23364) );
  AOI222_X1 U21462 ( .A1(n25084), .A2(n24244), .B1(n25078), .B2(n17829), .C1(
        n25072), .C2(n17828), .ZN(n23371) );
  OAI221_X1 U21463 ( .B1(n20677), .B2(n25096), .C1(n20997), .C2(n25090), .A(
        n23353), .ZN(n23346) );
  AOI222_X1 U21464 ( .A1(n25084), .A2(n24246), .B1(n25078), .B2(n17808), .C1(
        n25072), .C2(n17807), .ZN(n23353) );
  OAI221_X1 U21465 ( .B1(n20676), .B2(n25096), .C1(n20996), .C2(n25090), .A(
        n23335), .ZN(n23328) );
  AOI222_X1 U21466 ( .A1(n25084), .A2(n24248), .B1(n25078), .B2(n17787), .C1(
        n25072), .C2(n17786), .ZN(n23335) );
  OAI221_X1 U21467 ( .B1(n20675), .B2(n25096), .C1(n20995), .C2(n25090), .A(
        n23317), .ZN(n23310) );
  AOI222_X1 U21468 ( .A1(n25084), .A2(n24250), .B1(n25078), .B2(n17766), .C1(
        n25072), .C2(n17765), .ZN(n23317) );
  OAI221_X1 U21469 ( .B1(n20674), .B2(n25096), .C1(n20994), .C2(n25090), .A(
        n23299), .ZN(n23292) );
  AOI222_X1 U21470 ( .A1(n25084), .A2(n24252), .B1(n25078), .B2(n17745), .C1(
        n25072), .C2(n17744), .ZN(n23299) );
  OAI221_X1 U21471 ( .B1(n20673), .B2(n25097), .C1(n20993), .C2(n25091), .A(
        n23281), .ZN(n23274) );
  AOI222_X1 U21472 ( .A1(n25085), .A2(n24254), .B1(n25079), .B2(n17724), .C1(
        n25073), .C2(n17723), .ZN(n23281) );
  OAI221_X1 U21473 ( .B1(n20672), .B2(n25097), .C1(n20992), .C2(n25091), .A(
        n23263), .ZN(n23256) );
  AOI222_X1 U21474 ( .A1(n25085), .A2(n24256), .B1(n25079), .B2(n17703), .C1(
        n25073), .C2(n17702), .ZN(n23263) );
  OAI221_X1 U21475 ( .B1(n20671), .B2(n25097), .C1(n20991), .C2(n25091), .A(
        n23245), .ZN(n23238) );
  AOI222_X1 U21476 ( .A1(n25085), .A2(n24258), .B1(n25079), .B2(n17682), .C1(
        n25073), .C2(n17681), .ZN(n23245) );
  OAI221_X1 U21477 ( .B1(n20670), .B2(n25097), .C1(n20990), .C2(n25091), .A(
        n23227), .ZN(n23220) );
  AOI222_X1 U21478 ( .A1(n25085), .A2(n24260), .B1(n25079), .B2(n17661), .C1(
        n25073), .C2(n17660), .ZN(n23227) );
  OAI221_X1 U21479 ( .B1(n20669), .B2(n25097), .C1(n20989), .C2(n25091), .A(
        n23209), .ZN(n23202) );
  AOI222_X1 U21480 ( .A1(n25085), .A2(n24262), .B1(n25079), .B2(n17640), .C1(
        n25073), .C2(n17639), .ZN(n23209) );
  OAI221_X1 U21481 ( .B1(n20668), .B2(n25097), .C1(n20988), .C2(n25091), .A(
        n23191), .ZN(n23184) );
  AOI222_X1 U21482 ( .A1(n25085), .A2(n24264), .B1(n25079), .B2(n17619), .C1(
        n25073), .C2(n17618), .ZN(n23191) );
  OAI221_X1 U21483 ( .B1(n20667), .B2(n25097), .C1(n20987), .C2(n25091), .A(
        n23173), .ZN(n23166) );
  AOI222_X1 U21484 ( .A1(n25085), .A2(n24266), .B1(n25079), .B2(n17598), .C1(
        n25073), .C2(n17597), .ZN(n23173) );
  OAI221_X1 U21485 ( .B1(n20666), .B2(n25097), .C1(n20986), .C2(n25091), .A(
        n23155), .ZN(n23148) );
  AOI222_X1 U21486 ( .A1(n25085), .A2(n24268), .B1(n25079), .B2(n17577), .C1(
        n25073), .C2(n17576), .ZN(n23155) );
  OAI221_X1 U21487 ( .B1(n20665), .B2(n25097), .C1(n20985), .C2(n25091), .A(
        n23137), .ZN(n23130) );
  AOI222_X1 U21488 ( .A1(n25085), .A2(n24270), .B1(n25079), .B2(n17556), .C1(
        n25073), .C2(n17555), .ZN(n23137) );
  OAI221_X1 U21489 ( .B1(n20664), .B2(n25097), .C1(n20984), .C2(n25091), .A(
        n23119), .ZN(n23112) );
  AOI222_X1 U21490 ( .A1(n25085), .A2(n24272), .B1(n25079), .B2(n17535), .C1(
        n25073), .C2(n17534), .ZN(n23119) );
  OAI221_X1 U21491 ( .B1(n20663), .B2(n25097), .C1(n20983), .C2(n25091), .A(
        n23101), .ZN(n23094) );
  AOI222_X1 U21492 ( .A1(n25085), .A2(n24274), .B1(n25079), .B2(n17514), .C1(
        n25073), .C2(n17513), .ZN(n23101) );
  OAI221_X1 U21493 ( .B1(n20662), .B2(n25097), .C1(n20982), .C2(n25091), .A(
        n23083), .ZN(n23076) );
  AOI222_X1 U21494 ( .A1(n25085), .A2(n24276), .B1(n25079), .B2(n17493), .C1(
        n25073), .C2(n17492), .ZN(n23083) );
  OAI221_X1 U21495 ( .B1(n20661), .B2(n25098), .C1(n20981), .C2(n25092), .A(
        n23065), .ZN(n23058) );
  AOI222_X1 U21496 ( .A1(n25086), .A2(n24278), .B1(n25080), .B2(n17472), .C1(
        n25074), .C2(n17471), .ZN(n23065) );
  OAI221_X1 U21497 ( .B1(n20660), .B2(n25098), .C1(n20980), .C2(n25092), .A(
        n23047), .ZN(n23040) );
  AOI222_X1 U21498 ( .A1(n25086), .A2(n24280), .B1(n25080), .B2(n17451), .C1(
        n25074), .C2(n17450), .ZN(n23047) );
  OAI221_X1 U21499 ( .B1(n20659), .B2(n25098), .C1(n20979), .C2(n25092), .A(
        n23029), .ZN(n23022) );
  AOI222_X1 U21500 ( .A1(n25086), .A2(n24282), .B1(n25080), .B2(n17430), .C1(
        n25074), .C2(n17429), .ZN(n23029) );
  OAI221_X1 U21501 ( .B1(n20658), .B2(n25098), .C1(n20978), .C2(n25092), .A(
        n23011), .ZN(n23004) );
  AOI222_X1 U21502 ( .A1(n25086), .A2(n24284), .B1(n25080), .B2(n17409), .C1(
        n25074), .C2(n17408), .ZN(n23011) );
  OAI221_X1 U21503 ( .B1(n20657), .B2(n25098), .C1(n20977), .C2(n25092), .A(
        n22993), .ZN(n22986) );
  AOI222_X1 U21504 ( .A1(n25086), .A2(n24286), .B1(n25080), .B2(n17388), .C1(
        n25074), .C2(n17387), .ZN(n22993) );
  OAI221_X1 U21505 ( .B1(n20656), .B2(n25098), .C1(n20976), .C2(n25092), .A(
        n22975), .ZN(n22968) );
  AOI222_X1 U21506 ( .A1(n25086), .A2(n24288), .B1(n25080), .B2(n17367), .C1(
        n25074), .C2(n17366), .ZN(n22975) );
  OAI221_X1 U21507 ( .B1(n20655), .B2(n25098), .C1(n20975), .C2(n25092), .A(
        n22957), .ZN(n22950) );
  AOI222_X1 U21508 ( .A1(n25086), .A2(n24290), .B1(n25080), .B2(n17346), .C1(
        n25074), .C2(n17345), .ZN(n22957) );
  OAI221_X1 U21509 ( .B1(n20654), .B2(n25098), .C1(n20974), .C2(n25092), .A(
        n22939), .ZN(n22932) );
  AOI222_X1 U21510 ( .A1(n25086), .A2(n24292), .B1(n25080), .B2(n17325), .C1(
        n25074), .C2(n17324), .ZN(n22939) );
  OAI221_X1 U21511 ( .B1(n20653), .B2(n25098), .C1(n20973), .C2(n25092), .A(
        n22921), .ZN(n22914) );
  AOI222_X1 U21512 ( .A1(n25086), .A2(n24294), .B1(n25080), .B2(n17304), .C1(
        n25074), .C2(n17303), .ZN(n22921) );
  OAI221_X1 U21513 ( .B1(n20652), .B2(n25098), .C1(n20972), .C2(n25092), .A(
        n22903), .ZN(n22896) );
  AOI222_X1 U21514 ( .A1(n25086), .A2(n24296), .B1(n25080), .B2(n17283), .C1(
        n25074), .C2(n17282), .ZN(n22903) );
  OAI221_X1 U21515 ( .B1(n20651), .B2(n25098), .C1(n20971), .C2(n25092), .A(
        n22885), .ZN(n22878) );
  AOI222_X1 U21516 ( .A1(n25086), .A2(n24298), .B1(n25080), .B2(n17262), .C1(
        n25074), .C2(n17261), .ZN(n22885) );
  OAI221_X1 U21517 ( .B1(n20650), .B2(n25098), .C1(n20970), .C2(n25092), .A(
        n22867), .ZN(n22860) );
  AOI222_X1 U21518 ( .A1(n25086), .A2(n24300), .B1(n25080), .B2(n17241), .C1(
        n25074), .C2(n17240), .ZN(n22867) );
  OAI221_X1 U21519 ( .B1(n20697), .B2(n25293), .C1(n21017), .C2(n25287), .A(
        n22516), .ZN(n22509) );
  AOI222_X1 U21520 ( .A1(n25281), .A2(n24206), .B1(n25275), .B2(n18228), .C1(
        n25269), .C2(n18227), .ZN(n22516) );
  OAI221_X1 U21521 ( .B1(n20696), .B2(n25293), .C1(n21016), .C2(n25287), .A(
        n22498), .ZN(n22491) );
  AOI222_X1 U21522 ( .A1(n25281), .A2(n24208), .B1(n25275), .B2(n18207), .C1(
        n25269), .C2(n18206), .ZN(n22498) );
  OAI221_X1 U21523 ( .B1(n20695), .B2(n25293), .C1(n21015), .C2(n25287), .A(
        n22480), .ZN(n22473) );
  AOI222_X1 U21524 ( .A1(n25281), .A2(n24210), .B1(n25275), .B2(n18186), .C1(
        n25269), .C2(n18185), .ZN(n22480) );
  OAI221_X1 U21525 ( .B1(n20694), .B2(n25293), .C1(n21014), .C2(n25287), .A(
        n22462), .ZN(n22455) );
  AOI222_X1 U21526 ( .A1(n25281), .A2(n24212), .B1(n25275), .B2(n18165), .C1(
        n25269), .C2(n18164), .ZN(n22462) );
  OAI221_X1 U21527 ( .B1(n20693), .B2(n25293), .C1(n21013), .C2(n25287), .A(
        n22444), .ZN(n22437) );
  AOI222_X1 U21528 ( .A1(n25281), .A2(n24214), .B1(n25275), .B2(n18144), .C1(
        n25269), .C2(n18143), .ZN(n22444) );
  OAI221_X1 U21529 ( .B1(n20692), .B2(n25293), .C1(n21012), .C2(n25287), .A(
        n22426), .ZN(n22419) );
  AOI222_X1 U21530 ( .A1(n25281), .A2(n24216), .B1(n25275), .B2(n18123), .C1(
        n25269), .C2(n18122), .ZN(n22426) );
  OAI221_X1 U21531 ( .B1(n20691), .B2(n25293), .C1(n21011), .C2(n25287), .A(
        n22408), .ZN(n22401) );
  AOI222_X1 U21532 ( .A1(n25281), .A2(n24218), .B1(n25275), .B2(n18102), .C1(
        n25269), .C2(n18101), .ZN(n22408) );
  OAI221_X1 U21533 ( .B1(n20690), .B2(n25293), .C1(n21010), .C2(n25287), .A(
        n22390), .ZN(n22383) );
  AOI222_X1 U21534 ( .A1(n25281), .A2(n24220), .B1(n25275), .B2(n18081), .C1(
        n25269), .C2(n18080), .ZN(n22390) );
  OAI221_X1 U21535 ( .B1(n20689), .B2(n25293), .C1(n21009), .C2(n25287), .A(
        n22372), .ZN(n22365) );
  AOI222_X1 U21536 ( .A1(n25281), .A2(n24222), .B1(n25275), .B2(n18060), .C1(
        n25269), .C2(n18059), .ZN(n22372) );
  OAI221_X1 U21537 ( .B1(n20688), .B2(n25293), .C1(n21008), .C2(n25287), .A(
        n22354), .ZN(n22347) );
  AOI222_X1 U21538 ( .A1(n25281), .A2(n24224), .B1(n25275), .B2(n18039), .C1(
        n25269), .C2(n18038), .ZN(n22354) );
  OAI221_X1 U21539 ( .B1(n20687), .B2(n25293), .C1(n21007), .C2(n25287), .A(
        n22336), .ZN(n22329) );
  AOI222_X1 U21540 ( .A1(n25281), .A2(n24226), .B1(n25275), .B2(n18018), .C1(
        n25269), .C2(n18017), .ZN(n22336) );
  OAI221_X1 U21541 ( .B1(n20686), .B2(n25293), .C1(n21006), .C2(n25287), .A(
        n22318), .ZN(n22311) );
  AOI222_X1 U21542 ( .A1(n25281), .A2(n24228), .B1(n25275), .B2(n17997), .C1(
        n25269), .C2(n17996), .ZN(n22318) );
  OAI221_X1 U21543 ( .B1(n20685), .B2(n25294), .C1(n21005), .C2(n25288), .A(
        n22300), .ZN(n22293) );
  AOI222_X1 U21544 ( .A1(n25282), .A2(n24230), .B1(n25276), .B2(n17976), .C1(
        n25270), .C2(n17975), .ZN(n22300) );
  OAI221_X1 U21545 ( .B1(n20684), .B2(n25294), .C1(n21004), .C2(n25288), .A(
        n22282), .ZN(n22275) );
  AOI222_X1 U21546 ( .A1(n25282), .A2(n24232), .B1(n25276), .B2(n17955), .C1(
        n25270), .C2(n17954), .ZN(n22282) );
  OAI221_X1 U21547 ( .B1(n20683), .B2(n25294), .C1(n21003), .C2(n25288), .A(
        n22264), .ZN(n22257) );
  AOI222_X1 U21548 ( .A1(n25282), .A2(n24234), .B1(n25276), .B2(n17934), .C1(
        n25270), .C2(n17933), .ZN(n22264) );
  OAI221_X1 U21549 ( .B1(n20682), .B2(n25294), .C1(n21002), .C2(n25288), .A(
        n22246), .ZN(n22239) );
  AOI222_X1 U21550 ( .A1(n25282), .A2(n24236), .B1(n25276), .B2(n17913), .C1(
        n25270), .C2(n17912), .ZN(n22246) );
  OAI221_X1 U21551 ( .B1(n20681), .B2(n25294), .C1(n21001), .C2(n25288), .A(
        n22228), .ZN(n22221) );
  AOI222_X1 U21552 ( .A1(n25282), .A2(n24238), .B1(n25276), .B2(n17892), .C1(
        n25270), .C2(n17891), .ZN(n22228) );
  OAI221_X1 U21553 ( .B1(n20680), .B2(n25294), .C1(n21000), .C2(n25288), .A(
        n22210), .ZN(n22203) );
  AOI222_X1 U21554 ( .A1(n25282), .A2(n24240), .B1(n25276), .B2(n17871), .C1(
        n25270), .C2(n17870), .ZN(n22210) );
  OAI221_X1 U21555 ( .B1(n20679), .B2(n25294), .C1(n20999), .C2(n25288), .A(
        n22192), .ZN(n22185) );
  AOI222_X1 U21556 ( .A1(n25282), .A2(n24242), .B1(n25276), .B2(n17850), .C1(
        n25270), .C2(n17849), .ZN(n22192) );
  OAI221_X1 U21557 ( .B1(n20678), .B2(n25294), .C1(n20998), .C2(n25288), .A(
        n22174), .ZN(n22167) );
  AOI222_X1 U21558 ( .A1(n25282), .A2(n24244), .B1(n25276), .B2(n17829), .C1(
        n25270), .C2(n17828), .ZN(n22174) );
  OAI221_X1 U21559 ( .B1(n20677), .B2(n25294), .C1(n20997), .C2(n25288), .A(
        n22156), .ZN(n22149) );
  AOI222_X1 U21560 ( .A1(n25282), .A2(n24246), .B1(n25276), .B2(n17808), .C1(
        n25270), .C2(n17807), .ZN(n22156) );
  OAI221_X1 U21561 ( .B1(n20676), .B2(n25294), .C1(n20996), .C2(n25288), .A(
        n22138), .ZN(n22131) );
  AOI222_X1 U21562 ( .A1(n25282), .A2(n24248), .B1(n25276), .B2(n17787), .C1(
        n25270), .C2(n17786), .ZN(n22138) );
  OAI221_X1 U21563 ( .B1(n20675), .B2(n25294), .C1(n20995), .C2(n25288), .A(
        n22120), .ZN(n22113) );
  AOI222_X1 U21564 ( .A1(n25282), .A2(n24250), .B1(n25276), .B2(n17766), .C1(
        n25270), .C2(n17765), .ZN(n22120) );
  OAI221_X1 U21565 ( .B1(n20674), .B2(n25294), .C1(n20994), .C2(n25288), .A(
        n22102), .ZN(n22095) );
  AOI222_X1 U21566 ( .A1(n25282), .A2(n24252), .B1(n25276), .B2(n17745), .C1(
        n25270), .C2(n17744), .ZN(n22102) );
  OAI221_X1 U21567 ( .B1(n20673), .B2(n25295), .C1(n20993), .C2(n25289), .A(
        n22084), .ZN(n22077) );
  AOI222_X1 U21568 ( .A1(n25283), .A2(n24254), .B1(n25277), .B2(n17724), .C1(
        n25271), .C2(n17723), .ZN(n22084) );
  OAI221_X1 U21569 ( .B1(n20672), .B2(n25295), .C1(n20992), .C2(n25289), .A(
        n22066), .ZN(n22059) );
  AOI222_X1 U21570 ( .A1(n25283), .A2(n24256), .B1(n25277), .B2(n17703), .C1(
        n25271), .C2(n17702), .ZN(n22066) );
  OAI221_X1 U21571 ( .B1(n20671), .B2(n25295), .C1(n20991), .C2(n25289), .A(
        n22048), .ZN(n22041) );
  AOI222_X1 U21572 ( .A1(n25283), .A2(n24258), .B1(n25277), .B2(n17682), .C1(
        n25271), .C2(n17681), .ZN(n22048) );
  OAI221_X1 U21573 ( .B1(n20670), .B2(n25295), .C1(n20990), .C2(n25289), .A(
        n22030), .ZN(n22023) );
  AOI222_X1 U21574 ( .A1(n25283), .A2(n24260), .B1(n25277), .B2(n17661), .C1(
        n25271), .C2(n17660), .ZN(n22030) );
  OAI221_X1 U21575 ( .B1(n20669), .B2(n25295), .C1(n20989), .C2(n25289), .A(
        n22012), .ZN(n22005) );
  AOI222_X1 U21576 ( .A1(n25283), .A2(n24262), .B1(n25277), .B2(n17640), .C1(
        n25271), .C2(n17639), .ZN(n22012) );
  OAI221_X1 U21577 ( .B1(n20668), .B2(n25295), .C1(n20988), .C2(n25289), .A(
        n21994), .ZN(n21987) );
  AOI222_X1 U21578 ( .A1(n25283), .A2(n24264), .B1(n25277), .B2(n17619), .C1(
        n25271), .C2(n17618), .ZN(n21994) );
  OAI221_X1 U21579 ( .B1(n20667), .B2(n25295), .C1(n20987), .C2(n25289), .A(
        n21976), .ZN(n21969) );
  AOI222_X1 U21580 ( .A1(n25283), .A2(n24266), .B1(n25277), .B2(n17598), .C1(
        n25271), .C2(n17597), .ZN(n21976) );
  OAI221_X1 U21581 ( .B1(n20666), .B2(n25295), .C1(n20986), .C2(n25289), .A(
        n21958), .ZN(n21951) );
  AOI222_X1 U21582 ( .A1(n25283), .A2(n24268), .B1(n25277), .B2(n17577), .C1(
        n25271), .C2(n17576), .ZN(n21958) );
  OAI221_X1 U21583 ( .B1(n20665), .B2(n25295), .C1(n20985), .C2(n25289), .A(
        n21940), .ZN(n21933) );
  AOI222_X1 U21584 ( .A1(n25283), .A2(n24270), .B1(n25277), .B2(n17556), .C1(
        n25271), .C2(n17555), .ZN(n21940) );
  OAI221_X1 U21585 ( .B1(n20664), .B2(n25295), .C1(n20984), .C2(n25289), .A(
        n21922), .ZN(n21915) );
  AOI222_X1 U21586 ( .A1(n25283), .A2(n24272), .B1(n25277), .B2(n17535), .C1(
        n25271), .C2(n17534), .ZN(n21922) );
  OAI221_X1 U21587 ( .B1(n20663), .B2(n25295), .C1(n20983), .C2(n25289), .A(
        n21904), .ZN(n21897) );
  AOI222_X1 U21588 ( .A1(n25283), .A2(n24274), .B1(n25277), .B2(n17514), .C1(
        n25271), .C2(n17513), .ZN(n21904) );
  OAI221_X1 U21589 ( .B1(n20662), .B2(n25295), .C1(n20982), .C2(n25289), .A(
        n21886), .ZN(n21879) );
  AOI222_X1 U21590 ( .A1(n25283), .A2(n24276), .B1(n25277), .B2(n17493), .C1(
        n25271), .C2(n17492), .ZN(n21886) );
  OAI221_X1 U21591 ( .B1(n20661), .B2(n25296), .C1(n20981), .C2(n25290), .A(
        n21868), .ZN(n21861) );
  AOI222_X1 U21592 ( .A1(n25284), .A2(n24278), .B1(n25278), .B2(n17472), .C1(
        n25272), .C2(n17471), .ZN(n21868) );
  OAI221_X1 U21593 ( .B1(n20660), .B2(n25296), .C1(n20980), .C2(n25290), .A(
        n21850), .ZN(n21843) );
  AOI222_X1 U21594 ( .A1(n25284), .A2(n24280), .B1(n25278), .B2(n17451), .C1(
        n25272), .C2(n17450), .ZN(n21850) );
  OAI221_X1 U21595 ( .B1(n20659), .B2(n25296), .C1(n20979), .C2(n25290), .A(
        n21832), .ZN(n21825) );
  AOI222_X1 U21596 ( .A1(n25284), .A2(n24282), .B1(n25278), .B2(n17430), .C1(
        n25272), .C2(n17429), .ZN(n21832) );
  OAI221_X1 U21597 ( .B1(n20658), .B2(n25296), .C1(n20978), .C2(n25290), .A(
        n21814), .ZN(n21807) );
  AOI222_X1 U21598 ( .A1(n25284), .A2(n24284), .B1(n25278), .B2(n17409), .C1(
        n25272), .C2(n17408), .ZN(n21814) );
  OAI221_X1 U21599 ( .B1(n20657), .B2(n25296), .C1(n20977), .C2(n25290), .A(
        n21796), .ZN(n21789) );
  AOI222_X1 U21600 ( .A1(n25284), .A2(n24286), .B1(n25278), .B2(n17388), .C1(
        n25272), .C2(n17387), .ZN(n21796) );
  OAI221_X1 U21601 ( .B1(n20656), .B2(n25296), .C1(n20976), .C2(n25290), .A(
        n21778), .ZN(n21771) );
  AOI222_X1 U21602 ( .A1(n25284), .A2(n24288), .B1(n25278), .B2(n17367), .C1(
        n25272), .C2(n17366), .ZN(n21778) );
  OAI221_X1 U21603 ( .B1(n20655), .B2(n25296), .C1(n20975), .C2(n25290), .A(
        n21760), .ZN(n21753) );
  AOI222_X1 U21604 ( .A1(n25284), .A2(n24290), .B1(n25278), .B2(n17346), .C1(
        n25272), .C2(n17345), .ZN(n21760) );
  OAI221_X1 U21605 ( .B1(n20654), .B2(n25296), .C1(n20974), .C2(n25290), .A(
        n21742), .ZN(n21735) );
  AOI222_X1 U21606 ( .A1(n25284), .A2(n24292), .B1(n25278), .B2(n17325), .C1(
        n25272), .C2(n17324), .ZN(n21742) );
  OAI221_X1 U21607 ( .B1(n20653), .B2(n25296), .C1(n20973), .C2(n25290), .A(
        n21724), .ZN(n21717) );
  AOI222_X1 U21608 ( .A1(n25284), .A2(n24294), .B1(n25278), .B2(n17304), .C1(
        n25272), .C2(n17303), .ZN(n21724) );
  OAI221_X1 U21609 ( .B1(n20652), .B2(n25296), .C1(n20972), .C2(n25290), .A(
        n21706), .ZN(n21699) );
  AOI222_X1 U21610 ( .A1(n25284), .A2(n24296), .B1(n25278), .B2(n17283), .C1(
        n25272), .C2(n17282), .ZN(n21706) );
  OAI221_X1 U21611 ( .B1(n20651), .B2(n25296), .C1(n20971), .C2(n25290), .A(
        n21688), .ZN(n21681) );
  AOI222_X1 U21612 ( .A1(n25284), .A2(n24298), .B1(n25278), .B2(n17262), .C1(
        n25272), .C2(n17261), .ZN(n21688) );
  OAI221_X1 U21613 ( .B1(n20650), .B2(n25296), .C1(n20970), .C2(n25290), .A(
        n21670), .ZN(n21663) );
  AOI222_X1 U21614 ( .A1(n25284), .A2(n24300), .B1(n25278), .B2(n17241), .C1(
        n25272), .C2(n17240), .ZN(n21670) );
  OAI221_X1 U21615 ( .B1(n20646), .B2(n25099), .C1(n20966), .C2(n25093), .A(
        n22776), .ZN(n22755) );
  AOI222_X1 U21616 ( .A1(n25087), .A2(n24311), .B1(n25081), .B2(n17157), .C1(
        n25075), .C2(n17156), .ZN(n22776) );
  OAI221_X1 U21617 ( .B1(n20649), .B2(n25099), .C1(n20969), .C2(n25093), .A(
        n22849), .ZN(n22842) );
  AOI222_X1 U21618 ( .A1(n25087), .A2(n24302), .B1(n25081), .B2(n17220), .C1(
        n25075), .C2(n17219), .ZN(n22849) );
  OAI221_X1 U21619 ( .B1(n20648), .B2(n25099), .C1(n20968), .C2(n25093), .A(
        n22831), .ZN(n22824) );
  AOI222_X1 U21620 ( .A1(n25087), .A2(n24305), .B1(n25081), .B2(n17199), .C1(
        n25075), .C2(n17198), .ZN(n22831) );
  OAI221_X1 U21621 ( .B1(n20647), .B2(n25099), .C1(n20967), .C2(n25093), .A(
        n22813), .ZN(n22806) );
  AOI222_X1 U21622 ( .A1(n25087), .A2(n24308), .B1(n25081), .B2(n17178), .C1(
        n25075), .C2(n17177), .ZN(n22813) );
  OAI221_X1 U21623 ( .B1(n20649), .B2(n25297), .C1(n20969), .C2(n25291), .A(
        n21652), .ZN(n21645) );
  AOI222_X1 U21624 ( .A1(n25285), .A2(n24302), .B1(n25279), .B2(n17220), .C1(
        n25273), .C2(n17219), .ZN(n21652) );
  OAI221_X1 U21625 ( .B1(n20648), .B2(n25297), .C1(n20968), .C2(n25291), .A(
        n21634), .ZN(n21627) );
  AOI222_X1 U21626 ( .A1(n25285), .A2(n24305), .B1(n25279), .B2(n17199), .C1(
        n25273), .C2(n17198), .ZN(n21634) );
  OAI221_X1 U21627 ( .B1(n20647), .B2(n25297), .C1(n20967), .C2(n25291), .A(
        n21616), .ZN(n21609) );
  AOI222_X1 U21628 ( .A1(n25285), .A2(n24308), .B1(n25279), .B2(n17178), .C1(
        n25273), .C2(n17177), .ZN(n21616) );
  OAI221_X1 U21629 ( .B1(n20646), .B2(n25297), .C1(n20966), .C2(n25291), .A(
        n21579), .ZN(n21558) );
  AOI222_X1 U21630 ( .A1(n25285), .A2(n24311), .B1(n25279), .B2(n17157), .C1(
        n25273), .C2(n17156), .ZN(n21579) );
  OAI221_X1 U21631 ( .B1(n21413), .B2(n25016), .C1(n20333), .C2(n25010), .A(
        n23948), .ZN(n23942) );
  AOI22_X1 U21632 ( .A1(n25004), .A2(n24614), .B1(n24998), .B2(n18486), .ZN(
        n23948) );
  OAI221_X1 U21633 ( .B1(n21412), .B2(n25016), .C1(n20332), .C2(n25010), .A(
        n23918), .ZN(n23913) );
  AOI22_X1 U21634 ( .A1(n25004), .A2(n24615), .B1(n24998), .B2(n18465), .ZN(
        n23918) );
  OAI221_X1 U21635 ( .B1(n21411), .B2(n25016), .C1(n20331), .C2(n25010), .A(
        n23900), .ZN(n23895) );
  AOI22_X1 U21636 ( .A1(n25004), .A2(n24616), .B1(n24998), .B2(n18444), .ZN(
        n23900) );
  OAI221_X1 U21637 ( .B1(n21410), .B2(n25016), .C1(n20330), .C2(n25010), .A(
        n23882), .ZN(n23877) );
  AOI22_X1 U21638 ( .A1(n25004), .A2(n24617), .B1(n24998), .B2(n18423), .ZN(
        n23882) );
  OAI221_X1 U21639 ( .B1(n21409), .B2(n25016), .C1(n20329), .C2(n25010), .A(
        n23864), .ZN(n23859) );
  AOI22_X1 U21640 ( .A1(n25004), .A2(n24618), .B1(n24998), .B2(n18402), .ZN(
        n23864) );
  OAI221_X1 U21641 ( .B1(n21408), .B2(n25016), .C1(n20328), .C2(n25010), .A(
        n23846), .ZN(n23841) );
  AOI22_X1 U21642 ( .A1(n25004), .A2(n24619), .B1(n24998), .B2(n18381), .ZN(
        n23846) );
  OAI221_X1 U21643 ( .B1(n21407), .B2(n25016), .C1(n20327), .C2(n25010), .A(
        n23828), .ZN(n23823) );
  AOI22_X1 U21644 ( .A1(n25004), .A2(n24620), .B1(n24998), .B2(n18360), .ZN(
        n23828) );
  OAI221_X1 U21645 ( .B1(n21406), .B2(n25016), .C1(n20326), .C2(n25010), .A(
        n23810), .ZN(n23805) );
  AOI22_X1 U21646 ( .A1(n25004), .A2(n24621), .B1(n24998), .B2(n18339), .ZN(
        n23810) );
  OAI221_X1 U21647 ( .B1(n21405), .B2(n25016), .C1(n20325), .C2(n25010), .A(
        n23792), .ZN(n23787) );
  AOI22_X1 U21648 ( .A1(n25004), .A2(n24622), .B1(n24998), .B2(n18318), .ZN(
        n23792) );
  OAI221_X1 U21649 ( .B1(n21404), .B2(n25016), .C1(n20324), .C2(n25010), .A(
        n23774), .ZN(n23769) );
  AOI22_X1 U21650 ( .A1(n25004), .A2(n24623), .B1(n24998), .B2(n18297), .ZN(
        n23774) );
  OAI221_X1 U21651 ( .B1(n21403), .B2(n25016), .C1(n20323), .C2(n25010), .A(
        n23756), .ZN(n23751) );
  AOI22_X1 U21652 ( .A1(n25004), .A2(n24624), .B1(n24998), .B2(n18276), .ZN(
        n23756) );
  OAI221_X1 U21653 ( .B1(n21402), .B2(n25016), .C1(n20322), .C2(n25010), .A(
        n23738), .ZN(n23733) );
  AOI22_X1 U21654 ( .A1(n25004), .A2(n24625), .B1(n24998), .B2(n18255), .ZN(
        n23738) );
  OAI221_X1 U21655 ( .B1(n21413), .B2(n25214), .C1(n20333), .C2(n25208), .A(
        n22751), .ZN(n22745) );
  AOI22_X1 U21656 ( .A1(n25202), .A2(n24614), .B1(n25196), .B2(n18486), .ZN(
        n22751) );
  OAI221_X1 U21657 ( .B1(n21412), .B2(n25214), .C1(n20332), .C2(n25208), .A(
        n22721), .ZN(n22716) );
  AOI22_X1 U21658 ( .A1(n25202), .A2(n24615), .B1(n25196), .B2(n18465), .ZN(
        n22721) );
  OAI221_X1 U21659 ( .B1(n21411), .B2(n25214), .C1(n20331), .C2(n25208), .A(
        n22703), .ZN(n22698) );
  AOI22_X1 U21660 ( .A1(n25202), .A2(n24616), .B1(n25196), .B2(n18444), .ZN(
        n22703) );
  OAI221_X1 U21661 ( .B1(n21410), .B2(n25214), .C1(n20330), .C2(n25208), .A(
        n22685), .ZN(n22680) );
  AOI22_X1 U21662 ( .A1(n25202), .A2(n24617), .B1(n25196), .B2(n18423), .ZN(
        n22685) );
  OAI221_X1 U21663 ( .B1(n21409), .B2(n25214), .C1(n20329), .C2(n25208), .A(
        n22667), .ZN(n22662) );
  AOI22_X1 U21664 ( .A1(n25202), .A2(n24618), .B1(n25196), .B2(n18402), .ZN(
        n22667) );
  OAI221_X1 U21665 ( .B1(n21408), .B2(n25214), .C1(n20328), .C2(n25208), .A(
        n22649), .ZN(n22644) );
  AOI22_X1 U21666 ( .A1(n25202), .A2(n24619), .B1(n25196), .B2(n18381), .ZN(
        n22649) );
  OAI221_X1 U21667 ( .B1(n21407), .B2(n25214), .C1(n20327), .C2(n25208), .A(
        n22631), .ZN(n22626) );
  AOI22_X1 U21668 ( .A1(n25202), .A2(n24620), .B1(n25196), .B2(n18360), .ZN(
        n22631) );
  OAI221_X1 U21669 ( .B1(n21406), .B2(n25214), .C1(n20326), .C2(n25208), .A(
        n22613), .ZN(n22608) );
  AOI22_X1 U21670 ( .A1(n25202), .A2(n24621), .B1(n25196), .B2(n18339), .ZN(
        n22613) );
  OAI221_X1 U21671 ( .B1(n21405), .B2(n25214), .C1(n20325), .C2(n25208), .A(
        n22595), .ZN(n22590) );
  AOI22_X1 U21672 ( .A1(n25202), .A2(n24622), .B1(n25196), .B2(n18318), .ZN(
        n22595) );
  OAI221_X1 U21673 ( .B1(n21404), .B2(n25214), .C1(n20324), .C2(n25208), .A(
        n22577), .ZN(n22572) );
  AOI22_X1 U21674 ( .A1(n25202), .A2(n24623), .B1(n25196), .B2(n18297), .ZN(
        n22577) );
  OAI221_X1 U21675 ( .B1(n21403), .B2(n25214), .C1(n20323), .C2(n25208), .A(
        n22559), .ZN(n22554) );
  AOI22_X1 U21676 ( .A1(n25202), .A2(n24624), .B1(n25196), .B2(n18276), .ZN(
        n22559) );
  OAI221_X1 U21677 ( .B1(n21402), .B2(n25214), .C1(n20322), .C2(n25208), .A(
        n22541), .ZN(n22536) );
  AOI22_X1 U21678 ( .A1(n25202), .A2(n24625), .B1(n25196), .B2(n18255), .ZN(
        n22541) );
  OAI221_X1 U21679 ( .B1(n20709), .B2(n25094), .C1(n21029), .C2(n25088), .A(
        n23938), .ZN(n23922) );
  AOI222_X1 U21680 ( .A1(n25082), .A2(n24314), .B1(n25076), .B2(n18480), .C1(
        n25070), .C2(n18479), .ZN(n23938) );
  OAI221_X1 U21681 ( .B1(n20708), .B2(n25094), .C1(n21028), .C2(n25088), .A(
        n23911), .ZN(n23904) );
  AOI222_X1 U21682 ( .A1(n25082), .A2(n24316), .B1(n25076), .B2(n18459), .C1(
        n25070), .C2(n18458), .ZN(n23911) );
  OAI221_X1 U21683 ( .B1(n20707), .B2(n25094), .C1(n21027), .C2(n25088), .A(
        n23893), .ZN(n23886) );
  AOI222_X1 U21684 ( .A1(n25082), .A2(n24318), .B1(n25076), .B2(n18438), .C1(
        n25070), .C2(n18437), .ZN(n23893) );
  OAI221_X1 U21685 ( .B1(n20706), .B2(n25094), .C1(n21026), .C2(n25088), .A(
        n23875), .ZN(n23868) );
  AOI222_X1 U21686 ( .A1(n25082), .A2(n24320), .B1(n25076), .B2(n18417), .C1(
        n25070), .C2(n18416), .ZN(n23875) );
  OAI221_X1 U21687 ( .B1(n20705), .B2(n25094), .C1(n21025), .C2(n25088), .A(
        n23857), .ZN(n23850) );
  AOI222_X1 U21688 ( .A1(n25082), .A2(n24322), .B1(n25076), .B2(n18396), .C1(
        n25070), .C2(n18395), .ZN(n23857) );
  OAI221_X1 U21689 ( .B1(n20704), .B2(n25094), .C1(n21024), .C2(n25088), .A(
        n23839), .ZN(n23832) );
  AOI222_X1 U21690 ( .A1(n25082), .A2(n24324), .B1(n25076), .B2(n18375), .C1(
        n25070), .C2(n18374), .ZN(n23839) );
  OAI221_X1 U21691 ( .B1(n20703), .B2(n25094), .C1(n21023), .C2(n25088), .A(
        n23821), .ZN(n23814) );
  AOI222_X1 U21692 ( .A1(n25082), .A2(n24326), .B1(n25076), .B2(n18354), .C1(
        n25070), .C2(n18353), .ZN(n23821) );
  OAI221_X1 U21693 ( .B1(n20702), .B2(n25094), .C1(n21022), .C2(n25088), .A(
        n23803), .ZN(n23796) );
  AOI222_X1 U21694 ( .A1(n25082), .A2(n24328), .B1(n25076), .B2(n18333), .C1(
        n25070), .C2(n18332), .ZN(n23803) );
  OAI221_X1 U21695 ( .B1(n20701), .B2(n25094), .C1(n21021), .C2(n25088), .A(
        n23785), .ZN(n23778) );
  AOI222_X1 U21696 ( .A1(n25082), .A2(n24330), .B1(n25076), .B2(n18312), .C1(
        n25070), .C2(n18311), .ZN(n23785) );
  OAI221_X1 U21697 ( .B1(n20700), .B2(n25094), .C1(n21020), .C2(n25088), .A(
        n23767), .ZN(n23760) );
  AOI222_X1 U21698 ( .A1(n25082), .A2(n24332), .B1(n25076), .B2(n18291), .C1(
        n25070), .C2(n18290), .ZN(n23767) );
  OAI221_X1 U21699 ( .B1(n20699), .B2(n25094), .C1(n21019), .C2(n25088), .A(
        n23749), .ZN(n23742) );
  AOI222_X1 U21700 ( .A1(n25082), .A2(n24334), .B1(n25076), .B2(n18270), .C1(
        n25070), .C2(n18269), .ZN(n23749) );
  OAI221_X1 U21701 ( .B1(n20698), .B2(n25094), .C1(n21018), .C2(n25088), .A(
        n23731), .ZN(n23724) );
  AOI222_X1 U21702 ( .A1(n25082), .A2(n24336), .B1(n25076), .B2(n18249), .C1(
        n25070), .C2(n18248), .ZN(n23731) );
  OAI221_X1 U21703 ( .B1(n20709), .B2(n25292), .C1(n21029), .C2(n25286), .A(
        n22741), .ZN(n22725) );
  AOI222_X1 U21704 ( .A1(n25280), .A2(n24314), .B1(n25274), .B2(n18480), .C1(
        n25268), .C2(n18479), .ZN(n22741) );
  OAI221_X1 U21705 ( .B1(n20708), .B2(n25292), .C1(n21028), .C2(n25286), .A(
        n22714), .ZN(n22707) );
  AOI222_X1 U21706 ( .A1(n25280), .A2(n24316), .B1(n25274), .B2(n18459), .C1(
        n25268), .C2(n18458), .ZN(n22714) );
  OAI221_X1 U21707 ( .B1(n20707), .B2(n25292), .C1(n21027), .C2(n25286), .A(
        n22696), .ZN(n22689) );
  AOI222_X1 U21708 ( .A1(n25280), .A2(n24318), .B1(n25274), .B2(n18438), .C1(
        n25268), .C2(n18437), .ZN(n22696) );
  OAI221_X1 U21709 ( .B1(n20706), .B2(n25292), .C1(n21026), .C2(n25286), .A(
        n22678), .ZN(n22671) );
  AOI222_X1 U21710 ( .A1(n25280), .A2(n24320), .B1(n25274), .B2(n18417), .C1(
        n25268), .C2(n18416), .ZN(n22678) );
  OAI221_X1 U21711 ( .B1(n20705), .B2(n25292), .C1(n21025), .C2(n25286), .A(
        n22660), .ZN(n22653) );
  AOI222_X1 U21712 ( .A1(n25280), .A2(n24322), .B1(n25274), .B2(n18396), .C1(
        n25268), .C2(n18395), .ZN(n22660) );
  OAI221_X1 U21713 ( .B1(n20704), .B2(n25292), .C1(n21024), .C2(n25286), .A(
        n22642), .ZN(n22635) );
  AOI222_X1 U21714 ( .A1(n25280), .A2(n24324), .B1(n25274), .B2(n18375), .C1(
        n25268), .C2(n18374), .ZN(n22642) );
  OAI221_X1 U21715 ( .B1(n20703), .B2(n25292), .C1(n21023), .C2(n25286), .A(
        n22624), .ZN(n22617) );
  AOI222_X1 U21716 ( .A1(n25280), .A2(n24326), .B1(n25274), .B2(n18354), .C1(
        n25268), .C2(n18353), .ZN(n22624) );
  OAI221_X1 U21717 ( .B1(n20702), .B2(n25292), .C1(n21022), .C2(n25286), .A(
        n22606), .ZN(n22599) );
  AOI222_X1 U21718 ( .A1(n25280), .A2(n24328), .B1(n25274), .B2(n18333), .C1(
        n25268), .C2(n18332), .ZN(n22606) );
  OAI221_X1 U21719 ( .B1(n20701), .B2(n25292), .C1(n21021), .C2(n25286), .A(
        n22588), .ZN(n22581) );
  AOI222_X1 U21720 ( .A1(n25280), .A2(n24330), .B1(n25274), .B2(n18312), .C1(
        n25268), .C2(n18311), .ZN(n22588) );
  OAI221_X1 U21721 ( .B1(n20700), .B2(n25292), .C1(n21020), .C2(n25286), .A(
        n22570), .ZN(n22563) );
  AOI222_X1 U21722 ( .A1(n25280), .A2(n24332), .B1(n25274), .B2(n18291), .C1(
        n25268), .C2(n18290), .ZN(n22570) );
  OAI221_X1 U21723 ( .B1(n20699), .B2(n25292), .C1(n21019), .C2(n25286), .A(
        n22552), .ZN(n22545) );
  AOI222_X1 U21724 ( .A1(n25280), .A2(n24334), .B1(n25274), .B2(n18270), .C1(
        n25268), .C2(n18269), .ZN(n22552) );
  OAI221_X1 U21725 ( .B1(n20698), .B2(n25292), .C1(n21018), .C2(n25286), .A(
        n22534), .ZN(n22527) );
  AOI222_X1 U21726 ( .A1(n25280), .A2(n24336), .B1(n25274), .B2(n18249), .C1(
        n25268), .C2(n18248), .ZN(n22534) );
  OAI22_X1 U21727 ( .A1(n9466), .A2(n25776), .B1(n25770), .B2(n25817), .ZN(
        n7435) );
  OAI22_X1 U21728 ( .A1(n9465), .A2(n25776), .B1(n25770), .B2(n25820), .ZN(
        n7436) );
  OAI22_X1 U21729 ( .A1(n9464), .A2(n25776), .B1(n25770), .B2(n25823), .ZN(
        n7437) );
  OAI22_X1 U21730 ( .A1(n9463), .A2(n25776), .B1(n25770), .B2(n25826), .ZN(
        n7438) );
  OAI22_X1 U21731 ( .A1(n9462), .A2(n25776), .B1(n25770), .B2(n25829), .ZN(
        n7439) );
  OAI22_X1 U21732 ( .A1(n9461), .A2(n25776), .B1(n25770), .B2(n25832), .ZN(
        n7440) );
  OAI22_X1 U21733 ( .A1(n9460), .A2(n25776), .B1(n25770), .B2(n25835), .ZN(
        n7441) );
  OAI22_X1 U21734 ( .A1(n9459), .A2(n25776), .B1(n25770), .B2(n25838), .ZN(
        n7442) );
  OAI22_X1 U21735 ( .A1(n9458), .A2(n25776), .B1(n25770), .B2(n25841), .ZN(
        n7443) );
  OAI22_X1 U21736 ( .A1(n9457), .A2(n25776), .B1(n25770), .B2(n25844), .ZN(
        n7444) );
  OAI22_X1 U21737 ( .A1(n9456), .A2(n25776), .B1(n25770), .B2(n25847), .ZN(
        n7445) );
  OAI22_X1 U21738 ( .A1(n9455), .A2(n25777), .B1(n25770), .B2(n25850), .ZN(
        n7446) );
  OAI22_X1 U21739 ( .A1(n9454), .A2(n25777), .B1(n25771), .B2(n25853), .ZN(
        n7447) );
  OAI22_X1 U21740 ( .A1(n9453), .A2(n25777), .B1(n25771), .B2(n25856), .ZN(
        n7448) );
  OAI22_X1 U21741 ( .A1(n9452), .A2(n25777), .B1(n25771), .B2(n25859), .ZN(
        n7449) );
  OAI22_X1 U21742 ( .A1(n9451), .A2(n25777), .B1(n25771), .B2(n25862), .ZN(
        n7450) );
  OAI22_X1 U21743 ( .A1(n9450), .A2(n25777), .B1(n25771), .B2(n25865), .ZN(
        n7451) );
  OAI22_X1 U21744 ( .A1(n9449), .A2(n25777), .B1(n25771), .B2(n25868), .ZN(
        n7452) );
  OAI22_X1 U21745 ( .A1(n9448), .A2(n25777), .B1(n25771), .B2(n25871), .ZN(
        n7453) );
  OAI22_X1 U21746 ( .A1(n9447), .A2(n25777), .B1(n25771), .B2(n25874), .ZN(
        n7454) );
  OAI22_X1 U21747 ( .A1(n9446), .A2(n25777), .B1(n25771), .B2(n25877), .ZN(
        n7455) );
  OAI22_X1 U21748 ( .A1(n9445), .A2(n25777), .B1(n25771), .B2(n25880), .ZN(
        n7456) );
  OAI22_X1 U21749 ( .A1(n9444), .A2(n25777), .B1(n25771), .B2(n25883), .ZN(
        n7457) );
  OAI22_X1 U21750 ( .A1(n9443), .A2(n25778), .B1(n25771), .B2(n25886), .ZN(
        n7458) );
  OAI22_X1 U21751 ( .A1(n9442), .A2(n25778), .B1(n25772), .B2(n25889), .ZN(
        n7459) );
  OAI22_X1 U21752 ( .A1(n9441), .A2(n25778), .B1(n25772), .B2(n25892), .ZN(
        n7460) );
  OAI22_X1 U21753 ( .A1(n9440), .A2(n25778), .B1(n25772), .B2(n25895), .ZN(
        n7461) );
  OAI22_X1 U21754 ( .A1(n9439), .A2(n25778), .B1(n25772), .B2(n25898), .ZN(
        n7462) );
  OAI22_X1 U21755 ( .A1(n9438), .A2(n25778), .B1(n25772), .B2(n25901), .ZN(
        n7463) );
  OAI22_X1 U21756 ( .A1(n9437), .A2(n25778), .B1(n25772), .B2(n25904), .ZN(
        n7464) );
  OAI22_X1 U21757 ( .A1(n9436), .A2(n25778), .B1(n25772), .B2(n25907), .ZN(
        n7465) );
  OAI22_X1 U21758 ( .A1(n9435), .A2(n25778), .B1(n25772), .B2(n25910), .ZN(
        n7466) );
  OAI22_X1 U21759 ( .A1(n9434), .A2(n25778), .B1(n25772), .B2(n25913), .ZN(
        n7467) );
  OAI22_X1 U21760 ( .A1(n9433), .A2(n25778), .B1(n25772), .B2(n25916), .ZN(
        n7468) );
  OAI22_X1 U21761 ( .A1(n9432), .A2(n25778), .B1(n25772), .B2(n25919), .ZN(
        n7469) );
  OAI22_X1 U21762 ( .A1(n9431), .A2(n25779), .B1(n25772), .B2(n25922), .ZN(
        n7470) );
  OAI22_X1 U21763 ( .A1(n9430), .A2(n25779), .B1(n25773), .B2(n25925), .ZN(
        n7471) );
  OAI22_X1 U21764 ( .A1(n9429), .A2(n25779), .B1(n25773), .B2(n25928), .ZN(
        n7472) );
  OAI22_X1 U21765 ( .A1(n9428), .A2(n25779), .B1(n25773), .B2(n25931), .ZN(
        n7473) );
  OAI22_X1 U21766 ( .A1(n9427), .A2(n25779), .B1(n25773), .B2(n25934), .ZN(
        n7474) );
  OAI22_X1 U21767 ( .A1(n9426), .A2(n25779), .B1(n25773), .B2(n25937), .ZN(
        n7475) );
  OAI22_X1 U21768 ( .A1(n9425), .A2(n25779), .B1(n25773), .B2(n25940), .ZN(
        n7476) );
  OAI22_X1 U21769 ( .A1(n9424), .A2(n25779), .B1(n25773), .B2(n25943), .ZN(
        n7477) );
  OAI22_X1 U21770 ( .A1(n9423), .A2(n25779), .B1(n25773), .B2(n25946), .ZN(
        n7478) );
  OAI22_X1 U21771 ( .A1(n9422), .A2(n25779), .B1(n25773), .B2(n25949), .ZN(
        n7479) );
  OAI22_X1 U21772 ( .A1(n9421), .A2(n25779), .B1(n25773), .B2(n25952), .ZN(
        n7480) );
  OAI22_X1 U21773 ( .A1(n9420), .A2(n25779), .B1(n25773), .B2(n25955), .ZN(
        n7481) );
  OAI22_X1 U21774 ( .A1(n9419), .A2(n25780), .B1(n25773), .B2(n25958), .ZN(
        n7482) );
  OAI22_X1 U21775 ( .A1(n9418), .A2(n25780), .B1(n25774), .B2(n25961), .ZN(
        n7483) );
  OAI22_X1 U21776 ( .A1(n9417), .A2(n25780), .B1(n25774), .B2(n25964), .ZN(
        n7484) );
  OAI22_X1 U21777 ( .A1(n9416), .A2(n25780), .B1(n25774), .B2(n25967), .ZN(
        n7485) );
  OAI22_X1 U21778 ( .A1(n9415), .A2(n25780), .B1(n25774), .B2(n25970), .ZN(
        n7486) );
  OAI22_X1 U21779 ( .A1(n25601), .A2(n21417), .B1(n25962), .B2(n25594), .ZN(
        n6587) );
  OAI22_X1 U21780 ( .A1(n25601), .A2(n21416), .B1(n25965), .B2(n25594), .ZN(
        n6588) );
  OAI22_X1 U21781 ( .A1(n25601), .A2(n21415), .B1(n25968), .B2(n25594), .ZN(
        n6589) );
  OAI22_X1 U21782 ( .A1(n25601), .A2(n21414), .B1(n25971), .B2(n25594), .ZN(
        n6590) );
  OAI22_X1 U21783 ( .A1(n25473), .A2(n21289), .B1(n25962), .B2(n25466), .ZN(
        n5947) );
  OAI22_X1 U21784 ( .A1(n25473), .A2(n21288), .B1(n25965), .B2(n25466), .ZN(
        n5948) );
  OAI22_X1 U21785 ( .A1(n25473), .A2(n21287), .B1(n25968), .B2(n25466), .ZN(
        n5949) );
  OAI22_X1 U21786 ( .A1(n25473), .A2(n21286), .B1(n25971), .B2(n25466), .ZN(
        n5950) );
  OAI22_X1 U21787 ( .A1(n25486), .A2(n21033), .B1(n25962), .B2(n25479), .ZN(
        n6011) );
  OAI22_X1 U21788 ( .A1(n25486), .A2(n21032), .B1(n25965), .B2(n25479), .ZN(
        n6012) );
  OAI22_X1 U21789 ( .A1(n25486), .A2(n21031), .B1(n25968), .B2(n25479), .ZN(
        n6013) );
  OAI22_X1 U21790 ( .A1(n25486), .A2(n21030), .B1(n25971), .B2(n25479), .ZN(
        n6014) );
  OAI22_X1 U21791 ( .A1(n25576), .A2(n20905), .B1(n25962), .B2(n25569), .ZN(
        n6459) );
  OAI22_X1 U21792 ( .A1(n25576), .A2(n20904), .B1(n25965), .B2(n25569), .ZN(
        n6460) );
  OAI22_X1 U21793 ( .A1(n25576), .A2(n20903), .B1(n25968), .B2(n25569), .ZN(
        n6461) );
  OAI22_X1 U21794 ( .A1(n25576), .A2(n20902), .B1(n25971), .B2(n25569), .ZN(
        n6462) );
  OAI22_X1 U21795 ( .A1(n25460), .A2(n20781), .B1(n25963), .B2(n25453), .ZN(
        n5883) );
  OAI22_X1 U21796 ( .A1(n25460), .A2(n20780), .B1(n25966), .B2(n25453), .ZN(
        n5884) );
  OAI22_X1 U21797 ( .A1(n25460), .A2(n20779), .B1(n25969), .B2(n25453), .ZN(
        n5885) );
  OAI22_X1 U21798 ( .A1(n25460), .A2(n20778), .B1(n25972), .B2(n25453), .ZN(
        n5886) );
  OAI22_X1 U21799 ( .A1(n25653), .A2(n20585), .B1(n25961), .B2(n25646), .ZN(
        n6843) );
  OAI22_X1 U21800 ( .A1(n25653), .A2(n20584), .B1(n25964), .B2(n25646), .ZN(
        n6844) );
  OAI22_X1 U21801 ( .A1(n25653), .A2(n20583), .B1(n25967), .B2(n25646), .ZN(
        n6845) );
  OAI22_X1 U21802 ( .A1(n25653), .A2(n20582), .B1(n25970), .B2(n25646), .ZN(
        n6846) );
  OAI22_X1 U21803 ( .A1(n25421), .A2(n20269), .B1(n25963), .B2(n25414), .ZN(
        n5691) );
  OAI22_X1 U21804 ( .A1(n25421), .A2(n20268), .B1(n25966), .B2(n25414), .ZN(
        n5692) );
  OAI22_X1 U21805 ( .A1(n25421), .A2(n20267), .B1(n25969), .B2(n25414), .ZN(
        n5693) );
  OAI22_X1 U21806 ( .A1(n25421), .A2(n20266), .B1(n25972), .B2(n25414), .ZN(
        n5694) );
  OAI22_X1 U21807 ( .A1(n25395), .A2(n20265), .B1(n25963), .B2(n25388), .ZN(
        n5563) );
  OAI22_X1 U21808 ( .A1(n25395), .A2(n20264), .B1(n25966), .B2(n25388), .ZN(
        n5564) );
  OAI22_X1 U21809 ( .A1(n25395), .A2(n20263), .B1(n25969), .B2(n25388), .ZN(
        n5565) );
  OAI22_X1 U21810 ( .A1(n25395), .A2(n20262), .B1(n25972), .B2(n25388), .ZN(
        n5566) );
  OAI22_X1 U21811 ( .A1(n25743), .A2(n20201), .B1(n25961), .B2(n25736), .ZN(
        n7291) );
  OAI22_X1 U21812 ( .A1(n25743), .A2(n20200), .B1(n25964), .B2(n25736), .ZN(
        n7292) );
  OAI22_X1 U21813 ( .A1(n25743), .A2(n20199), .B1(n25967), .B2(n25736), .ZN(
        n7293) );
  OAI22_X1 U21814 ( .A1(n25743), .A2(n20198), .B1(n25970), .B2(n25736), .ZN(
        n7294) );
  OAI22_X1 U21815 ( .A1(n9226), .A2(n25588), .B1(n25962), .B2(n25582), .ZN(
        n6523) );
  OAI22_X1 U21816 ( .A1(n9225), .A2(n25588), .B1(n25965), .B2(n25582), .ZN(
        n6524) );
  OAI22_X1 U21817 ( .A1(n9224), .A2(n25588), .B1(n25968), .B2(n25582), .ZN(
        n6525) );
  OAI22_X1 U21818 ( .A1(n9223), .A2(n25588), .B1(n25971), .B2(n25582), .ZN(
        n6526) );
  OAI22_X1 U21819 ( .A1(n8970), .A2(n25511), .B1(n25962), .B2(n25505), .ZN(
        n6139) );
  OAI22_X1 U21820 ( .A1(n8969), .A2(n25511), .B1(n25965), .B2(n25505), .ZN(
        n6140) );
  OAI22_X1 U21821 ( .A1(n8968), .A2(n25511), .B1(n25968), .B2(n25505), .ZN(
        n6141) );
  OAI22_X1 U21822 ( .A1(n8967), .A2(n25511), .B1(n25971), .B2(n25505), .ZN(
        n6142) );
  OAI22_X1 U21823 ( .A1(n9034), .A2(n25755), .B1(n25961), .B2(n25749), .ZN(
        n7355) );
  OAI22_X1 U21824 ( .A1(n9033), .A2(n25755), .B1(n25964), .B2(n25749), .ZN(
        n7356) );
  OAI22_X1 U21825 ( .A1(n9032), .A2(n25755), .B1(n25967), .B2(n25749), .ZN(
        n7357) );
  OAI22_X1 U21826 ( .A1(n9031), .A2(n25755), .B1(n25970), .B2(n25749), .ZN(
        n7358) );
  OAI22_X1 U21827 ( .A1(n9290), .A2(n25691), .B1(n25961), .B2(n25685), .ZN(
        n7035) );
  OAI22_X1 U21828 ( .A1(n9289), .A2(n25691), .B1(n25964), .B2(n25685), .ZN(
        n7036) );
  OAI22_X1 U21829 ( .A1(n9288), .A2(n25691), .B1(n25967), .B2(n25685), .ZN(
        n7037) );
  OAI22_X1 U21830 ( .A1(n9287), .A2(n25691), .B1(n25970), .B2(n25685), .ZN(
        n7038) );
  OAI22_X1 U21831 ( .A1(n25499), .A2(n19880), .B1(n25962), .B2(n25492), .ZN(
        n6075) );
  OAI22_X1 U21832 ( .A1(n25499), .A2(n19879), .B1(n25965), .B2(n25492), .ZN(
        n6076) );
  OAI22_X1 U21833 ( .A1(n25499), .A2(n19878), .B1(n25968), .B2(n25492), .ZN(
        n6077) );
  OAI22_X1 U21834 ( .A1(n25499), .A2(n19877), .B1(n25971), .B2(n25492), .ZN(
        n6078) );
  OAI22_X1 U21835 ( .A1(n25679), .A2(n19689), .B1(n25961), .B2(n25672), .ZN(
        n6971) );
  OAI22_X1 U21836 ( .A1(n25679), .A2(n19688), .B1(n25964), .B2(n25672), .ZN(
        n6972) );
  OAI22_X1 U21837 ( .A1(n25679), .A2(n19687), .B1(n25967), .B2(n25672), .ZN(
        n6973) );
  OAI22_X1 U21838 ( .A1(n25679), .A2(n19686), .B1(n25970), .B2(n25672), .ZN(
        n6974) );
  OAI22_X1 U21839 ( .A1(n25704), .A2(n19625), .B1(n25961), .B2(n25697), .ZN(
        n7099) );
  OAI22_X1 U21840 ( .A1(n25704), .A2(n19624), .B1(n25964), .B2(n25697), .ZN(
        n7100) );
  OAI22_X1 U21841 ( .A1(n25704), .A2(n19623), .B1(n25967), .B2(n25697), .ZN(
        n7101) );
  OAI22_X1 U21842 ( .A1(n25704), .A2(n19622), .B1(n25970), .B2(n25697), .ZN(
        n7102) );
  AOI22_X1 U21843 ( .A1(n24985), .A2(n19941), .B1(n24979), .B2(n24477), .ZN(
        n22801) );
  AOI22_X1 U21844 ( .A1(n24980), .A2(n20004), .B1(n24974), .B2(n24794), .ZN(
        n23949) );
  AOI22_X1 U21845 ( .A1(n24980), .A2(n20003), .B1(n24974), .B2(n24795), .ZN(
        n23919) );
  AOI22_X1 U21846 ( .A1(n24980), .A2(n20002), .B1(n24974), .B2(n24796), .ZN(
        n23901) );
  AOI22_X1 U21847 ( .A1(n24980), .A2(n20001), .B1(n24974), .B2(n24797), .ZN(
        n23883) );
  AOI22_X1 U21848 ( .A1(n24980), .A2(n20000), .B1(n24974), .B2(n24798), .ZN(
        n23865) );
  AOI22_X1 U21849 ( .A1(n24980), .A2(n19999), .B1(n24974), .B2(n24799), .ZN(
        n23847) );
  AOI22_X1 U21850 ( .A1(n24980), .A2(n19998), .B1(n24974), .B2(n24800), .ZN(
        n23829) );
  AOI22_X1 U21851 ( .A1(n24980), .A2(n19997), .B1(n24974), .B2(n24801), .ZN(
        n23811) );
  AOI22_X1 U21852 ( .A1(n24980), .A2(n19996), .B1(n24974), .B2(n24802), .ZN(
        n23793) );
  AOI22_X1 U21853 ( .A1(n24980), .A2(n19995), .B1(n24974), .B2(n24803), .ZN(
        n23775) );
  AOI22_X1 U21854 ( .A1(n24980), .A2(n19994), .B1(n24974), .B2(n24804), .ZN(
        n23757) );
  AOI22_X1 U21855 ( .A1(n24980), .A2(n19993), .B1(n24974), .B2(n24805), .ZN(
        n23739) );
  AOI22_X1 U21856 ( .A1(n24981), .A2(n19992), .B1(n24975), .B2(n24806), .ZN(
        n23721) );
  AOI22_X1 U21857 ( .A1(n24981), .A2(n19991), .B1(n24975), .B2(n24807), .ZN(
        n23703) );
  AOI22_X1 U21858 ( .A1(n24981), .A2(n19990), .B1(n24975), .B2(n24808), .ZN(
        n23685) );
  AOI22_X1 U21859 ( .A1(n24981), .A2(n19989), .B1(n24975), .B2(n24809), .ZN(
        n23667) );
  AOI22_X1 U21860 ( .A1(n24981), .A2(n19988), .B1(n24975), .B2(n24810), .ZN(
        n23649) );
  AOI22_X1 U21861 ( .A1(n24981), .A2(n19987), .B1(n24975), .B2(n24811), .ZN(
        n23631) );
  AOI22_X1 U21862 ( .A1(n24981), .A2(n19986), .B1(n24975), .B2(n24812), .ZN(
        n23613) );
  AOI22_X1 U21863 ( .A1(n24981), .A2(n19985), .B1(n24975), .B2(n24813), .ZN(
        n23595) );
  AOI22_X1 U21864 ( .A1(n24981), .A2(n19984), .B1(n24975), .B2(n24814), .ZN(
        n23577) );
  AOI22_X1 U21865 ( .A1(n24981), .A2(n19983), .B1(n24975), .B2(n24815), .ZN(
        n23559) );
  AOI22_X1 U21866 ( .A1(n24981), .A2(n19982), .B1(n24975), .B2(n24816), .ZN(
        n23541) );
  AOI22_X1 U21867 ( .A1(n24981), .A2(n19981), .B1(n24975), .B2(n24817), .ZN(
        n23523) );
  AOI22_X1 U21868 ( .A1(n24982), .A2(n19980), .B1(n24976), .B2(n24818), .ZN(
        n23505) );
  AOI22_X1 U21869 ( .A1(n24982), .A2(n19979), .B1(n24976), .B2(n24819), .ZN(
        n23487) );
  AOI22_X1 U21870 ( .A1(n24982), .A2(n19978), .B1(n24976), .B2(n24820), .ZN(
        n23469) );
  AOI22_X1 U21871 ( .A1(n24982), .A2(n19977), .B1(n24976), .B2(n24821), .ZN(
        n23451) );
  AOI22_X1 U21872 ( .A1(n24982), .A2(n19976), .B1(n24976), .B2(n24822), .ZN(
        n23433) );
  AOI22_X1 U21873 ( .A1(n24982), .A2(n19975), .B1(n24976), .B2(n24823), .ZN(
        n23415) );
  AOI22_X1 U21874 ( .A1(n24982), .A2(n19974), .B1(n24976), .B2(n24824), .ZN(
        n23397) );
  AOI22_X1 U21875 ( .A1(n24982), .A2(n19973), .B1(n24976), .B2(n24825), .ZN(
        n23379) );
  AOI22_X1 U21876 ( .A1(n24982), .A2(n19972), .B1(n24976), .B2(n24826), .ZN(
        n23361) );
  AOI22_X1 U21877 ( .A1(n24982), .A2(n19971), .B1(n24976), .B2(n24827), .ZN(
        n23343) );
  AOI22_X1 U21878 ( .A1(n24982), .A2(n19970), .B1(n24976), .B2(n24828), .ZN(
        n23325) );
  AOI22_X1 U21879 ( .A1(n24982), .A2(n19969), .B1(n24976), .B2(n24829), .ZN(
        n23307) );
  AOI22_X1 U21880 ( .A1(n24983), .A2(n19968), .B1(n24977), .B2(n24830), .ZN(
        n23289) );
  AOI22_X1 U21881 ( .A1(n24983), .A2(n19967), .B1(n24977), .B2(n24831), .ZN(
        n23271) );
  AOI22_X1 U21882 ( .A1(n24983), .A2(n19966), .B1(n24977), .B2(n24832), .ZN(
        n23253) );
  AOI22_X1 U21883 ( .A1(n24983), .A2(n19965), .B1(n24977), .B2(n24833), .ZN(
        n23235) );
  AOI22_X1 U21884 ( .A1(n24983), .A2(n19964), .B1(n24977), .B2(n24834), .ZN(
        n23217) );
  AOI22_X1 U21885 ( .A1(n24983), .A2(n19963), .B1(n24977), .B2(n24835), .ZN(
        n23199) );
  AOI22_X1 U21886 ( .A1(n24983), .A2(n19962), .B1(n24977), .B2(n24836), .ZN(
        n23181) );
  AOI22_X1 U21887 ( .A1(n24983), .A2(n19961), .B1(n24977), .B2(n24837), .ZN(
        n23163) );
  AOI22_X1 U21888 ( .A1(n24983), .A2(n19960), .B1(n24977), .B2(n24838), .ZN(
        n23145) );
  AOI22_X1 U21889 ( .A1(n24983), .A2(n19959), .B1(n24977), .B2(n24839), .ZN(
        n23127) );
  AOI22_X1 U21890 ( .A1(n24983), .A2(n19958), .B1(n24977), .B2(n24840), .ZN(
        n23109) );
  AOI22_X1 U21891 ( .A1(n24983), .A2(n19957), .B1(n24977), .B2(n24841), .ZN(
        n23091) );
  AOI22_X1 U21892 ( .A1(n24984), .A2(n19956), .B1(n24978), .B2(n24842), .ZN(
        n23073) );
  AOI22_X1 U21893 ( .A1(n24984), .A2(n19955), .B1(n24978), .B2(n24843), .ZN(
        n23055) );
  AOI22_X1 U21894 ( .A1(n24984), .A2(n19954), .B1(n24978), .B2(n24844), .ZN(
        n23037) );
  AOI22_X1 U21895 ( .A1(n24984), .A2(n19953), .B1(n24978), .B2(n24845), .ZN(
        n23019) );
  AOI22_X1 U21896 ( .A1(n24984), .A2(n19952), .B1(n24978), .B2(n24846), .ZN(
        n23001) );
  AOI22_X1 U21897 ( .A1(n24984), .A2(n19951), .B1(n24978), .B2(n24847), .ZN(
        n22983) );
  AOI22_X1 U21898 ( .A1(n24984), .A2(n19950), .B1(n24978), .B2(n24848), .ZN(
        n22965) );
  AOI22_X1 U21899 ( .A1(n24984), .A2(n19949), .B1(n24978), .B2(n24849), .ZN(
        n22947) );
  AOI22_X1 U21900 ( .A1(n24984), .A2(n19948), .B1(n24978), .B2(n24850), .ZN(
        n22929) );
  AOI22_X1 U21901 ( .A1(n24984), .A2(n19947), .B1(n24978), .B2(n24851), .ZN(
        n22911) );
  AOI22_X1 U21902 ( .A1(n24984), .A2(n19946), .B1(n24978), .B2(n24852), .ZN(
        n22893) );
  AOI22_X1 U21903 ( .A1(n24984), .A2(n19945), .B1(n24978), .B2(n24853), .ZN(
        n22875) );
  AOI22_X1 U21904 ( .A1(n24985), .A2(n19944), .B1(n24979), .B2(n24474), .ZN(
        n22857) );
  AOI22_X1 U21905 ( .A1(n24985), .A2(n19943), .B1(n24979), .B2(n24475), .ZN(
        n22839) );
  AOI22_X1 U21906 ( .A1(n24985), .A2(n19942), .B1(n24979), .B2(n24476), .ZN(
        n22821) );
  AOI22_X1 U21907 ( .A1(n25178), .A2(n20004), .B1(n25172), .B2(n24794), .ZN(
        n22752) );
  AOI22_X1 U21908 ( .A1(n25178), .A2(n20003), .B1(n25172), .B2(n24795), .ZN(
        n22722) );
  AOI22_X1 U21909 ( .A1(n25178), .A2(n20002), .B1(n25172), .B2(n24796), .ZN(
        n22704) );
  AOI22_X1 U21910 ( .A1(n25178), .A2(n20001), .B1(n25172), .B2(n24797), .ZN(
        n22686) );
  AOI22_X1 U21911 ( .A1(n25178), .A2(n20000), .B1(n25172), .B2(n24798), .ZN(
        n22668) );
  AOI22_X1 U21912 ( .A1(n25178), .A2(n19999), .B1(n25172), .B2(n24799), .ZN(
        n22650) );
  AOI22_X1 U21913 ( .A1(n25178), .A2(n19998), .B1(n25172), .B2(n24800), .ZN(
        n22632) );
  AOI22_X1 U21914 ( .A1(n25178), .A2(n19997), .B1(n25172), .B2(n24801), .ZN(
        n22614) );
  AOI22_X1 U21915 ( .A1(n25178), .A2(n19996), .B1(n25172), .B2(n24802), .ZN(
        n22596) );
  AOI22_X1 U21916 ( .A1(n25178), .A2(n19995), .B1(n25172), .B2(n24803), .ZN(
        n22578) );
  AOI22_X1 U21917 ( .A1(n25178), .A2(n19994), .B1(n25172), .B2(n24804), .ZN(
        n22560) );
  AOI22_X1 U21918 ( .A1(n25178), .A2(n19993), .B1(n25172), .B2(n24805), .ZN(
        n22542) );
  AOI22_X1 U21919 ( .A1(n25179), .A2(n19992), .B1(n25173), .B2(n24806), .ZN(
        n22524) );
  AOI22_X1 U21920 ( .A1(n25179), .A2(n19991), .B1(n25173), .B2(n24807), .ZN(
        n22506) );
  AOI22_X1 U21921 ( .A1(n25179), .A2(n19990), .B1(n25173), .B2(n24808), .ZN(
        n22488) );
  AOI22_X1 U21922 ( .A1(n25179), .A2(n19989), .B1(n25173), .B2(n24809), .ZN(
        n22470) );
  AOI22_X1 U21923 ( .A1(n25179), .A2(n19988), .B1(n25173), .B2(n24810), .ZN(
        n22452) );
  AOI22_X1 U21924 ( .A1(n25179), .A2(n19987), .B1(n25173), .B2(n24811), .ZN(
        n22434) );
  AOI22_X1 U21925 ( .A1(n25179), .A2(n19986), .B1(n25173), .B2(n24812), .ZN(
        n22416) );
  AOI22_X1 U21926 ( .A1(n25179), .A2(n19985), .B1(n25173), .B2(n24813), .ZN(
        n22398) );
  AOI22_X1 U21927 ( .A1(n25179), .A2(n19984), .B1(n25173), .B2(n24814), .ZN(
        n22380) );
  AOI22_X1 U21928 ( .A1(n25179), .A2(n19983), .B1(n25173), .B2(n24815), .ZN(
        n22362) );
  AOI22_X1 U21929 ( .A1(n25179), .A2(n19982), .B1(n25173), .B2(n24816), .ZN(
        n22344) );
  AOI22_X1 U21930 ( .A1(n25179), .A2(n19981), .B1(n25173), .B2(n24817), .ZN(
        n22326) );
  AOI22_X1 U21931 ( .A1(n25180), .A2(n19980), .B1(n25174), .B2(n24818), .ZN(
        n22308) );
  AOI22_X1 U21932 ( .A1(n25180), .A2(n19979), .B1(n25174), .B2(n24819), .ZN(
        n22290) );
  AOI22_X1 U21933 ( .A1(n25180), .A2(n19978), .B1(n25174), .B2(n24820), .ZN(
        n22272) );
  AOI22_X1 U21934 ( .A1(n25180), .A2(n19977), .B1(n25174), .B2(n24821), .ZN(
        n22254) );
  AOI22_X1 U21935 ( .A1(n25180), .A2(n19976), .B1(n25174), .B2(n24822), .ZN(
        n22236) );
  AOI22_X1 U21936 ( .A1(n25180), .A2(n19975), .B1(n25174), .B2(n24823), .ZN(
        n22218) );
  AOI22_X1 U21937 ( .A1(n25180), .A2(n19974), .B1(n25174), .B2(n24824), .ZN(
        n22200) );
  AOI22_X1 U21938 ( .A1(n25180), .A2(n19973), .B1(n25174), .B2(n24825), .ZN(
        n22182) );
  AOI22_X1 U21939 ( .A1(n25180), .A2(n19972), .B1(n25174), .B2(n24826), .ZN(
        n22164) );
  AOI22_X1 U21940 ( .A1(n25180), .A2(n19971), .B1(n25174), .B2(n24827), .ZN(
        n22146) );
  AOI22_X1 U21941 ( .A1(n25180), .A2(n19970), .B1(n25174), .B2(n24828), .ZN(
        n22128) );
  AOI22_X1 U21942 ( .A1(n25180), .A2(n19969), .B1(n25174), .B2(n24829), .ZN(
        n22110) );
  AOI22_X1 U21943 ( .A1(n25181), .A2(n19968), .B1(n25175), .B2(n24830), .ZN(
        n22092) );
  AOI22_X1 U21944 ( .A1(n25181), .A2(n19967), .B1(n25175), .B2(n24831), .ZN(
        n22074) );
  AOI22_X1 U21945 ( .A1(n25181), .A2(n19966), .B1(n25175), .B2(n24832), .ZN(
        n22056) );
  AOI22_X1 U21946 ( .A1(n25181), .A2(n19965), .B1(n25175), .B2(n24833), .ZN(
        n22038) );
  AOI22_X1 U21947 ( .A1(n25181), .A2(n19964), .B1(n25175), .B2(n24834), .ZN(
        n22020) );
  AOI22_X1 U21948 ( .A1(n25181), .A2(n19963), .B1(n25175), .B2(n24835), .ZN(
        n22002) );
  AOI22_X1 U21949 ( .A1(n25181), .A2(n19962), .B1(n25175), .B2(n24836), .ZN(
        n21984) );
  AOI22_X1 U21950 ( .A1(n25181), .A2(n19961), .B1(n25175), .B2(n24837), .ZN(
        n21966) );
  AOI22_X1 U21951 ( .A1(n25181), .A2(n19960), .B1(n25175), .B2(n24838), .ZN(
        n21948) );
  AOI22_X1 U21952 ( .A1(n25181), .A2(n19959), .B1(n25175), .B2(n24839), .ZN(
        n21930) );
  AOI22_X1 U21953 ( .A1(n25181), .A2(n19958), .B1(n25175), .B2(n24840), .ZN(
        n21912) );
  AOI22_X1 U21954 ( .A1(n25181), .A2(n19957), .B1(n25175), .B2(n24841), .ZN(
        n21894) );
  AOI22_X1 U21955 ( .A1(n25182), .A2(n19956), .B1(n25176), .B2(n24842), .ZN(
        n21876) );
  AOI22_X1 U21956 ( .A1(n25182), .A2(n19955), .B1(n25176), .B2(n24843), .ZN(
        n21858) );
  AOI22_X1 U21957 ( .A1(n25182), .A2(n19954), .B1(n25176), .B2(n24844), .ZN(
        n21840) );
  AOI22_X1 U21958 ( .A1(n25182), .A2(n19953), .B1(n25176), .B2(n24845), .ZN(
        n21822) );
  AOI22_X1 U21959 ( .A1(n25182), .A2(n19952), .B1(n25176), .B2(n24846), .ZN(
        n21804) );
  AOI22_X1 U21960 ( .A1(n25182), .A2(n19951), .B1(n25176), .B2(n24847), .ZN(
        n21786) );
  AOI22_X1 U21961 ( .A1(n25182), .A2(n19950), .B1(n25176), .B2(n24848), .ZN(
        n21768) );
  AOI22_X1 U21962 ( .A1(n25182), .A2(n19949), .B1(n25176), .B2(n24849), .ZN(
        n21750) );
  AOI22_X1 U21963 ( .A1(n25182), .A2(n19948), .B1(n25176), .B2(n24850), .ZN(
        n21732) );
  AOI22_X1 U21964 ( .A1(n25182), .A2(n19947), .B1(n25176), .B2(n24851), .ZN(
        n21714) );
  AOI22_X1 U21965 ( .A1(n25182), .A2(n19946), .B1(n25176), .B2(n24852), .ZN(
        n21696) );
  AOI22_X1 U21966 ( .A1(n25182), .A2(n19945), .B1(n25176), .B2(n24853), .ZN(
        n21678) );
  AOI22_X1 U21967 ( .A1(n25183), .A2(n19944), .B1(n25177), .B2(n24474), .ZN(
        n21660) );
  AOI22_X1 U21968 ( .A1(n25183), .A2(n19943), .B1(n25177), .B2(n24475), .ZN(
        n21642) );
  AOI22_X1 U21969 ( .A1(n25183), .A2(n19942), .B1(n25177), .B2(n24476), .ZN(
        n21624) );
  AOI22_X1 U21970 ( .A1(n25183), .A2(n19941), .B1(n25177), .B2(n24477), .ZN(
        n21604) );
  OAI221_X1 U21971 ( .B1(n21285), .B2(n25118), .C1(n19621), .C2(n25112), .A(
        n23936), .ZN(n23923) );
  AOI22_X1 U21972 ( .A1(n25106), .A2(n24854), .B1(n25100), .B2(n20068), .ZN(
        n23936) );
  OAI221_X1 U21973 ( .B1(n21221), .B2(n25064), .C1(n20197), .C2(n25058), .A(
        n23945), .ZN(n23944) );
  AOI22_X1 U21974 ( .A1(n25052), .A2(n24087), .B1(n25046), .B2(OUT2[0]), .ZN(
        n23945) );
  OAI221_X1 U21975 ( .B1(n21284), .B2(n25118), .C1(n19620), .C2(n25112), .A(
        n23910), .ZN(n23905) );
  AOI22_X1 U21976 ( .A1(n25106), .A2(n24855), .B1(n25100), .B2(n20067), .ZN(
        n23910) );
  OAI221_X1 U21977 ( .B1(n21220), .B2(n25064), .C1(n20196), .C2(n25058), .A(
        n23916), .ZN(n23915) );
  AOI22_X1 U21978 ( .A1(n25052), .A2(n24089), .B1(n25051), .B2(OUT2[1]), .ZN(
        n23916) );
  OAI221_X1 U21979 ( .B1(n21283), .B2(n25118), .C1(n19619), .C2(n25112), .A(
        n23892), .ZN(n23887) );
  AOI22_X1 U21980 ( .A1(n25106), .A2(n24856), .B1(n25100), .B2(n20066), .ZN(
        n23892) );
  OAI221_X1 U21981 ( .B1(n21219), .B2(n25064), .C1(n20195), .C2(n25058), .A(
        n23898), .ZN(n23897) );
  AOI22_X1 U21982 ( .A1(n25052), .A2(n24091), .B1(n25051), .B2(OUT2[2]), .ZN(
        n23898) );
  OAI221_X1 U21983 ( .B1(n21282), .B2(n25118), .C1(n19618), .C2(n25112), .A(
        n23874), .ZN(n23869) );
  AOI22_X1 U21984 ( .A1(n25106), .A2(n24857), .B1(n25100), .B2(n20065), .ZN(
        n23874) );
  OAI221_X1 U21985 ( .B1(n21218), .B2(n25064), .C1(n20194), .C2(n25058), .A(
        n23880), .ZN(n23879) );
  AOI22_X1 U21986 ( .A1(n25052), .A2(n24093), .B1(n25051), .B2(OUT2[3]), .ZN(
        n23880) );
  OAI221_X1 U21987 ( .B1(n21281), .B2(n25118), .C1(n19617), .C2(n25112), .A(
        n23856), .ZN(n23851) );
  AOI22_X1 U21988 ( .A1(n25106), .A2(n24858), .B1(n25100), .B2(n20064), .ZN(
        n23856) );
  OAI221_X1 U21989 ( .B1(n21217), .B2(n25064), .C1(n20193), .C2(n25058), .A(
        n23862), .ZN(n23861) );
  AOI22_X1 U21990 ( .A1(n25052), .A2(n24095), .B1(n25050), .B2(OUT2[4]), .ZN(
        n23862) );
  OAI221_X1 U21991 ( .B1(n21280), .B2(n25118), .C1(n19616), .C2(n25112), .A(
        n23838), .ZN(n23833) );
  AOI22_X1 U21992 ( .A1(n25106), .A2(n24859), .B1(n25100), .B2(n20063), .ZN(
        n23838) );
  OAI221_X1 U21993 ( .B1(n21216), .B2(n25064), .C1(n20192), .C2(n25058), .A(
        n23844), .ZN(n23843) );
  AOI22_X1 U21994 ( .A1(n25052), .A2(n24097), .B1(n25050), .B2(OUT2[5]), .ZN(
        n23844) );
  OAI221_X1 U21995 ( .B1(n21279), .B2(n25118), .C1(n19615), .C2(n25112), .A(
        n23820), .ZN(n23815) );
  AOI22_X1 U21996 ( .A1(n25106), .A2(n24860), .B1(n25100), .B2(n20062), .ZN(
        n23820) );
  OAI221_X1 U21997 ( .B1(n21215), .B2(n25064), .C1(n20191), .C2(n25058), .A(
        n23826), .ZN(n23825) );
  AOI22_X1 U21998 ( .A1(n25052), .A2(n24099), .B1(n25050), .B2(OUT2[6]), .ZN(
        n23826) );
  OAI221_X1 U21999 ( .B1(n21278), .B2(n25118), .C1(n19614), .C2(n25112), .A(
        n23802), .ZN(n23797) );
  AOI22_X1 U22000 ( .A1(n25106), .A2(n24861), .B1(n25100), .B2(n20061), .ZN(
        n23802) );
  OAI221_X1 U22001 ( .B1(n21214), .B2(n25064), .C1(n20190), .C2(n25058), .A(
        n23808), .ZN(n23807) );
  AOI22_X1 U22002 ( .A1(n25052), .A2(n24101), .B1(n25050), .B2(OUT2[7]), .ZN(
        n23808) );
  OAI221_X1 U22003 ( .B1(n21277), .B2(n25118), .C1(n19613), .C2(n25112), .A(
        n23784), .ZN(n23779) );
  AOI22_X1 U22004 ( .A1(n25106), .A2(n24862), .B1(n25100), .B2(n20060), .ZN(
        n23784) );
  OAI221_X1 U22005 ( .B1(n21213), .B2(n25064), .C1(n20189), .C2(n25058), .A(
        n23790), .ZN(n23789) );
  AOI22_X1 U22006 ( .A1(n25052), .A2(n24103), .B1(n25050), .B2(OUT2[8]), .ZN(
        n23790) );
  OAI221_X1 U22007 ( .B1(n21276), .B2(n25118), .C1(n19612), .C2(n25112), .A(
        n23766), .ZN(n23761) );
  AOI22_X1 U22008 ( .A1(n25106), .A2(n24863), .B1(n25100), .B2(n20059), .ZN(
        n23766) );
  OAI221_X1 U22009 ( .B1(n21212), .B2(n25064), .C1(n20188), .C2(n25058), .A(
        n23772), .ZN(n23771) );
  AOI22_X1 U22010 ( .A1(n25052), .A2(n24105), .B1(n25050), .B2(OUT2[9]), .ZN(
        n23772) );
  OAI221_X1 U22011 ( .B1(n21275), .B2(n25118), .C1(n19611), .C2(n25112), .A(
        n23748), .ZN(n23743) );
  AOI22_X1 U22012 ( .A1(n25106), .A2(n24864), .B1(n25100), .B2(n20058), .ZN(
        n23748) );
  OAI221_X1 U22013 ( .B1(n21211), .B2(n25064), .C1(n20187), .C2(n25058), .A(
        n23754), .ZN(n23753) );
  AOI22_X1 U22014 ( .A1(n25052), .A2(n24107), .B1(n25050), .B2(OUT2[10]), .ZN(
        n23754) );
  OAI221_X1 U22015 ( .B1(n21274), .B2(n25118), .C1(n19610), .C2(n25112), .A(
        n23730), .ZN(n23725) );
  AOI22_X1 U22016 ( .A1(n25106), .A2(n24865), .B1(n25100), .B2(n20057), .ZN(
        n23730) );
  OAI221_X1 U22017 ( .B1(n21210), .B2(n25064), .C1(n20186), .C2(n25058), .A(
        n23736), .ZN(n23735) );
  AOI22_X1 U22018 ( .A1(n25052), .A2(n24109), .B1(n25050), .B2(OUT2[11]), .ZN(
        n23736) );
  OAI221_X1 U22019 ( .B1(n21273), .B2(n25119), .C1(n19609), .C2(n25113), .A(
        n23712), .ZN(n23707) );
  AOI22_X1 U22020 ( .A1(n25107), .A2(n24866), .B1(n25101), .B2(n20056), .ZN(
        n23712) );
  OAI221_X1 U22021 ( .B1(n21209), .B2(n25065), .C1(n20185), .C2(n25059), .A(
        n23718), .ZN(n23717) );
  AOI22_X1 U22022 ( .A1(n25053), .A2(n24111), .B1(n25050), .B2(OUT2[12]), .ZN(
        n23718) );
  OAI221_X1 U22023 ( .B1(n21272), .B2(n25119), .C1(n19608), .C2(n25113), .A(
        n23694), .ZN(n23689) );
  AOI22_X1 U22024 ( .A1(n25107), .A2(n24867), .B1(n25101), .B2(n20055), .ZN(
        n23694) );
  OAI221_X1 U22025 ( .B1(n21208), .B2(n25065), .C1(n20184), .C2(n25059), .A(
        n23700), .ZN(n23699) );
  AOI22_X1 U22026 ( .A1(n25053), .A2(n24113), .B1(n25050), .B2(OUT2[13]), .ZN(
        n23700) );
  OAI221_X1 U22027 ( .B1(n21271), .B2(n25119), .C1(n19607), .C2(n25113), .A(
        n23676), .ZN(n23671) );
  AOI22_X1 U22028 ( .A1(n25107), .A2(n24868), .B1(n25101), .B2(n20054), .ZN(
        n23676) );
  OAI221_X1 U22029 ( .B1(n21207), .B2(n25065), .C1(n20183), .C2(n25059), .A(
        n23682), .ZN(n23681) );
  AOI22_X1 U22030 ( .A1(n25053), .A2(n24115), .B1(n25050), .B2(OUT2[14]), .ZN(
        n23682) );
  OAI221_X1 U22031 ( .B1(n21270), .B2(n25119), .C1(n19606), .C2(n25113), .A(
        n23658), .ZN(n23653) );
  AOI22_X1 U22032 ( .A1(n25107), .A2(n24869), .B1(n25101), .B2(n20053), .ZN(
        n23658) );
  OAI221_X1 U22033 ( .B1(n21206), .B2(n25065), .C1(n20182), .C2(n25059), .A(
        n23664), .ZN(n23663) );
  AOI22_X1 U22034 ( .A1(n25053), .A2(n24117), .B1(n25050), .B2(OUT2[15]), .ZN(
        n23664) );
  OAI221_X1 U22035 ( .B1(n21269), .B2(n25119), .C1(n19605), .C2(n25113), .A(
        n23640), .ZN(n23635) );
  AOI22_X1 U22036 ( .A1(n25107), .A2(n24870), .B1(n25101), .B2(n20052), .ZN(
        n23640) );
  OAI221_X1 U22037 ( .B1(n21205), .B2(n25065), .C1(n20181), .C2(n25059), .A(
        n23646), .ZN(n23645) );
  AOI22_X1 U22038 ( .A1(n25053), .A2(n24119), .B1(n25050), .B2(OUT2[16]), .ZN(
        n23646) );
  OAI221_X1 U22039 ( .B1(n21268), .B2(n25119), .C1(n19604), .C2(n25113), .A(
        n23622), .ZN(n23617) );
  AOI22_X1 U22040 ( .A1(n25107), .A2(n24871), .B1(n25101), .B2(n20051), .ZN(
        n23622) );
  OAI221_X1 U22041 ( .B1(n21204), .B2(n25065), .C1(n20180), .C2(n25059), .A(
        n23628), .ZN(n23627) );
  AOI22_X1 U22042 ( .A1(n25053), .A2(n24121), .B1(n25049), .B2(OUT2[17]), .ZN(
        n23628) );
  OAI221_X1 U22043 ( .B1(n21267), .B2(n25119), .C1(n19603), .C2(n25113), .A(
        n23604), .ZN(n23599) );
  AOI22_X1 U22044 ( .A1(n25107), .A2(n24872), .B1(n25101), .B2(n20050), .ZN(
        n23604) );
  OAI221_X1 U22045 ( .B1(n21203), .B2(n25065), .C1(n20179), .C2(n25059), .A(
        n23610), .ZN(n23609) );
  AOI22_X1 U22046 ( .A1(n25053), .A2(n24123), .B1(n25049), .B2(OUT2[18]), .ZN(
        n23610) );
  OAI221_X1 U22047 ( .B1(n21266), .B2(n25119), .C1(n19602), .C2(n25113), .A(
        n23586), .ZN(n23581) );
  AOI22_X1 U22048 ( .A1(n25107), .A2(n24873), .B1(n25101), .B2(n20049), .ZN(
        n23586) );
  OAI221_X1 U22049 ( .B1(n21202), .B2(n25065), .C1(n20178), .C2(n25059), .A(
        n23592), .ZN(n23591) );
  AOI22_X1 U22050 ( .A1(n25053), .A2(n24125), .B1(n25049), .B2(OUT2[19]), .ZN(
        n23592) );
  OAI221_X1 U22051 ( .B1(n21265), .B2(n25119), .C1(n19601), .C2(n25113), .A(
        n23568), .ZN(n23563) );
  AOI22_X1 U22052 ( .A1(n25107), .A2(n24874), .B1(n25101), .B2(n20048), .ZN(
        n23568) );
  OAI221_X1 U22053 ( .B1(n21201), .B2(n25065), .C1(n20177), .C2(n25059), .A(
        n23574), .ZN(n23573) );
  AOI22_X1 U22054 ( .A1(n25053), .A2(n24127), .B1(n25049), .B2(OUT2[20]), .ZN(
        n23574) );
  OAI221_X1 U22055 ( .B1(n21264), .B2(n25119), .C1(n19600), .C2(n25113), .A(
        n23550), .ZN(n23545) );
  AOI22_X1 U22056 ( .A1(n25107), .A2(n24875), .B1(n25101), .B2(n20047), .ZN(
        n23550) );
  OAI221_X1 U22057 ( .B1(n21200), .B2(n25065), .C1(n20176), .C2(n25059), .A(
        n23556), .ZN(n23555) );
  AOI22_X1 U22058 ( .A1(n25053), .A2(n24129), .B1(n25049), .B2(OUT2[21]), .ZN(
        n23556) );
  OAI221_X1 U22059 ( .B1(n21263), .B2(n25119), .C1(n19599), .C2(n25113), .A(
        n23532), .ZN(n23527) );
  AOI22_X1 U22060 ( .A1(n25107), .A2(n24876), .B1(n25101), .B2(n20046), .ZN(
        n23532) );
  OAI221_X1 U22061 ( .B1(n21199), .B2(n25065), .C1(n20175), .C2(n25059), .A(
        n23538), .ZN(n23537) );
  AOI22_X1 U22062 ( .A1(n25053), .A2(n24131), .B1(n25049), .B2(OUT2[22]), .ZN(
        n23538) );
  OAI221_X1 U22063 ( .B1(n21262), .B2(n25119), .C1(n19598), .C2(n25113), .A(
        n23514), .ZN(n23509) );
  AOI22_X1 U22064 ( .A1(n25107), .A2(n24877), .B1(n25101), .B2(n20045), .ZN(
        n23514) );
  OAI221_X1 U22065 ( .B1(n21198), .B2(n25065), .C1(n20174), .C2(n25059), .A(
        n23520), .ZN(n23519) );
  AOI22_X1 U22066 ( .A1(n25053), .A2(n24133), .B1(n25049), .B2(OUT2[23]), .ZN(
        n23520) );
  OAI221_X1 U22067 ( .B1(n21261), .B2(n25120), .C1(n19597), .C2(n25114), .A(
        n23496), .ZN(n23491) );
  AOI22_X1 U22068 ( .A1(n25108), .A2(n24878), .B1(n25102), .B2(n20044), .ZN(
        n23496) );
  OAI221_X1 U22069 ( .B1(n21197), .B2(n25066), .C1(n20173), .C2(n25060), .A(
        n23502), .ZN(n23501) );
  AOI22_X1 U22070 ( .A1(n25054), .A2(n24135), .B1(n25049), .B2(OUT2[24]), .ZN(
        n23502) );
  OAI221_X1 U22071 ( .B1(n21260), .B2(n25120), .C1(n19596), .C2(n25114), .A(
        n23478), .ZN(n23473) );
  AOI22_X1 U22072 ( .A1(n25108), .A2(n24879), .B1(n25102), .B2(n20043), .ZN(
        n23478) );
  OAI221_X1 U22073 ( .B1(n21196), .B2(n25066), .C1(n20172), .C2(n25060), .A(
        n23484), .ZN(n23483) );
  AOI22_X1 U22074 ( .A1(n25054), .A2(n24137), .B1(n25049), .B2(OUT2[25]), .ZN(
        n23484) );
  OAI221_X1 U22075 ( .B1(n21259), .B2(n25120), .C1(n19595), .C2(n25114), .A(
        n23460), .ZN(n23455) );
  AOI22_X1 U22076 ( .A1(n25108), .A2(n24880), .B1(n25102), .B2(n20042), .ZN(
        n23460) );
  OAI221_X1 U22077 ( .B1(n21195), .B2(n25066), .C1(n20171), .C2(n25060), .A(
        n23466), .ZN(n23465) );
  AOI22_X1 U22078 ( .A1(n25054), .A2(n24139), .B1(n25049), .B2(OUT2[26]), .ZN(
        n23466) );
  OAI221_X1 U22079 ( .B1(n21258), .B2(n25120), .C1(n19594), .C2(n25114), .A(
        n23442), .ZN(n23437) );
  AOI22_X1 U22080 ( .A1(n25108), .A2(n24881), .B1(n25102), .B2(n20041), .ZN(
        n23442) );
  OAI221_X1 U22081 ( .B1(n21194), .B2(n25066), .C1(n20170), .C2(n25060), .A(
        n23448), .ZN(n23447) );
  AOI22_X1 U22082 ( .A1(n25054), .A2(n24141), .B1(n25049), .B2(OUT2[27]), .ZN(
        n23448) );
  OAI221_X1 U22083 ( .B1(n21257), .B2(n25120), .C1(n19593), .C2(n25114), .A(
        n23424), .ZN(n23419) );
  AOI22_X1 U22084 ( .A1(n25108), .A2(n24882), .B1(n25102), .B2(n20040), .ZN(
        n23424) );
  OAI221_X1 U22085 ( .B1(n21193), .B2(n25066), .C1(n20169), .C2(n25060), .A(
        n23430), .ZN(n23429) );
  AOI22_X1 U22086 ( .A1(n25054), .A2(n24143), .B1(n25049), .B2(OUT2[28]), .ZN(
        n23430) );
  OAI221_X1 U22087 ( .B1(n21256), .B2(n25120), .C1(n19592), .C2(n25114), .A(
        n23406), .ZN(n23401) );
  AOI22_X1 U22088 ( .A1(n25108), .A2(n24883), .B1(n25102), .B2(n20039), .ZN(
        n23406) );
  OAI221_X1 U22089 ( .B1(n21192), .B2(n25066), .C1(n20168), .C2(n25060), .A(
        n23412), .ZN(n23411) );
  AOI22_X1 U22090 ( .A1(n25054), .A2(n24145), .B1(n25049), .B2(OUT2[29]), .ZN(
        n23412) );
  OAI221_X1 U22091 ( .B1(n21255), .B2(n25120), .C1(n19591), .C2(n25114), .A(
        n23388), .ZN(n23383) );
  AOI22_X1 U22092 ( .A1(n25108), .A2(n24884), .B1(n25102), .B2(n20038), .ZN(
        n23388) );
  OAI221_X1 U22093 ( .B1(n21191), .B2(n25066), .C1(n20167), .C2(n25060), .A(
        n23394), .ZN(n23393) );
  AOI22_X1 U22094 ( .A1(n25054), .A2(n24147), .B1(n25048), .B2(OUT2[30]), .ZN(
        n23394) );
  OAI221_X1 U22095 ( .B1(n21254), .B2(n25120), .C1(n19590), .C2(n25114), .A(
        n23370), .ZN(n23365) );
  AOI22_X1 U22096 ( .A1(n25108), .A2(n24885), .B1(n25102), .B2(n20037), .ZN(
        n23370) );
  OAI221_X1 U22097 ( .B1(n21190), .B2(n25066), .C1(n20166), .C2(n25060), .A(
        n23376), .ZN(n23375) );
  AOI22_X1 U22098 ( .A1(n25054), .A2(n24149), .B1(n25048), .B2(OUT2[31]), .ZN(
        n23376) );
  OAI221_X1 U22099 ( .B1(n21253), .B2(n25120), .C1(n19589), .C2(n25114), .A(
        n23352), .ZN(n23347) );
  AOI22_X1 U22100 ( .A1(n25108), .A2(n24886), .B1(n25102), .B2(n20036), .ZN(
        n23352) );
  OAI221_X1 U22101 ( .B1(n21189), .B2(n25066), .C1(n20165), .C2(n25060), .A(
        n23358), .ZN(n23357) );
  AOI22_X1 U22102 ( .A1(n25054), .A2(n24151), .B1(n25048), .B2(OUT2[32]), .ZN(
        n23358) );
  OAI221_X1 U22103 ( .B1(n21252), .B2(n25120), .C1(n19588), .C2(n25114), .A(
        n23334), .ZN(n23329) );
  AOI22_X1 U22104 ( .A1(n25108), .A2(n24887), .B1(n25102), .B2(n20035), .ZN(
        n23334) );
  OAI221_X1 U22105 ( .B1(n21188), .B2(n25066), .C1(n20164), .C2(n25060), .A(
        n23340), .ZN(n23339) );
  AOI22_X1 U22106 ( .A1(n25054), .A2(n24153), .B1(n25048), .B2(OUT2[33]), .ZN(
        n23340) );
  OAI221_X1 U22107 ( .B1(n21251), .B2(n25120), .C1(n19587), .C2(n25114), .A(
        n23316), .ZN(n23311) );
  AOI22_X1 U22108 ( .A1(n25108), .A2(n24888), .B1(n25102), .B2(n20034), .ZN(
        n23316) );
  OAI221_X1 U22109 ( .B1(n21187), .B2(n25066), .C1(n20163), .C2(n25060), .A(
        n23322), .ZN(n23321) );
  AOI22_X1 U22110 ( .A1(n25054), .A2(n24155), .B1(n25048), .B2(OUT2[34]), .ZN(
        n23322) );
  OAI221_X1 U22111 ( .B1(n21250), .B2(n25120), .C1(n19586), .C2(n25114), .A(
        n23298), .ZN(n23293) );
  AOI22_X1 U22112 ( .A1(n25108), .A2(n24889), .B1(n25102), .B2(n20033), .ZN(
        n23298) );
  OAI221_X1 U22113 ( .B1(n21186), .B2(n25066), .C1(n20162), .C2(n25060), .A(
        n23304), .ZN(n23303) );
  AOI22_X1 U22114 ( .A1(n25054), .A2(n24157), .B1(n25048), .B2(OUT2[35]), .ZN(
        n23304) );
  OAI221_X1 U22115 ( .B1(n21249), .B2(n25121), .C1(n19585), .C2(n25115), .A(
        n23280), .ZN(n23275) );
  AOI22_X1 U22116 ( .A1(n25109), .A2(n24890), .B1(n25103), .B2(n20032), .ZN(
        n23280) );
  OAI221_X1 U22117 ( .B1(n21185), .B2(n25067), .C1(n20161), .C2(n25061), .A(
        n23286), .ZN(n23285) );
  AOI22_X1 U22118 ( .A1(n25055), .A2(n24159), .B1(n25048), .B2(OUT2[36]), .ZN(
        n23286) );
  OAI221_X1 U22119 ( .B1(n21248), .B2(n25121), .C1(n19584), .C2(n25115), .A(
        n23262), .ZN(n23257) );
  AOI22_X1 U22120 ( .A1(n25109), .A2(n24891), .B1(n25103), .B2(n20031), .ZN(
        n23262) );
  OAI221_X1 U22121 ( .B1(n21184), .B2(n25067), .C1(n20160), .C2(n25061), .A(
        n23268), .ZN(n23267) );
  AOI22_X1 U22122 ( .A1(n25055), .A2(n24161), .B1(n25048), .B2(OUT2[37]), .ZN(
        n23268) );
  OAI221_X1 U22123 ( .B1(n21247), .B2(n25121), .C1(n19583), .C2(n25115), .A(
        n23244), .ZN(n23239) );
  AOI22_X1 U22124 ( .A1(n25109), .A2(n24892), .B1(n25103), .B2(n20030), .ZN(
        n23244) );
  OAI221_X1 U22125 ( .B1(n21183), .B2(n25067), .C1(n20159), .C2(n25061), .A(
        n23250), .ZN(n23249) );
  AOI22_X1 U22126 ( .A1(n25055), .A2(n24163), .B1(n25048), .B2(OUT2[38]), .ZN(
        n23250) );
  OAI221_X1 U22127 ( .B1(n21246), .B2(n25121), .C1(n19582), .C2(n25115), .A(
        n23226), .ZN(n23221) );
  AOI22_X1 U22128 ( .A1(n25109), .A2(n24893), .B1(n25103), .B2(n20029), .ZN(
        n23226) );
  OAI221_X1 U22129 ( .B1(n21182), .B2(n25067), .C1(n20158), .C2(n25061), .A(
        n23232), .ZN(n23231) );
  AOI22_X1 U22130 ( .A1(n25055), .A2(n24165), .B1(n25048), .B2(OUT2[39]), .ZN(
        n23232) );
  OAI221_X1 U22131 ( .B1(n21245), .B2(n25121), .C1(n19581), .C2(n25115), .A(
        n23208), .ZN(n23203) );
  AOI22_X1 U22132 ( .A1(n25109), .A2(n24894), .B1(n25103), .B2(n20028), .ZN(
        n23208) );
  OAI221_X1 U22133 ( .B1(n21181), .B2(n25067), .C1(n20157), .C2(n25061), .A(
        n23214), .ZN(n23213) );
  AOI22_X1 U22134 ( .A1(n25055), .A2(n24167), .B1(n25048), .B2(OUT2[40]), .ZN(
        n23214) );
  OAI221_X1 U22135 ( .B1(n21244), .B2(n25121), .C1(n19580), .C2(n25115), .A(
        n23190), .ZN(n23185) );
  AOI22_X1 U22136 ( .A1(n25109), .A2(n24895), .B1(n25103), .B2(n20027), .ZN(
        n23190) );
  OAI221_X1 U22137 ( .B1(n21180), .B2(n25067), .C1(n20156), .C2(n25061), .A(
        n23196), .ZN(n23195) );
  AOI22_X1 U22138 ( .A1(n25055), .A2(n24169), .B1(n25048), .B2(OUT2[41]), .ZN(
        n23196) );
  OAI221_X1 U22139 ( .B1(n21243), .B2(n25121), .C1(n19579), .C2(n25115), .A(
        n23172), .ZN(n23167) );
  AOI22_X1 U22140 ( .A1(n25109), .A2(n24896), .B1(n25103), .B2(n20026), .ZN(
        n23172) );
  OAI221_X1 U22141 ( .B1(n21179), .B2(n25067), .C1(n20155), .C2(n25061), .A(
        n23178), .ZN(n23177) );
  AOI22_X1 U22142 ( .A1(n25055), .A2(n24171), .B1(n25047), .B2(OUT2[42]), .ZN(
        n23178) );
  OAI221_X1 U22143 ( .B1(n21242), .B2(n25121), .C1(n19578), .C2(n25115), .A(
        n23154), .ZN(n23149) );
  AOI22_X1 U22144 ( .A1(n25109), .A2(n24897), .B1(n25103), .B2(n20025), .ZN(
        n23154) );
  OAI221_X1 U22145 ( .B1(n21178), .B2(n25067), .C1(n20154), .C2(n25061), .A(
        n23160), .ZN(n23159) );
  AOI22_X1 U22146 ( .A1(n25055), .A2(n24173), .B1(n25047), .B2(OUT2[43]), .ZN(
        n23160) );
  OAI221_X1 U22147 ( .B1(n21241), .B2(n25121), .C1(n19577), .C2(n25115), .A(
        n23136), .ZN(n23131) );
  AOI22_X1 U22148 ( .A1(n25109), .A2(n24898), .B1(n25103), .B2(n20024), .ZN(
        n23136) );
  OAI221_X1 U22149 ( .B1(n21177), .B2(n25067), .C1(n20153), .C2(n25061), .A(
        n23142), .ZN(n23141) );
  AOI22_X1 U22150 ( .A1(n25055), .A2(n24175), .B1(n25047), .B2(OUT2[44]), .ZN(
        n23142) );
  OAI221_X1 U22151 ( .B1(n21240), .B2(n25121), .C1(n19576), .C2(n25115), .A(
        n23118), .ZN(n23113) );
  AOI22_X1 U22152 ( .A1(n25109), .A2(n24899), .B1(n25103), .B2(n20023), .ZN(
        n23118) );
  OAI221_X1 U22153 ( .B1(n21176), .B2(n25067), .C1(n20152), .C2(n25061), .A(
        n23124), .ZN(n23123) );
  AOI22_X1 U22154 ( .A1(n25055), .A2(n24177), .B1(n25047), .B2(OUT2[45]), .ZN(
        n23124) );
  OAI221_X1 U22155 ( .B1(n21239), .B2(n25121), .C1(n19575), .C2(n25115), .A(
        n23100), .ZN(n23095) );
  AOI22_X1 U22156 ( .A1(n25109), .A2(n24900), .B1(n25103), .B2(n20022), .ZN(
        n23100) );
  OAI221_X1 U22157 ( .B1(n21175), .B2(n25067), .C1(n20151), .C2(n25061), .A(
        n23106), .ZN(n23105) );
  AOI22_X1 U22158 ( .A1(n25055), .A2(n24179), .B1(n25047), .B2(OUT2[46]), .ZN(
        n23106) );
  OAI221_X1 U22159 ( .B1(n21238), .B2(n25121), .C1(n19574), .C2(n25115), .A(
        n23082), .ZN(n23077) );
  AOI22_X1 U22160 ( .A1(n25109), .A2(n24901), .B1(n25103), .B2(n20021), .ZN(
        n23082) );
  OAI221_X1 U22161 ( .B1(n21174), .B2(n25067), .C1(n20150), .C2(n25061), .A(
        n23088), .ZN(n23087) );
  AOI22_X1 U22162 ( .A1(n25055), .A2(n24181), .B1(n25047), .B2(OUT2[47]), .ZN(
        n23088) );
  OAI221_X1 U22163 ( .B1(n21237), .B2(n25122), .C1(n19573), .C2(n25116), .A(
        n23064), .ZN(n23059) );
  AOI22_X1 U22164 ( .A1(n25110), .A2(n24902), .B1(n25104), .B2(n20020), .ZN(
        n23064) );
  OAI221_X1 U22165 ( .B1(n21173), .B2(n25068), .C1(n20149), .C2(n25062), .A(
        n23070), .ZN(n23069) );
  AOI22_X1 U22166 ( .A1(n25056), .A2(n24183), .B1(n25047), .B2(OUT2[48]), .ZN(
        n23070) );
  OAI221_X1 U22167 ( .B1(n21236), .B2(n25122), .C1(n19572), .C2(n25116), .A(
        n23046), .ZN(n23041) );
  AOI22_X1 U22168 ( .A1(n25110), .A2(n24903), .B1(n25104), .B2(n20019), .ZN(
        n23046) );
  OAI221_X1 U22169 ( .B1(n21172), .B2(n25068), .C1(n20148), .C2(n25062), .A(
        n23052), .ZN(n23051) );
  AOI22_X1 U22170 ( .A1(n25056), .A2(n24185), .B1(n25047), .B2(OUT2[49]), .ZN(
        n23052) );
  OAI221_X1 U22171 ( .B1(n21235), .B2(n25122), .C1(n19571), .C2(n25116), .A(
        n23028), .ZN(n23023) );
  AOI22_X1 U22172 ( .A1(n25110), .A2(n24904), .B1(n25104), .B2(n20018), .ZN(
        n23028) );
  OAI221_X1 U22173 ( .B1(n21171), .B2(n25068), .C1(n20147), .C2(n25062), .A(
        n23034), .ZN(n23033) );
  AOI22_X1 U22174 ( .A1(n25056), .A2(n24187), .B1(n25047), .B2(OUT2[50]), .ZN(
        n23034) );
  OAI221_X1 U22175 ( .B1(n21234), .B2(n25122), .C1(n19570), .C2(n25116), .A(
        n23010), .ZN(n23005) );
  AOI22_X1 U22176 ( .A1(n25110), .A2(n24905), .B1(n25104), .B2(n20017), .ZN(
        n23010) );
  OAI221_X1 U22177 ( .B1(n21170), .B2(n25068), .C1(n20146), .C2(n25062), .A(
        n23016), .ZN(n23015) );
  AOI22_X1 U22178 ( .A1(n25056), .A2(n24189), .B1(n25047), .B2(OUT2[51]), .ZN(
        n23016) );
  OAI221_X1 U22179 ( .B1(n21233), .B2(n25122), .C1(n19569), .C2(n25116), .A(
        n22992), .ZN(n22987) );
  AOI22_X1 U22180 ( .A1(n25110), .A2(n24906), .B1(n25104), .B2(n20016), .ZN(
        n22992) );
  OAI221_X1 U22181 ( .B1(n21169), .B2(n25068), .C1(n20145), .C2(n25062), .A(
        n22998), .ZN(n22997) );
  AOI22_X1 U22182 ( .A1(n25056), .A2(n24191), .B1(n25047), .B2(OUT2[52]), .ZN(
        n22998) );
  OAI221_X1 U22183 ( .B1(n21232), .B2(n25122), .C1(n19568), .C2(n25116), .A(
        n22974), .ZN(n22969) );
  AOI22_X1 U22184 ( .A1(n25110), .A2(n24907), .B1(n25104), .B2(n20015), .ZN(
        n22974) );
  OAI221_X1 U22185 ( .B1(n21168), .B2(n25068), .C1(n20144), .C2(n25062), .A(
        n22980), .ZN(n22979) );
  AOI22_X1 U22186 ( .A1(n25056), .A2(n24193), .B1(n25047), .B2(OUT2[53]), .ZN(
        n22980) );
  OAI221_X1 U22187 ( .B1(n21231), .B2(n25122), .C1(n19567), .C2(n25116), .A(
        n22956), .ZN(n22951) );
  AOI22_X1 U22188 ( .A1(n25110), .A2(n24908), .B1(n25104), .B2(n20014), .ZN(
        n22956) );
  OAI221_X1 U22189 ( .B1(n21167), .B2(n25068), .C1(n20143), .C2(n25062), .A(
        n22962), .ZN(n22961) );
  AOI22_X1 U22190 ( .A1(n25056), .A2(n24195), .B1(n25047), .B2(OUT2[54]), .ZN(
        n22962) );
  OAI221_X1 U22191 ( .B1(n21230), .B2(n25122), .C1(n19566), .C2(n25116), .A(
        n22938), .ZN(n22933) );
  AOI22_X1 U22192 ( .A1(n25110), .A2(n24909), .B1(n25104), .B2(n20013), .ZN(
        n22938) );
  OAI221_X1 U22193 ( .B1(n21166), .B2(n25068), .C1(n20142), .C2(n25062), .A(
        n22944), .ZN(n22943) );
  AOI22_X1 U22194 ( .A1(n25056), .A2(n24197), .B1(n25046), .B2(OUT2[55]), .ZN(
        n22944) );
  OAI221_X1 U22195 ( .B1(n21229), .B2(n25122), .C1(n19565), .C2(n25116), .A(
        n22920), .ZN(n22915) );
  AOI22_X1 U22196 ( .A1(n25110), .A2(n24910), .B1(n25104), .B2(n20012), .ZN(
        n22920) );
  OAI221_X1 U22197 ( .B1(n21165), .B2(n25068), .C1(n20141), .C2(n25062), .A(
        n22926), .ZN(n22925) );
  AOI22_X1 U22198 ( .A1(n25056), .A2(n24199), .B1(n25046), .B2(OUT2[56]), .ZN(
        n22926) );
  OAI221_X1 U22199 ( .B1(n21228), .B2(n25122), .C1(n19564), .C2(n25116), .A(
        n22902), .ZN(n22897) );
  AOI22_X1 U22200 ( .A1(n25110), .A2(n24911), .B1(n25104), .B2(n20011), .ZN(
        n22902) );
  OAI221_X1 U22201 ( .B1(n21164), .B2(n25068), .C1(n20140), .C2(n25062), .A(
        n22908), .ZN(n22907) );
  AOI22_X1 U22202 ( .A1(n25056), .A2(n24201), .B1(n25046), .B2(OUT2[57]), .ZN(
        n22908) );
  OAI221_X1 U22203 ( .B1(n21227), .B2(n25122), .C1(n19563), .C2(n25116), .A(
        n22884), .ZN(n22879) );
  AOI22_X1 U22204 ( .A1(n25110), .A2(n24912), .B1(n25104), .B2(n20010), .ZN(
        n22884) );
  OAI221_X1 U22205 ( .B1(n21163), .B2(n25068), .C1(n20139), .C2(n25062), .A(
        n22890), .ZN(n22889) );
  AOI22_X1 U22206 ( .A1(n25056), .A2(n24203), .B1(n25046), .B2(OUT2[58]), .ZN(
        n22890) );
  OAI221_X1 U22207 ( .B1(n21226), .B2(n25122), .C1(n19562), .C2(n25116), .A(
        n22866), .ZN(n22861) );
  AOI22_X1 U22208 ( .A1(n25110), .A2(n24913), .B1(n25104), .B2(n20009), .ZN(
        n22866) );
  OAI221_X1 U22209 ( .B1(n21162), .B2(n25068), .C1(n20138), .C2(n25062), .A(
        n22872), .ZN(n22871) );
  AOI22_X1 U22210 ( .A1(n25056), .A2(n24205), .B1(n25046), .B2(OUT2[59]), .ZN(
        n22872) );
  OAI221_X1 U22211 ( .B1(n21285), .B2(n25316), .C1(n19621), .C2(n25310), .A(
        n22739), .ZN(n22726) );
  AOI22_X1 U22212 ( .A1(n25304), .A2(n24854), .B1(n25298), .B2(n20068), .ZN(
        n22739) );
  OAI221_X1 U22213 ( .B1(n21221), .B2(n25262), .C1(n20197), .C2(n25256), .A(
        n22748), .ZN(n22747) );
  AOI22_X1 U22214 ( .A1(n25250), .A2(n24087), .B1(n25244), .B2(OUT1[0]), .ZN(
        n22748) );
  OAI221_X1 U22215 ( .B1(n21284), .B2(n25316), .C1(n19620), .C2(n25310), .A(
        n22713), .ZN(n22708) );
  AOI22_X1 U22216 ( .A1(n25304), .A2(n24855), .B1(n25298), .B2(n20067), .ZN(
        n22713) );
  OAI221_X1 U22217 ( .B1(n21220), .B2(n25262), .C1(n20196), .C2(n25256), .A(
        n22719), .ZN(n22718) );
  AOI22_X1 U22218 ( .A1(n25250), .A2(n24089), .B1(n25249), .B2(OUT1[1]), .ZN(
        n22719) );
  OAI221_X1 U22219 ( .B1(n21283), .B2(n25316), .C1(n19619), .C2(n25310), .A(
        n22695), .ZN(n22690) );
  AOI22_X1 U22220 ( .A1(n25304), .A2(n24856), .B1(n25298), .B2(n20066), .ZN(
        n22695) );
  OAI221_X1 U22221 ( .B1(n21219), .B2(n25262), .C1(n20195), .C2(n25256), .A(
        n22701), .ZN(n22700) );
  AOI22_X1 U22222 ( .A1(n25250), .A2(n24091), .B1(n25249), .B2(OUT1[2]), .ZN(
        n22701) );
  OAI221_X1 U22223 ( .B1(n21282), .B2(n25316), .C1(n19618), .C2(n25310), .A(
        n22677), .ZN(n22672) );
  AOI22_X1 U22224 ( .A1(n25304), .A2(n24857), .B1(n25298), .B2(n20065), .ZN(
        n22677) );
  OAI221_X1 U22225 ( .B1(n21218), .B2(n25262), .C1(n20194), .C2(n25256), .A(
        n22683), .ZN(n22682) );
  AOI22_X1 U22226 ( .A1(n25250), .A2(n24093), .B1(n25249), .B2(OUT1[3]), .ZN(
        n22683) );
  OAI221_X1 U22227 ( .B1(n21281), .B2(n25316), .C1(n19617), .C2(n25310), .A(
        n22659), .ZN(n22654) );
  AOI22_X1 U22228 ( .A1(n25304), .A2(n24858), .B1(n25298), .B2(n20064), .ZN(
        n22659) );
  OAI221_X1 U22229 ( .B1(n21217), .B2(n25262), .C1(n20193), .C2(n25256), .A(
        n22665), .ZN(n22664) );
  AOI22_X1 U22230 ( .A1(n25250), .A2(n24095), .B1(n25248), .B2(OUT1[4]), .ZN(
        n22665) );
  OAI221_X1 U22231 ( .B1(n21280), .B2(n25316), .C1(n19616), .C2(n25310), .A(
        n22641), .ZN(n22636) );
  AOI22_X1 U22232 ( .A1(n25304), .A2(n24859), .B1(n25298), .B2(n20063), .ZN(
        n22641) );
  OAI221_X1 U22233 ( .B1(n21216), .B2(n25262), .C1(n20192), .C2(n25256), .A(
        n22647), .ZN(n22646) );
  AOI22_X1 U22234 ( .A1(n25250), .A2(n24097), .B1(n25248), .B2(OUT1[5]), .ZN(
        n22647) );
  OAI221_X1 U22235 ( .B1(n21279), .B2(n25316), .C1(n19615), .C2(n25310), .A(
        n22623), .ZN(n22618) );
  AOI22_X1 U22236 ( .A1(n25304), .A2(n24860), .B1(n25298), .B2(n20062), .ZN(
        n22623) );
  OAI221_X1 U22237 ( .B1(n21215), .B2(n25262), .C1(n20191), .C2(n25256), .A(
        n22629), .ZN(n22628) );
  AOI22_X1 U22238 ( .A1(n25250), .A2(n24099), .B1(n25248), .B2(OUT1[6]), .ZN(
        n22629) );
  OAI221_X1 U22239 ( .B1(n21278), .B2(n25316), .C1(n19614), .C2(n25310), .A(
        n22605), .ZN(n22600) );
  AOI22_X1 U22240 ( .A1(n25304), .A2(n24861), .B1(n25298), .B2(n20061), .ZN(
        n22605) );
  OAI221_X1 U22241 ( .B1(n21214), .B2(n25262), .C1(n20190), .C2(n25256), .A(
        n22611), .ZN(n22610) );
  AOI22_X1 U22242 ( .A1(n25250), .A2(n24101), .B1(n25248), .B2(OUT1[7]), .ZN(
        n22611) );
  OAI221_X1 U22243 ( .B1(n21277), .B2(n25316), .C1(n19613), .C2(n25310), .A(
        n22587), .ZN(n22582) );
  AOI22_X1 U22244 ( .A1(n25304), .A2(n24862), .B1(n25298), .B2(n20060), .ZN(
        n22587) );
  OAI221_X1 U22245 ( .B1(n21213), .B2(n25262), .C1(n20189), .C2(n25256), .A(
        n22593), .ZN(n22592) );
  AOI22_X1 U22246 ( .A1(n25250), .A2(n24103), .B1(n25248), .B2(OUT1[8]), .ZN(
        n22593) );
  OAI221_X1 U22247 ( .B1(n21276), .B2(n25316), .C1(n19612), .C2(n25310), .A(
        n22569), .ZN(n22564) );
  AOI22_X1 U22248 ( .A1(n25304), .A2(n24863), .B1(n25298), .B2(n20059), .ZN(
        n22569) );
  OAI221_X1 U22249 ( .B1(n21212), .B2(n25262), .C1(n20188), .C2(n25256), .A(
        n22575), .ZN(n22574) );
  AOI22_X1 U22250 ( .A1(n25250), .A2(n24105), .B1(n25248), .B2(OUT1[9]), .ZN(
        n22575) );
  OAI221_X1 U22251 ( .B1(n21275), .B2(n25316), .C1(n19611), .C2(n25310), .A(
        n22551), .ZN(n22546) );
  AOI22_X1 U22252 ( .A1(n25304), .A2(n24864), .B1(n25298), .B2(n20058), .ZN(
        n22551) );
  OAI221_X1 U22253 ( .B1(n21211), .B2(n25262), .C1(n20187), .C2(n25256), .A(
        n22557), .ZN(n22556) );
  AOI22_X1 U22254 ( .A1(n25250), .A2(n24107), .B1(n25248), .B2(OUT1[10]), .ZN(
        n22557) );
  OAI221_X1 U22255 ( .B1(n21274), .B2(n25316), .C1(n19610), .C2(n25310), .A(
        n22533), .ZN(n22528) );
  AOI22_X1 U22256 ( .A1(n25304), .A2(n24865), .B1(n25298), .B2(n20057), .ZN(
        n22533) );
  OAI221_X1 U22257 ( .B1(n21210), .B2(n25262), .C1(n20186), .C2(n25256), .A(
        n22539), .ZN(n22538) );
  AOI22_X1 U22258 ( .A1(n25250), .A2(n24109), .B1(n25248), .B2(OUT1[11]), .ZN(
        n22539) );
  OAI221_X1 U22259 ( .B1(n21273), .B2(n25317), .C1(n19609), .C2(n25311), .A(
        n22515), .ZN(n22510) );
  AOI22_X1 U22260 ( .A1(n25305), .A2(n24866), .B1(n25299), .B2(n20056), .ZN(
        n22515) );
  OAI221_X1 U22261 ( .B1(n21209), .B2(n25263), .C1(n20185), .C2(n25257), .A(
        n22521), .ZN(n22520) );
  AOI22_X1 U22262 ( .A1(n25251), .A2(n24111), .B1(n25248), .B2(OUT1[12]), .ZN(
        n22521) );
  OAI221_X1 U22263 ( .B1(n21272), .B2(n25317), .C1(n19608), .C2(n25311), .A(
        n22497), .ZN(n22492) );
  AOI22_X1 U22264 ( .A1(n25305), .A2(n24867), .B1(n25299), .B2(n20055), .ZN(
        n22497) );
  OAI221_X1 U22265 ( .B1(n21208), .B2(n25263), .C1(n20184), .C2(n25257), .A(
        n22503), .ZN(n22502) );
  AOI22_X1 U22266 ( .A1(n25251), .A2(n24113), .B1(n25248), .B2(OUT1[13]), .ZN(
        n22503) );
  OAI221_X1 U22267 ( .B1(n21271), .B2(n25317), .C1(n19607), .C2(n25311), .A(
        n22479), .ZN(n22474) );
  AOI22_X1 U22268 ( .A1(n25305), .A2(n24868), .B1(n25299), .B2(n20054), .ZN(
        n22479) );
  OAI221_X1 U22269 ( .B1(n21207), .B2(n25263), .C1(n20183), .C2(n25257), .A(
        n22485), .ZN(n22484) );
  AOI22_X1 U22270 ( .A1(n25251), .A2(n24115), .B1(n25248), .B2(OUT1[14]), .ZN(
        n22485) );
  OAI221_X1 U22271 ( .B1(n21270), .B2(n25317), .C1(n19606), .C2(n25311), .A(
        n22461), .ZN(n22456) );
  AOI22_X1 U22272 ( .A1(n25305), .A2(n24869), .B1(n25299), .B2(n20053), .ZN(
        n22461) );
  OAI221_X1 U22273 ( .B1(n21206), .B2(n25263), .C1(n20182), .C2(n25257), .A(
        n22467), .ZN(n22466) );
  AOI22_X1 U22274 ( .A1(n25251), .A2(n24117), .B1(n25248), .B2(OUT1[15]), .ZN(
        n22467) );
  OAI221_X1 U22275 ( .B1(n21269), .B2(n25317), .C1(n19605), .C2(n25311), .A(
        n22443), .ZN(n22438) );
  AOI22_X1 U22276 ( .A1(n25305), .A2(n24870), .B1(n25299), .B2(n20052), .ZN(
        n22443) );
  OAI221_X1 U22277 ( .B1(n21205), .B2(n25263), .C1(n20181), .C2(n25257), .A(
        n22449), .ZN(n22448) );
  AOI22_X1 U22278 ( .A1(n25251), .A2(n24119), .B1(n25248), .B2(OUT1[16]), .ZN(
        n22449) );
  OAI221_X1 U22279 ( .B1(n21268), .B2(n25317), .C1(n19604), .C2(n25311), .A(
        n22425), .ZN(n22420) );
  AOI22_X1 U22280 ( .A1(n25305), .A2(n24871), .B1(n25299), .B2(n20051), .ZN(
        n22425) );
  OAI221_X1 U22281 ( .B1(n21204), .B2(n25263), .C1(n20180), .C2(n25257), .A(
        n22431), .ZN(n22430) );
  AOI22_X1 U22282 ( .A1(n25251), .A2(n24121), .B1(n25247), .B2(OUT1[17]), .ZN(
        n22431) );
  OAI221_X1 U22283 ( .B1(n21267), .B2(n25317), .C1(n19603), .C2(n25311), .A(
        n22407), .ZN(n22402) );
  AOI22_X1 U22284 ( .A1(n25305), .A2(n24872), .B1(n25299), .B2(n20050), .ZN(
        n22407) );
  OAI221_X1 U22285 ( .B1(n21203), .B2(n25263), .C1(n20179), .C2(n25257), .A(
        n22413), .ZN(n22412) );
  AOI22_X1 U22286 ( .A1(n25251), .A2(n24123), .B1(n25247), .B2(OUT1[18]), .ZN(
        n22413) );
  OAI221_X1 U22287 ( .B1(n21266), .B2(n25317), .C1(n19602), .C2(n25311), .A(
        n22389), .ZN(n22384) );
  AOI22_X1 U22288 ( .A1(n25305), .A2(n24873), .B1(n25299), .B2(n20049), .ZN(
        n22389) );
  OAI221_X1 U22289 ( .B1(n21202), .B2(n25263), .C1(n20178), .C2(n25257), .A(
        n22395), .ZN(n22394) );
  AOI22_X1 U22290 ( .A1(n25251), .A2(n24125), .B1(n25247), .B2(OUT1[19]), .ZN(
        n22395) );
  OAI221_X1 U22291 ( .B1(n21265), .B2(n25317), .C1(n19601), .C2(n25311), .A(
        n22371), .ZN(n22366) );
  AOI22_X1 U22292 ( .A1(n25305), .A2(n24874), .B1(n25299), .B2(n20048), .ZN(
        n22371) );
  OAI221_X1 U22293 ( .B1(n21201), .B2(n25263), .C1(n20177), .C2(n25257), .A(
        n22377), .ZN(n22376) );
  AOI22_X1 U22294 ( .A1(n25251), .A2(n24127), .B1(n25247), .B2(OUT1[20]), .ZN(
        n22377) );
  OAI221_X1 U22295 ( .B1(n21264), .B2(n25317), .C1(n19600), .C2(n25311), .A(
        n22353), .ZN(n22348) );
  AOI22_X1 U22296 ( .A1(n25305), .A2(n24875), .B1(n25299), .B2(n20047), .ZN(
        n22353) );
  OAI221_X1 U22297 ( .B1(n21200), .B2(n25263), .C1(n20176), .C2(n25257), .A(
        n22359), .ZN(n22358) );
  AOI22_X1 U22298 ( .A1(n25251), .A2(n24129), .B1(n25247), .B2(OUT1[21]), .ZN(
        n22359) );
  OAI221_X1 U22299 ( .B1(n21263), .B2(n25317), .C1(n19599), .C2(n25311), .A(
        n22335), .ZN(n22330) );
  AOI22_X1 U22300 ( .A1(n25305), .A2(n24876), .B1(n25299), .B2(n20046), .ZN(
        n22335) );
  OAI221_X1 U22301 ( .B1(n21199), .B2(n25263), .C1(n20175), .C2(n25257), .A(
        n22341), .ZN(n22340) );
  AOI22_X1 U22302 ( .A1(n25251), .A2(n24131), .B1(n25247), .B2(OUT1[22]), .ZN(
        n22341) );
  OAI221_X1 U22303 ( .B1(n21262), .B2(n25317), .C1(n19598), .C2(n25311), .A(
        n22317), .ZN(n22312) );
  AOI22_X1 U22304 ( .A1(n25305), .A2(n24877), .B1(n25299), .B2(n20045), .ZN(
        n22317) );
  OAI221_X1 U22305 ( .B1(n21198), .B2(n25263), .C1(n20174), .C2(n25257), .A(
        n22323), .ZN(n22322) );
  AOI22_X1 U22306 ( .A1(n25251), .A2(n24133), .B1(n25247), .B2(OUT1[23]), .ZN(
        n22323) );
  OAI221_X1 U22307 ( .B1(n21261), .B2(n25318), .C1(n19597), .C2(n25312), .A(
        n22299), .ZN(n22294) );
  AOI22_X1 U22308 ( .A1(n25306), .A2(n24878), .B1(n25300), .B2(n20044), .ZN(
        n22299) );
  OAI221_X1 U22309 ( .B1(n21197), .B2(n25264), .C1(n20173), .C2(n25258), .A(
        n22305), .ZN(n22304) );
  AOI22_X1 U22310 ( .A1(n25252), .A2(n24135), .B1(n25247), .B2(OUT1[24]), .ZN(
        n22305) );
  OAI221_X1 U22311 ( .B1(n21260), .B2(n25318), .C1(n19596), .C2(n25312), .A(
        n22281), .ZN(n22276) );
  AOI22_X1 U22312 ( .A1(n25306), .A2(n24879), .B1(n25300), .B2(n20043), .ZN(
        n22281) );
  OAI221_X1 U22313 ( .B1(n21196), .B2(n25264), .C1(n20172), .C2(n25258), .A(
        n22287), .ZN(n22286) );
  AOI22_X1 U22314 ( .A1(n25252), .A2(n24137), .B1(n25247), .B2(OUT1[25]), .ZN(
        n22287) );
  OAI221_X1 U22315 ( .B1(n21259), .B2(n25318), .C1(n19595), .C2(n25312), .A(
        n22263), .ZN(n22258) );
  AOI22_X1 U22316 ( .A1(n25306), .A2(n24880), .B1(n25300), .B2(n20042), .ZN(
        n22263) );
  OAI221_X1 U22317 ( .B1(n21195), .B2(n25264), .C1(n20171), .C2(n25258), .A(
        n22269), .ZN(n22268) );
  AOI22_X1 U22318 ( .A1(n25252), .A2(n24139), .B1(n25247), .B2(OUT1[26]), .ZN(
        n22269) );
  OAI221_X1 U22319 ( .B1(n21258), .B2(n25318), .C1(n19594), .C2(n25312), .A(
        n22245), .ZN(n22240) );
  AOI22_X1 U22320 ( .A1(n25306), .A2(n24881), .B1(n25300), .B2(n20041), .ZN(
        n22245) );
  OAI221_X1 U22321 ( .B1(n21194), .B2(n25264), .C1(n20170), .C2(n25258), .A(
        n22251), .ZN(n22250) );
  AOI22_X1 U22322 ( .A1(n25252), .A2(n24141), .B1(n25247), .B2(OUT1[27]), .ZN(
        n22251) );
  OAI221_X1 U22323 ( .B1(n21257), .B2(n25318), .C1(n19593), .C2(n25312), .A(
        n22227), .ZN(n22222) );
  AOI22_X1 U22324 ( .A1(n25306), .A2(n24882), .B1(n25300), .B2(n20040), .ZN(
        n22227) );
  OAI221_X1 U22325 ( .B1(n21193), .B2(n25264), .C1(n20169), .C2(n25258), .A(
        n22233), .ZN(n22232) );
  AOI22_X1 U22326 ( .A1(n25252), .A2(n24143), .B1(n25247), .B2(OUT1[28]), .ZN(
        n22233) );
  OAI221_X1 U22327 ( .B1(n21256), .B2(n25318), .C1(n19592), .C2(n25312), .A(
        n22209), .ZN(n22204) );
  AOI22_X1 U22328 ( .A1(n25306), .A2(n24883), .B1(n25300), .B2(n20039), .ZN(
        n22209) );
  OAI221_X1 U22329 ( .B1(n21192), .B2(n25264), .C1(n20168), .C2(n25258), .A(
        n22215), .ZN(n22214) );
  AOI22_X1 U22330 ( .A1(n25252), .A2(n24145), .B1(n25247), .B2(OUT1[29]), .ZN(
        n22215) );
  OAI221_X1 U22331 ( .B1(n21255), .B2(n25318), .C1(n19591), .C2(n25312), .A(
        n22191), .ZN(n22186) );
  AOI22_X1 U22332 ( .A1(n25306), .A2(n24884), .B1(n25300), .B2(n20038), .ZN(
        n22191) );
  OAI221_X1 U22333 ( .B1(n21191), .B2(n25264), .C1(n20167), .C2(n25258), .A(
        n22197), .ZN(n22196) );
  AOI22_X1 U22334 ( .A1(n25252), .A2(n24147), .B1(n25246), .B2(OUT1[30]), .ZN(
        n22197) );
  OAI221_X1 U22335 ( .B1(n21254), .B2(n25318), .C1(n19590), .C2(n25312), .A(
        n22173), .ZN(n22168) );
  AOI22_X1 U22336 ( .A1(n25306), .A2(n24885), .B1(n25300), .B2(n20037), .ZN(
        n22173) );
  OAI221_X1 U22337 ( .B1(n21190), .B2(n25264), .C1(n20166), .C2(n25258), .A(
        n22179), .ZN(n22178) );
  AOI22_X1 U22338 ( .A1(n25252), .A2(n24149), .B1(n25246), .B2(OUT1[31]), .ZN(
        n22179) );
  OAI221_X1 U22339 ( .B1(n21253), .B2(n25318), .C1(n19589), .C2(n25312), .A(
        n22155), .ZN(n22150) );
  AOI22_X1 U22340 ( .A1(n25306), .A2(n24886), .B1(n25300), .B2(n20036), .ZN(
        n22155) );
  OAI221_X1 U22341 ( .B1(n21189), .B2(n25264), .C1(n20165), .C2(n25258), .A(
        n22161), .ZN(n22160) );
  AOI22_X1 U22342 ( .A1(n25252), .A2(n24151), .B1(n25246), .B2(OUT1[32]), .ZN(
        n22161) );
  OAI221_X1 U22343 ( .B1(n21252), .B2(n25318), .C1(n19588), .C2(n25312), .A(
        n22137), .ZN(n22132) );
  AOI22_X1 U22344 ( .A1(n25306), .A2(n24887), .B1(n25300), .B2(n20035), .ZN(
        n22137) );
  OAI221_X1 U22345 ( .B1(n21188), .B2(n25264), .C1(n20164), .C2(n25258), .A(
        n22143), .ZN(n22142) );
  AOI22_X1 U22346 ( .A1(n25252), .A2(n24153), .B1(n25246), .B2(OUT1[33]), .ZN(
        n22143) );
  OAI221_X1 U22347 ( .B1(n21251), .B2(n25318), .C1(n19587), .C2(n25312), .A(
        n22119), .ZN(n22114) );
  AOI22_X1 U22348 ( .A1(n25306), .A2(n24888), .B1(n25300), .B2(n20034), .ZN(
        n22119) );
  OAI221_X1 U22349 ( .B1(n21187), .B2(n25264), .C1(n20163), .C2(n25258), .A(
        n22125), .ZN(n22124) );
  AOI22_X1 U22350 ( .A1(n25252), .A2(n24155), .B1(n25246), .B2(OUT1[34]), .ZN(
        n22125) );
  OAI221_X1 U22351 ( .B1(n21250), .B2(n25318), .C1(n19586), .C2(n25312), .A(
        n22101), .ZN(n22096) );
  AOI22_X1 U22352 ( .A1(n25306), .A2(n24889), .B1(n25300), .B2(n20033), .ZN(
        n22101) );
  OAI221_X1 U22353 ( .B1(n21186), .B2(n25264), .C1(n20162), .C2(n25258), .A(
        n22107), .ZN(n22106) );
  AOI22_X1 U22354 ( .A1(n25252), .A2(n24157), .B1(n25246), .B2(OUT1[35]), .ZN(
        n22107) );
  OAI221_X1 U22355 ( .B1(n21249), .B2(n25319), .C1(n19585), .C2(n25313), .A(
        n22083), .ZN(n22078) );
  AOI22_X1 U22356 ( .A1(n25307), .A2(n24890), .B1(n25301), .B2(n20032), .ZN(
        n22083) );
  OAI221_X1 U22357 ( .B1(n21185), .B2(n25265), .C1(n20161), .C2(n25259), .A(
        n22089), .ZN(n22088) );
  AOI22_X1 U22358 ( .A1(n25253), .A2(n24159), .B1(n25246), .B2(OUT1[36]), .ZN(
        n22089) );
  OAI221_X1 U22359 ( .B1(n21248), .B2(n25319), .C1(n19584), .C2(n25313), .A(
        n22065), .ZN(n22060) );
  AOI22_X1 U22360 ( .A1(n25307), .A2(n24891), .B1(n25301), .B2(n20031), .ZN(
        n22065) );
  OAI221_X1 U22361 ( .B1(n21184), .B2(n25265), .C1(n20160), .C2(n25259), .A(
        n22071), .ZN(n22070) );
  AOI22_X1 U22362 ( .A1(n25253), .A2(n24161), .B1(n25246), .B2(OUT1[37]), .ZN(
        n22071) );
  OAI221_X1 U22363 ( .B1(n21247), .B2(n25319), .C1(n19583), .C2(n25313), .A(
        n22047), .ZN(n22042) );
  AOI22_X1 U22364 ( .A1(n25307), .A2(n24892), .B1(n25301), .B2(n20030), .ZN(
        n22047) );
  OAI221_X1 U22365 ( .B1(n21183), .B2(n25265), .C1(n20159), .C2(n25259), .A(
        n22053), .ZN(n22052) );
  AOI22_X1 U22366 ( .A1(n25253), .A2(n24163), .B1(n25246), .B2(OUT1[38]), .ZN(
        n22053) );
  OAI221_X1 U22367 ( .B1(n21246), .B2(n25319), .C1(n19582), .C2(n25313), .A(
        n22029), .ZN(n22024) );
  AOI22_X1 U22368 ( .A1(n25307), .A2(n24893), .B1(n25301), .B2(n20029), .ZN(
        n22029) );
  OAI221_X1 U22369 ( .B1(n21182), .B2(n25265), .C1(n20158), .C2(n25259), .A(
        n22035), .ZN(n22034) );
  AOI22_X1 U22370 ( .A1(n25253), .A2(n24165), .B1(n25246), .B2(OUT1[39]), .ZN(
        n22035) );
  OAI221_X1 U22371 ( .B1(n21245), .B2(n25319), .C1(n19581), .C2(n25313), .A(
        n22011), .ZN(n22006) );
  AOI22_X1 U22372 ( .A1(n25307), .A2(n24894), .B1(n25301), .B2(n20028), .ZN(
        n22011) );
  OAI221_X1 U22373 ( .B1(n21181), .B2(n25265), .C1(n20157), .C2(n25259), .A(
        n22017), .ZN(n22016) );
  AOI22_X1 U22374 ( .A1(n25253), .A2(n24167), .B1(n25246), .B2(OUT1[40]), .ZN(
        n22017) );
  OAI221_X1 U22375 ( .B1(n21244), .B2(n25319), .C1(n19580), .C2(n25313), .A(
        n21993), .ZN(n21988) );
  AOI22_X1 U22376 ( .A1(n25307), .A2(n24895), .B1(n25301), .B2(n20027), .ZN(
        n21993) );
  OAI221_X1 U22377 ( .B1(n21180), .B2(n25265), .C1(n20156), .C2(n25259), .A(
        n21999), .ZN(n21998) );
  AOI22_X1 U22378 ( .A1(n25253), .A2(n24169), .B1(n25246), .B2(OUT1[41]), .ZN(
        n21999) );
  OAI221_X1 U22379 ( .B1(n21243), .B2(n25319), .C1(n19579), .C2(n25313), .A(
        n21975), .ZN(n21970) );
  AOI22_X1 U22380 ( .A1(n25307), .A2(n24896), .B1(n25301), .B2(n20026), .ZN(
        n21975) );
  OAI221_X1 U22381 ( .B1(n21179), .B2(n25265), .C1(n20155), .C2(n25259), .A(
        n21981), .ZN(n21980) );
  AOI22_X1 U22382 ( .A1(n25253), .A2(n24171), .B1(n25245), .B2(OUT1[42]), .ZN(
        n21981) );
  OAI221_X1 U22383 ( .B1(n21242), .B2(n25319), .C1(n19578), .C2(n25313), .A(
        n21957), .ZN(n21952) );
  AOI22_X1 U22384 ( .A1(n25307), .A2(n24897), .B1(n25301), .B2(n20025), .ZN(
        n21957) );
  OAI221_X1 U22385 ( .B1(n21178), .B2(n25265), .C1(n20154), .C2(n25259), .A(
        n21963), .ZN(n21962) );
  AOI22_X1 U22386 ( .A1(n25253), .A2(n24173), .B1(n25245), .B2(OUT1[43]), .ZN(
        n21963) );
  OAI221_X1 U22387 ( .B1(n21241), .B2(n25319), .C1(n19577), .C2(n25313), .A(
        n21939), .ZN(n21934) );
  AOI22_X1 U22388 ( .A1(n25307), .A2(n24898), .B1(n25301), .B2(n20024), .ZN(
        n21939) );
  OAI221_X1 U22389 ( .B1(n21177), .B2(n25265), .C1(n20153), .C2(n25259), .A(
        n21945), .ZN(n21944) );
  AOI22_X1 U22390 ( .A1(n25253), .A2(n24175), .B1(n25245), .B2(OUT1[44]), .ZN(
        n21945) );
  OAI221_X1 U22391 ( .B1(n21240), .B2(n25319), .C1(n19576), .C2(n25313), .A(
        n21921), .ZN(n21916) );
  AOI22_X1 U22392 ( .A1(n25307), .A2(n24899), .B1(n25301), .B2(n20023), .ZN(
        n21921) );
  OAI221_X1 U22393 ( .B1(n21176), .B2(n25265), .C1(n20152), .C2(n25259), .A(
        n21927), .ZN(n21926) );
  AOI22_X1 U22394 ( .A1(n25253), .A2(n24177), .B1(n25245), .B2(OUT1[45]), .ZN(
        n21927) );
  OAI221_X1 U22395 ( .B1(n21239), .B2(n25319), .C1(n19575), .C2(n25313), .A(
        n21903), .ZN(n21898) );
  AOI22_X1 U22396 ( .A1(n25307), .A2(n24900), .B1(n25301), .B2(n20022), .ZN(
        n21903) );
  OAI221_X1 U22397 ( .B1(n21175), .B2(n25265), .C1(n20151), .C2(n25259), .A(
        n21909), .ZN(n21908) );
  AOI22_X1 U22398 ( .A1(n25253), .A2(n24179), .B1(n25245), .B2(OUT1[46]), .ZN(
        n21909) );
  OAI221_X1 U22399 ( .B1(n21238), .B2(n25319), .C1(n19574), .C2(n25313), .A(
        n21885), .ZN(n21880) );
  AOI22_X1 U22400 ( .A1(n25307), .A2(n24901), .B1(n25301), .B2(n20021), .ZN(
        n21885) );
  OAI221_X1 U22401 ( .B1(n21174), .B2(n25265), .C1(n20150), .C2(n25259), .A(
        n21891), .ZN(n21890) );
  AOI22_X1 U22402 ( .A1(n25253), .A2(n24181), .B1(n25245), .B2(OUT1[47]), .ZN(
        n21891) );
  OAI221_X1 U22403 ( .B1(n21237), .B2(n25320), .C1(n19573), .C2(n25314), .A(
        n21867), .ZN(n21862) );
  AOI22_X1 U22404 ( .A1(n25308), .A2(n24902), .B1(n25302), .B2(n20020), .ZN(
        n21867) );
  OAI221_X1 U22405 ( .B1(n21173), .B2(n25266), .C1(n20149), .C2(n25260), .A(
        n21873), .ZN(n21872) );
  AOI22_X1 U22406 ( .A1(n25254), .A2(n24183), .B1(n25245), .B2(OUT1[48]), .ZN(
        n21873) );
  OAI221_X1 U22407 ( .B1(n21236), .B2(n25320), .C1(n19572), .C2(n25314), .A(
        n21849), .ZN(n21844) );
  AOI22_X1 U22408 ( .A1(n25308), .A2(n24903), .B1(n25302), .B2(n20019), .ZN(
        n21849) );
  OAI221_X1 U22409 ( .B1(n21172), .B2(n25266), .C1(n20148), .C2(n25260), .A(
        n21855), .ZN(n21854) );
  AOI22_X1 U22410 ( .A1(n25254), .A2(n24185), .B1(n25245), .B2(OUT1[49]), .ZN(
        n21855) );
  OAI221_X1 U22411 ( .B1(n21235), .B2(n25320), .C1(n19571), .C2(n25314), .A(
        n21831), .ZN(n21826) );
  AOI22_X1 U22412 ( .A1(n25308), .A2(n24904), .B1(n25302), .B2(n20018), .ZN(
        n21831) );
  OAI221_X1 U22413 ( .B1(n21171), .B2(n25266), .C1(n20147), .C2(n25260), .A(
        n21837), .ZN(n21836) );
  AOI22_X1 U22414 ( .A1(n25254), .A2(n24187), .B1(n25245), .B2(OUT1[50]), .ZN(
        n21837) );
  OAI221_X1 U22415 ( .B1(n21234), .B2(n25320), .C1(n19570), .C2(n25314), .A(
        n21813), .ZN(n21808) );
  AOI22_X1 U22416 ( .A1(n25308), .A2(n24905), .B1(n25302), .B2(n20017), .ZN(
        n21813) );
  OAI221_X1 U22417 ( .B1(n21170), .B2(n25266), .C1(n20146), .C2(n25260), .A(
        n21819), .ZN(n21818) );
  AOI22_X1 U22418 ( .A1(n25254), .A2(n24189), .B1(n25245), .B2(OUT1[51]), .ZN(
        n21819) );
  OAI221_X1 U22419 ( .B1(n21233), .B2(n25320), .C1(n19569), .C2(n25314), .A(
        n21795), .ZN(n21790) );
  AOI22_X1 U22420 ( .A1(n25308), .A2(n24906), .B1(n25302), .B2(n20016), .ZN(
        n21795) );
  OAI221_X1 U22421 ( .B1(n21169), .B2(n25266), .C1(n20145), .C2(n25260), .A(
        n21801), .ZN(n21800) );
  AOI22_X1 U22422 ( .A1(n25254), .A2(n24191), .B1(n25245), .B2(OUT1[52]), .ZN(
        n21801) );
  OAI221_X1 U22423 ( .B1(n21232), .B2(n25320), .C1(n19568), .C2(n25314), .A(
        n21777), .ZN(n21772) );
  AOI22_X1 U22424 ( .A1(n25308), .A2(n24907), .B1(n25302), .B2(n20015), .ZN(
        n21777) );
  OAI221_X1 U22425 ( .B1(n21168), .B2(n25266), .C1(n20144), .C2(n25260), .A(
        n21783), .ZN(n21782) );
  AOI22_X1 U22426 ( .A1(n25254), .A2(n24193), .B1(n25245), .B2(OUT1[53]), .ZN(
        n21783) );
  OAI221_X1 U22427 ( .B1(n21231), .B2(n25320), .C1(n19567), .C2(n25314), .A(
        n21759), .ZN(n21754) );
  AOI22_X1 U22428 ( .A1(n25308), .A2(n24908), .B1(n25302), .B2(n20014), .ZN(
        n21759) );
  OAI221_X1 U22429 ( .B1(n21167), .B2(n25266), .C1(n20143), .C2(n25260), .A(
        n21765), .ZN(n21764) );
  AOI22_X1 U22430 ( .A1(n25254), .A2(n24195), .B1(n25245), .B2(OUT1[54]), .ZN(
        n21765) );
  OAI221_X1 U22431 ( .B1(n21230), .B2(n25320), .C1(n19566), .C2(n25314), .A(
        n21741), .ZN(n21736) );
  AOI22_X1 U22432 ( .A1(n25308), .A2(n24909), .B1(n25302), .B2(n20013), .ZN(
        n21741) );
  OAI221_X1 U22433 ( .B1(n21166), .B2(n25266), .C1(n20142), .C2(n25260), .A(
        n21747), .ZN(n21746) );
  AOI22_X1 U22434 ( .A1(n25254), .A2(n24197), .B1(n25244), .B2(OUT1[55]), .ZN(
        n21747) );
  OAI221_X1 U22435 ( .B1(n21229), .B2(n25320), .C1(n19565), .C2(n25314), .A(
        n21723), .ZN(n21718) );
  AOI22_X1 U22436 ( .A1(n25308), .A2(n24910), .B1(n25302), .B2(n20012), .ZN(
        n21723) );
  OAI221_X1 U22437 ( .B1(n21165), .B2(n25266), .C1(n20141), .C2(n25260), .A(
        n21729), .ZN(n21728) );
  AOI22_X1 U22438 ( .A1(n25254), .A2(n24199), .B1(n25244), .B2(OUT1[56]), .ZN(
        n21729) );
  OAI221_X1 U22439 ( .B1(n21228), .B2(n25320), .C1(n19564), .C2(n25314), .A(
        n21705), .ZN(n21700) );
  AOI22_X1 U22440 ( .A1(n25308), .A2(n24911), .B1(n25302), .B2(n20011), .ZN(
        n21705) );
  OAI221_X1 U22441 ( .B1(n21164), .B2(n25266), .C1(n20140), .C2(n25260), .A(
        n21711), .ZN(n21710) );
  AOI22_X1 U22442 ( .A1(n25254), .A2(n24201), .B1(n25244), .B2(OUT1[57]), .ZN(
        n21711) );
  OAI221_X1 U22443 ( .B1(n21227), .B2(n25320), .C1(n19563), .C2(n25314), .A(
        n21687), .ZN(n21682) );
  AOI22_X1 U22444 ( .A1(n25308), .A2(n24912), .B1(n25302), .B2(n20010), .ZN(
        n21687) );
  OAI221_X1 U22445 ( .B1(n21163), .B2(n25266), .C1(n20139), .C2(n25260), .A(
        n21693), .ZN(n21692) );
  AOI22_X1 U22446 ( .A1(n25254), .A2(n24203), .B1(n25244), .B2(OUT1[58]), .ZN(
        n21693) );
  OAI221_X1 U22447 ( .B1(n21226), .B2(n25320), .C1(n19562), .C2(n25314), .A(
        n21669), .ZN(n21664) );
  AOI22_X1 U22448 ( .A1(n25308), .A2(n24913), .B1(n25302), .B2(n20009), .ZN(
        n21669) );
  OAI221_X1 U22449 ( .B1(n21162), .B2(n25266), .C1(n20138), .C2(n25260), .A(
        n21675), .ZN(n21674) );
  AOI22_X1 U22450 ( .A1(n25254), .A2(n24205), .B1(n25244), .B2(OUT1[59]), .ZN(
        n21675) );
  OAI22_X1 U22451 ( .A1(n25456), .A2(n20901), .B1(n25783), .B2(n25448), .ZN(
        n5823) );
  OAI22_X1 U22452 ( .A1(n25456), .A2(n20900), .B1(n25786), .B2(n25448), .ZN(
        n5824) );
  OAI22_X1 U22453 ( .A1(n25456), .A2(n20899), .B1(n25789), .B2(n25448), .ZN(
        n5825) );
  OAI22_X1 U22454 ( .A1(n25456), .A2(n20898), .B1(n25792), .B2(n25448), .ZN(
        n5826) );
  OAI22_X1 U22455 ( .A1(n25456), .A2(n20897), .B1(n25795), .B2(n25448), .ZN(
        n5827) );
  OAI22_X1 U22456 ( .A1(n25456), .A2(n20896), .B1(n25798), .B2(n25448), .ZN(
        n5828) );
  OAI22_X1 U22457 ( .A1(n25456), .A2(n20895), .B1(n25801), .B2(n25448), .ZN(
        n5829) );
  OAI22_X1 U22458 ( .A1(n25456), .A2(n20894), .B1(n25804), .B2(n25448), .ZN(
        n5830) );
  OAI22_X1 U22459 ( .A1(n25456), .A2(n20893), .B1(n25807), .B2(n25448), .ZN(
        n5831) );
  OAI22_X1 U22460 ( .A1(n25456), .A2(n20892), .B1(n25810), .B2(n25448), .ZN(
        n5832) );
  OAI22_X1 U22461 ( .A1(n25456), .A2(n20891), .B1(n25813), .B2(n25448), .ZN(
        n5833) );
  OAI22_X1 U22462 ( .A1(n25456), .A2(n20890), .B1(n25816), .B2(n25448), .ZN(
        n5834) );
  OAI22_X1 U22463 ( .A1(n25457), .A2(n20889), .B1(n25819), .B2(n25449), .ZN(
        n5835) );
  OAI22_X1 U22464 ( .A1(n25457), .A2(n20888), .B1(n25822), .B2(n25449), .ZN(
        n5836) );
  OAI22_X1 U22465 ( .A1(n25457), .A2(n20887), .B1(n25825), .B2(n25449), .ZN(
        n5837) );
  OAI22_X1 U22466 ( .A1(n25457), .A2(n20886), .B1(n25828), .B2(n25449), .ZN(
        n5838) );
  OAI22_X1 U22467 ( .A1(n25457), .A2(n20885), .B1(n25831), .B2(n25449), .ZN(
        n5839) );
  OAI22_X1 U22468 ( .A1(n25457), .A2(n20884), .B1(n25834), .B2(n25449), .ZN(
        n5840) );
  OAI22_X1 U22469 ( .A1(n25457), .A2(n20883), .B1(n25837), .B2(n25449), .ZN(
        n5841) );
  OAI22_X1 U22470 ( .A1(n25457), .A2(n20882), .B1(n25840), .B2(n25449), .ZN(
        n5842) );
  OAI22_X1 U22471 ( .A1(n25457), .A2(n20881), .B1(n25843), .B2(n25449), .ZN(
        n5843) );
  OAI22_X1 U22472 ( .A1(n25457), .A2(n20880), .B1(n25846), .B2(n25449), .ZN(
        n5844) );
  OAI22_X1 U22473 ( .A1(n25457), .A2(n20879), .B1(n25849), .B2(n25449), .ZN(
        n5845) );
  OAI22_X1 U22474 ( .A1(n25457), .A2(n20878), .B1(n25852), .B2(n25449), .ZN(
        n5846) );
  OAI22_X1 U22475 ( .A1(n25457), .A2(n20877), .B1(n25855), .B2(n25450), .ZN(
        n5847) );
  OAI22_X1 U22476 ( .A1(n25458), .A2(n20876), .B1(n25858), .B2(n25450), .ZN(
        n5848) );
  OAI22_X1 U22477 ( .A1(n25458), .A2(n20875), .B1(n25861), .B2(n25450), .ZN(
        n5849) );
  OAI22_X1 U22478 ( .A1(n25458), .A2(n20874), .B1(n25864), .B2(n25450), .ZN(
        n5850) );
  OAI22_X1 U22479 ( .A1(n25458), .A2(n20873), .B1(n25867), .B2(n25450), .ZN(
        n5851) );
  OAI22_X1 U22480 ( .A1(n25458), .A2(n20872), .B1(n25870), .B2(n25450), .ZN(
        n5852) );
  OAI22_X1 U22481 ( .A1(n25458), .A2(n20871), .B1(n25873), .B2(n25450), .ZN(
        n5853) );
  OAI22_X1 U22482 ( .A1(n25458), .A2(n20870), .B1(n25876), .B2(n25450), .ZN(
        n5854) );
  OAI22_X1 U22483 ( .A1(n25458), .A2(n20869), .B1(n25879), .B2(n25450), .ZN(
        n5855) );
  OAI22_X1 U22484 ( .A1(n25458), .A2(n20868), .B1(n25882), .B2(n25450), .ZN(
        n5856) );
  OAI22_X1 U22485 ( .A1(n25458), .A2(n20867), .B1(n25885), .B2(n25450), .ZN(
        n5857) );
  OAI22_X1 U22486 ( .A1(n25458), .A2(n20866), .B1(n25888), .B2(n25450), .ZN(
        n5858) );
  OAI22_X1 U22487 ( .A1(n25458), .A2(n20865), .B1(n25891), .B2(n25451), .ZN(
        n5859) );
  OAI22_X1 U22488 ( .A1(n25458), .A2(n20864), .B1(n25894), .B2(n25451), .ZN(
        n5860) );
  OAI22_X1 U22489 ( .A1(n25459), .A2(n20863), .B1(n25897), .B2(n25451), .ZN(
        n5861) );
  OAI22_X1 U22490 ( .A1(n25459), .A2(n20862), .B1(n25900), .B2(n25451), .ZN(
        n5862) );
  OAI22_X1 U22491 ( .A1(n25459), .A2(n20861), .B1(n25903), .B2(n25451), .ZN(
        n5863) );
  OAI22_X1 U22492 ( .A1(n25459), .A2(n20860), .B1(n25906), .B2(n25451), .ZN(
        n5864) );
  OAI22_X1 U22493 ( .A1(n25459), .A2(n20859), .B1(n25909), .B2(n25451), .ZN(
        n5865) );
  OAI22_X1 U22494 ( .A1(n25459), .A2(n20858), .B1(n25912), .B2(n25451), .ZN(
        n5866) );
  OAI22_X1 U22495 ( .A1(n25459), .A2(n20857), .B1(n25915), .B2(n25451), .ZN(
        n5867) );
  OAI22_X1 U22496 ( .A1(n25459), .A2(n20856), .B1(n25918), .B2(n25451), .ZN(
        n5868) );
  OAI22_X1 U22497 ( .A1(n25459), .A2(n20855), .B1(n25921), .B2(n25451), .ZN(
        n5869) );
  OAI22_X1 U22498 ( .A1(n25459), .A2(n20854), .B1(n25924), .B2(n25451), .ZN(
        n5870) );
  OAI22_X1 U22499 ( .A1(n25459), .A2(n20853), .B1(n25927), .B2(n25452), .ZN(
        n5871) );
  OAI22_X1 U22500 ( .A1(n25459), .A2(n20852), .B1(n25930), .B2(n25452), .ZN(
        n5872) );
  OAI22_X1 U22501 ( .A1(n25459), .A2(n20851), .B1(n25933), .B2(n25452), .ZN(
        n5873) );
  OAI22_X1 U22502 ( .A1(n25460), .A2(n20850), .B1(n25936), .B2(n25452), .ZN(
        n5874) );
  OAI22_X1 U22503 ( .A1(n25460), .A2(n20849), .B1(n25939), .B2(n25452), .ZN(
        n5875) );
  OAI22_X1 U22504 ( .A1(n25460), .A2(n20848), .B1(n25942), .B2(n25452), .ZN(
        n5876) );
  OAI22_X1 U22505 ( .A1(n25460), .A2(n20847), .B1(n25945), .B2(n25452), .ZN(
        n5877) );
  OAI22_X1 U22506 ( .A1(n25460), .A2(n20846), .B1(n25948), .B2(n25452), .ZN(
        n5878) );
  OAI22_X1 U22507 ( .A1(n25460), .A2(n20845), .B1(n25951), .B2(n25452), .ZN(
        n5879) );
  OAI22_X1 U22508 ( .A1(n25460), .A2(n20844), .B1(n25954), .B2(n25452), .ZN(
        n5880) );
  OAI22_X1 U22509 ( .A1(n25460), .A2(n20843), .B1(n25957), .B2(n25452), .ZN(
        n5881) );
  OAI22_X1 U22510 ( .A1(n25460), .A2(n20842), .B1(n25960), .B2(n25452), .ZN(
        n5882) );
  OAI22_X1 U22511 ( .A1(n25378), .A2(n20841), .B1(n25783), .B2(n25370), .ZN(
        n5439) );
  OAI22_X1 U22512 ( .A1(n25378), .A2(n20840), .B1(n25786), .B2(n25370), .ZN(
        n5440) );
  OAI22_X1 U22513 ( .A1(n25378), .A2(n20839), .B1(n25789), .B2(n25370), .ZN(
        n5441) );
  OAI22_X1 U22514 ( .A1(n25378), .A2(n20838), .B1(n25792), .B2(n25370), .ZN(
        n5442) );
  OAI22_X1 U22515 ( .A1(n25378), .A2(n20837), .B1(n25795), .B2(n25370), .ZN(
        n5443) );
  OAI22_X1 U22516 ( .A1(n25378), .A2(n20836), .B1(n25798), .B2(n25370), .ZN(
        n5444) );
  OAI22_X1 U22517 ( .A1(n25378), .A2(n20835), .B1(n25801), .B2(n25370), .ZN(
        n5445) );
  OAI22_X1 U22518 ( .A1(n25378), .A2(n20834), .B1(n25804), .B2(n25370), .ZN(
        n5446) );
  OAI22_X1 U22519 ( .A1(n25378), .A2(n20833), .B1(n25807), .B2(n25370), .ZN(
        n5447) );
  OAI22_X1 U22520 ( .A1(n25378), .A2(n20832), .B1(n25810), .B2(n25370), .ZN(
        n5448) );
  OAI22_X1 U22521 ( .A1(n25378), .A2(n20831), .B1(n25813), .B2(n25370), .ZN(
        n5449) );
  OAI22_X1 U22522 ( .A1(n25378), .A2(n20830), .B1(n25816), .B2(n25370), .ZN(
        n5450) );
  OAI22_X1 U22523 ( .A1(n25379), .A2(n20829), .B1(n25819), .B2(n25371), .ZN(
        n5451) );
  OAI22_X1 U22524 ( .A1(n25379), .A2(n20828), .B1(n25822), .B2(n25371), .ZN(
        n5452) );
  OAI22_X1 U22525 ( .A1(n25379), .A2(n20827), .B1(n25825), .B2(n25371), .ZN(
        n5453) );
  OAI22_X1 U22526 ( .A1(n25379), .A2(n20826), .B1(n25828), .B2(n25371), .ZN(
        n5454) );
  OAI22_X1 U22527 ( .A1(n25379), .A2(n20825), .B1(n25831), .B2(n25371), .ZN(
        n5455) );
  OAI22_X1 U22528 ( .A1(n25379), .A2(n20824), .B1(n25834), .B2(n25371), .ZN(
        n5456) );
  OAI22_X1 U22529 ( .A1(n25379), .A2(n20823), .B1(n25837), .B2(n25371), .ZN(
        n5457) );
  OAI22_X1 U22530 ( .A1(n25379), .A2(n20822), .B1(n25840), .B2(n25371), .ZN(
        n5458) );
  OAI22_X1 U22531 ( .A1(n25379), .A2(n20821), .B1(n25843), .B2(n25371), .ZN(
        n5459) );
  OAI22_X1 U22532 ( .A1(n25379), .A2(n20820), .B1(n25846), .B2(n25371), .ZN(
        n5460) );
  OAI22_X1 U22533 ( .A1(n25379), .A2(n20819), .B1(n25849), .B2(n25371), .ZN(
        n5461) );
  OAI22_X1 U22534 ( .A1(n25379), .A2(n20818), .B1(n25852), .B2(n25371), .ZN(
        n5462) );
  OAI22_X1 U22535 ( .A1(n25379), .A2(n20817), .B1(n25855), .B2(n25372), .ZN(
        n5463) );
  OAI22_X1 U22536 ( .A1(n25380), .A2(n20816), .B1(n25858), .B2(n25372), .ZN(
        n5464) );
  OAI22_X1 U22537 ( .A1(n25380), .A2(n20815), .B1(n25861), .B2(n25372), .ZN(
        n5465) );
  OAI22_X1 U22538 ( .A1(n25380), .A2(n20814), .B1(n25864), .B2(n25372), .ZN(
        n5466) );
  OAI22_X1 U22539 ( .A1(n25380), .A2(n20813), .B1(n25867), .B2(n25372), .ZN(
        n5467) );
  OAI22_X1 U22540 ( .A1(n25380), .A2(n20812), .B1(n25870), .B2(n25372), .ZN(
        n5468) );
  OAI22_X1 U22541 ( .A1(n25380), .A2(n20811), .B1(n25873), .B2(n25372), .ZN(
        n5469) );
  OAI22_X1 U22542 ( .A1(n25380), .A2(n20810), .B1(n25876), .B2(n25372), .ZN(
        n5470) );
  OAI22_X1 U22543 ( .A1(n25380), .A2(n20809), .B1(n25879), .B2(n25372), .ZN(
        n5471) );
  OAI22_X1 U22544 ( .A1(n25380), .A2(n20808), .B1(n25882), .B2(n25372), .ZN(
        n5472) );
  OAI22_X1 U22545 ( .A1(n25380), .A2(n20807), .B1(n25885), .B2(n25372), .ZN(
        n5473) );
  OAI22_X1 U22546 ( .A1(n25380), .A2(n20806), .B1(n25888), .B2(n25372), .ZN(
        n5474) );
  OAI22_X1 U22547 ( .A1(n25380), .A2(n20805), .B1(n25891), .B2(n25373), .ZN(
        n5475) );
  OAI22_X1 U22548 ( .A1(n25380), .A2(n20804), .B1(n25894), .B2(n25373), .ZN(
        n5476) );
  OAI22_X1 U22549 ( .A1(n25381), .A2(n20803), .B1(n25897), .B2(n25373), .ZN(
        n5477) );
  OAI22_X1 U22550 ( .A1(n25381), .A2(n20802), .B1(n25900), .B2(n25373), .ZN(
        n5478) );
  OAI22_X1 U22551 ( .A1(n25381), .A2(n20801), .B1(n25903), .B2(n25373), .ZN(
        n5479) );
  OAI22_X1 U22552 ( .A1(n25381), .A2(n20800), .B1(n25906), .B2(n25373), .ZN(
        n5480) );
  OAI22_X1 U22553 ( .A1(n25381), .A2(n20799), .B1(n25909), .B2(n25373), .ZN(
        n5481) );
  OAI22_X1 U22554 ( .A1(n25381), .A2(n20798), .B1(n25912), .B2(n25373), .ZN(
        n5482) );
  OAI22_X1 U22555 ( .A1(n25381), .A2(n20797), .B1(n25915), .B2(n25373), .ZN(
        n5483) );
  OAI22_X1 U22556 ( .A1(n25381), .A2(n20796), .B1(n25918), .B2(n25373), .ZN(
        n5484) );
  OAI22_X1 U22557 ( .A1(n25381), .A2(n20795), .B1(n25921), .B2(n25373), .ZN(
        n5485) );
  OAI22_X1 U22558 ( .A1(n25381), .A2(n20794), .B1(n25924), .B2(n25373), .ZN(
        n5486) );
  OAI22_X1 U22559 ( .A1(n25381), .A2(n20793), .B1(n25927), .B2(n25374), .ZN(
        n5487) );
  OAI22_X1 U22560 ( .A1(n25381), .A2(n20792), .B1(n25930), .B2(n25374), .ZN(
        n5488) );
  OAI22_X1 U22561 ( .A1(n25381), .A2(n20791), .B1(n25933), .B2(n25374), .ZN(
        n5489) );
  OAI22_X1 U22562 ( .A1(n25382), .A2(n20790), .B1(n25936), .B2(n25374), .ZN(
        n5490) );
  OAI22_X1 U22563 ( .A1(n25382), .A2(n20789), .B1(n25939), .B2(n25374), .ZN(
        n5491) );
  OAI22_X1 U22564 ( .A1(n25382), .A2(n20788), .B1(n25942), .B2(n25374), .ZN(
        n5492) );
  OAI22_X1 U22565 ( .A1(n25382), .A2(n20787), .B1(n25945), .B2(n25374), .ZN(
        n5493) );
  OAI22_X1 U22566 ( .A1(n25382), .A2(n20786), .B1(n25948), .B2(n25374), .ZN(
        n5494) );
  OAI22_X1 U22567 ( .A1(n25382), .A2(n20785), .B1(n25951), .B2(n25374), .ZN(
        n5495) );
  OAI22_X1 U22568 ( .A1(n25382), .A2(n20784), .B1(n25954), .B2(n25374), .ZN(
        n5496) );
  OAI22_X1 U22569 ( .A1(n25382), .A2(n20783), .B1(n25957), .B2(n25374), .ZN(
        n5497) );
  OAI22_X1 U22570 ( .A1(n25382), .A2(n20782), .B1(n25960), .B2(n25374), .ZN(
        n5498) );
  OAI22_X1 U22571 ( .A1(n25417), .A2(n20581), .B1(n25783), .B2(n25409), .ZN(
        n5631) );
  OAI22_X1 U22572 ( .A1(n25417), .A2(n20580), .B1(n25786), .B2(n25409), .ZN(
        n5632) );
  OAI22_X1 U22573 ( .A1(n25417), .A2(n20579), .B1(n25789), .B2(n25409), .ZN(
        n5633) );
  OAI22_X1 U22574 ( .A1(n25417), .A2(n20578), .B1(n25792), .B2(n25409), .ZN(
        n5634) );
  OAI22_X1 U22575 ( .A1(n25417), .A2(n20577), .B1(n25795), .B2(n25409), .ZN(
        n5635) );
  OAI22_X1 U22576 ( .A1(n25417), .A2(n20576), .B1(n25798), .B2(n25409), .ZN(
        n5636) );
  OAI22_X1 U22577 ( .A1(n25417), .A2(n20575), .B1(n25801), .B2(n25409), .ZN(
        n5637) );
  OAI22_X1 U22578 ( .A1(n25417), .A2(n20574), .B1(n25804), .B2(n25409), .ZN(
        n5638) );
  OAI22_X1 U22579 ( .A1(n25417), .A2(n20573), .B1(n25807), .B2(n25409), .ZN(
        n5639) );
  OAI22_X1 U22580 ( .A1(n25417), .A2(n20572), .B1(n25810), .B2(n25409), .ZN(
        n5640) );
  OAI22_X1 U22581 ( .A1(n25417), .A2(n20571), .B1(n25813), .B2(n25409), .ZN(
        n5641) );
  OAI22_X1 U22582 ( .A1(n25417), .A2(n20570), .B1(n25816), .B2(n25409), .ZN(
        n5642) );
  OAI22_X1 U22583 ( .A1(n25418), .A2(n20569), .B1(n25819), .B2(n25410), .ZN(
        n5643) );
  OAI22_X1 U22584 ( .A1(n25418), .A2(n20568), .B1(n25822), .B2(n25410), .ZN(
        n5644) );
  OAI22_X1 U22585 ( .A1(n25418), .A2(n20567), .B1(n25825), .B2(n25410), .ZN(
        n5645) );
  OAI22_X1 U22586 ( .A1(n25418), .A2(n20566), .B1(n25828), .B2(n25410), .ZN(
        n5646) );
  OAI22_X1 U22587 ( .A1(n25418), .A2(n20565), .B1(n25831), .B2(n25410), .ZN(
        n5647) );
  OAI22_X1 U22588 ( .A1(n25418), .A2(n20564), .B1(n25834), .B2(n25410), .ZN(
        n5648) );
  OAI22_X1 U22589 ( .A1(n25418), .A2(n20563), .B1(n25837), .B2(n25410), .ZN(
        n5649) );
  OAI22_X1 U22590 ( .A1(n25418), .A2(n20562), .B1(n25840), .B2(n25410), .ZN(
        n5650) );
  OAI22_X1 U22591 ( .A1(n25418), .A2(n20561), .B1(n25843), .B2(n25410), .ZN(
        n5651) );
  OAI22_X1 U22592 ( .A1(n25418), .A2(n20560), .B1(n25846), .B2(n25410), .ZN(
        n5652) );
  OAI22_X1 U22593 ( .A1(n25418), .A2(n20559), .B1(n25849), .B2(n25410), .ZN(
        n5653) );
  OAI22_X1 U22594 ( .A1(n25418), .A2(n20558), .B1(n25852), .B2(n25410), .ZN(
        n5654) );
  OAI22_X1 U22595 ( .A1(n25418), .A2(n20557), .B1(n25855), .B2(n25411), .ZN(
        n5655) );
  OAI22_X1 U22596 ( .A1(n25419), .A2(n20556), .B1(n25858), .B2(n25411), .ZN(
        n5656) );
  OAI22_X1 U22597 ( .A1(n25419), .A2(n20555), .B1(n25861), .B2(n25411), .ZN(
        n5657) );
  OAI22_X1 U22598 ( .A1(n25419), .A2(n20554), .B1(n25864), .B2(n25411), .ZN(
        n5658) );
  OAI22_X1 U22599 ( .A1(n25419), .A2(n20553), .B1(n25867), .B2(n25411), .ZN(
        n5659) );
  OAI22_X1 U22600 ( .A1(n25419), .A2(n20552), .B1(n25870), .B2(n25411), .ZN(
        n5660) );
  OAI22_X1 U22601 ( .A1(n25419), .A2(n20551), .B1(n25873), .B2(n25411), .ZN(
        n5661) );
  OAI22_X1 U22602 ( .A1(n25419), .A2(n20550), .B1(n25876), .B2(n25411), .ZN(
        n5662) );
  OAI22_X1 U22603 ( .A1(n25419), .A2(n20549), .B1(n25879), .B2(n25411), .ZN(
        n5663) );
  OAI22_X1 U22604 ( .A1(n25419), .A2(n20548), .B1(n25882), .B2(n25411), .ZN(
        n5664) );
  OAI22_X1 U22605 ( .A1(n25419), .A2(n20547), .B1(n25885), .B2(n25411), .ZN(
        n5665) );
  OAI22_X1 U22606 ( .A1(n25419), .A2(n20546), .B1(n25888), .B2(n25411), .ZN(
        n5666) );
  OAI22_X1 U22607 ( .A1(n25419), .A2(n20545), .B1(n25891), .B2(n25412), .ZN(
        n5667) );
  OAI22_X1 U22608 ( .A1(n25419), .A2(n20544), .B1(n25894), .B2(n25412), .ZN(
        n5668) );
  OAI22_X1 U22609 ( .A1(n25420), .A2(n20543), .B1(n25897), .B2(n25412), .ZN(
        n5669) );
  OAI22_X1 U22610 ( .A1(n25420), .A2(n20542), .B1(n25900), .B2(n25412), .ZN(
        n5670) );
  OAI22_X1 U22611 ( .A1(n25420), .A2(n20541), .B1(n25903), .B2(n25412), .ZN(
        n5671) );
  OAI22_X1 U22612 ( .A1(n25420), .A2(n20540), .B1(n25906), .B2(n25412), .ZN(
        n5672) );
  OAI22_X1 U22613 ( .A1(n25420), .A2(n20539), .B1(n25909), .B2(n25412), .ZN(
        n5673) );
  OAI22_X1 U22614 ( .A1(n25420), .A2(n20538), .B1(n25912), .B2(n25412), .ZN(
        n5674) );
  OAI22_X1 U22615 ( .A1(n25420), .A2(n20537), .B1(n25915), .B2(n25412), .ZN(
        n5675) );
  OAI22_X1 U22616 ( .A1(n25420), .A2(n20536), .B1(n25918), .B2(n25412), .ZN(
        n5676) );
  OAI22_X1 U22617 ( .A1(n25420), .A2(n20535), .B1(n25921), .B2(n25412), .ZN(
        n5677) );
  OAI22_X1 U22618 ( .A1(n25420), .A2(n20534), .B1(n25924), .B2(n25412), .ZN(
        n5678) );
  OAI22_X1 U22619 ( .A1(n25420), .A2(n20533), .B1(n25927), .B2(n25413), .ZN(
        n5679) );
  OAI22_X1 U22620 ( .A1(n25420), .A2(n20532), .B1(n25930), .B2(n25413), .ZN(
        n5680) );
  OAI22_X1 U22621 ( .A1(n25420), .A2(n20531), .B1(n25933), .B2(n25413), .ZN(
        n5681) );
  OAI22_X1 U22622 ( .A1(n25421), .A2(n20530), .B1(n25936), .B2(n25413), .ZN(
        n5682) );
  OAI22_X1 U22623 ( .A1(n25421), .A2(n20529), .B1(n25939), .B2(n25413), .ZN(
        n5683) );
  OAI22_X1 U22624 ( .A1(n25421), .A2(n20528), .B1(n25942), .B2(n25413), .ZN(
        n5684) );
  OAI22_X1 U22625 ( .A1(n25421), .A2(n20527), .B1(n25945), .B2(n25413), .ZN(
        n5685) );
  OAI22_X1 U22626 ( .A1(n25421), .A2(n20526), .B1(n25948), .B2(n25413), .ZN(
        n5686) );
  OAI22_X1 U22627 ( .A1(n25421), .A2(n20525), .B1(n25951), .B2(n25413), .ZN(
        n5687) );
  OAI22_X1 U22628 ( .A1(n25421), .A2(n20524), .B1(n25954), .B2(n25413), .ZN(
        n5688) );
  OAI22_X1 U22629 ( .A1(n25421), .A2(n20523), .B1(n25957), .B2(n25413), .ZN(
        n5689) );
  OAI22_X1 U22630 ( .A1(n25421), .A2(n20522), .B1(n25960), .B2(n25413), .ZN(
        n5690) );
  OAI22_X1 U22631 ( .A1(n25391), .A2(n20521), .B1(n25783), .B2(n25383), .ZN(
        n5503) );
  OAI22_X1 U22632 ( .A1(n25391), .A2(n20520), .B1(n25786), .B2(n25383), .ZN(
        n5504) );
  OAI22_X1 U22633 ( .A1(n25391), .A2(n20519), .B1(n25789), .B2(n25383), .ZN(
        n5505) );
  OAI22_X1 U22634 ( .A1(n25391), .A2(n20518), .B1(n25792), .B2(n25383), .ZN(
        n5506) );
  OAI22_X1 U22635 ( .A1(n25391), .A2(n20517), .B1(n25795), .B2(n25383), .ZN(
        n5507) );
  OAI22_X1 U22636 ( .A1(n25391), .A2(n20516), .B1(n25798), .B2(n25383), .ZN(
        n5508) );
  OAI22_X1 U22637 ( .A1(n25391), .A2(n20515), .B1(n25801), .B2(n25383), .ZN(
        n5509) );
  OAI22_X1 U22638 ( .A1(n25391), .A2(n20514), .B1(n25804), .B2(n25383), .ZN(
        n5510) );
  OAI22_X1 U22639 ( .A1(n25391), .A2(n20513), .B1(n25807), .B2(n25383), .ZN(
        n5511) );
  OAI22_X1 U22640 ( .A1(n25391), .A2(n20512), .B1(n25810), .B2(n25383), .ZN(
        n5512) );
  OAI22_X1 U22641 ( .A1(n25391), .A2(n20511), .B1(n25813), .B2(n25383), .ZN(
        n5513) );
  OAI22_X1 U22642 ( .A1(n25391), .A2(n20510), .B1(n25816), .B2(n25383), .ZN(
        n5514) );
  OAI22_X1 U22643 ( .A1(n25392), .A2(n20509), .B1(n25819), .B2(n25384), .ZN(
        n5515) );
  OAI22_X1 U22644 ( .A1(n25392), .A2(n20508), .B1(n25822), .B2(n25384), .ZN(
        n5516) );
  OAI22_X1 U22645 ( .A1(n25392), .A2(n20507), .B1(n25825), .B2(n25384), .ZN(
        n5517) );
  OAI22_X1 U22646 ( .A1(n25392), .A2(n20506), .B1(n25828), .B2(n25384), .ZN(
        n5518) );
  OAI22_X1 U22647 ( .A1(n25392), .A2(n20505), .B1(n25831), .B2(n25384), .ZN(
        n5519) );
  OAI22_X1 U22648 ( .A1(n25392), .A2(n20504), .B1(n25834), .B2(n25384), .ZN(
        n5520) );
  OAI22_X1 U22649 ( .A1(n25392), .A2(n20503), .B1(n25837), .B2(n25384), .ZN(
        n5521) );
  OAI22_X1 U22650 ( .A1(n25392), .A2(n20502), .B1(n25840), .B2(n25384), .ZN(
        n5522) );
  OAI22_X1 U22651 ( .A1(n25392), .A2(n20501), .B1(n25843), .B2(n25384), .ZN(
        n5523) );
  OAI22_X1 U22652 ( .A1(n25392), .A2(n20500), .B1(n25846), .B2(n25384), .ZN(
        n5524) );
  OAI22_X1 U22653 ( .A1(n25392), .A2(n20499), .B1(n25849), .B2(n25384), .ZN(
        n5525) );
  OAI22_X1 U22654 ( .A1(n25392), .A2(n20498), .B1(n25852), .B2(n25384), .ZN(
        n5526) );
  OAI22_X1 U22655 ( .A1(n25392), .A2(n20497), .B1(n25855), .B2(n25385), .ZN(
        n5527) );
  OAI22_X1 U22656 ( .A1(n25393), .A2(n20496), .B1(n25858), .B2(n25385), .ZN(
        n5528) );
  OAI22_X1 U22657 ( .A1(n25393), .A2(n20495), .B1(n25861), .B2(n25385), .ZN(
        n5529) );
  OAI22_X1 U22658 ( .A1(n25393), .A2(n20494), .B1(n25864), .B2(n25385), .ZN(
        n5530) );
  OAI22_X1 U22659 ( .A1(n25393), .A2(n20493), .B1(n25867), .B2(n25385), .ZN(
        n5531) );
  OAI22_X1 U22660 ( .A1(n25393), .A2(n20492), .B1(n25870), .B2(n25385), .ZN(
        n5532) );
  OAI22_X1 U22661 ( .A1(n25393), .A2(n20491), .B1(n25873), .B2(n25385), .ZN(
        n5533) );
  OAI22_X1 U22662 ( .A1(n25393), .A2(n20490), .B1(n25876), .B2(n25385), .ZN(
        n5534) );
  OAI22_X1 U22663 ( .A1(n25393), .A2(n20489), .B1(n25879), .B2(n25385), .ZN(
        n5535) );
  OAI22_X1 U22664 ( .A1(n25393), .A2(n20488), .B1(n25882), .B2(n25385), .ZN(
        n5536) );
  OAI22_X1 U22665 ( .A1(n25393), .A2(n20487), .B1(n25885), .B2(n25385), .ZN(
        n5537) );
  OAI22_X1 U22666 ( .A1(n25393), .A2(n20486), .B1(n25888), .B2(n25385), .ZN(
        n5538) );
  OAI22_X1 U22667 ( .A1(n25393), .A2(n20485), .B1(n25891), .B2(n25386), .ZN(
        n5539) );
  OAI22_X1 U22668 ( .A1(n25393), .A2(n20484), .B1(n25894), .B2(n25386), .ZN(
        n5540) );
  OAI22_X1 U22669 ( .A1(n25394), .A2(n20483), .B1(n25897), .B2(n25386), .ZN(
        n5541) );
  OAI22_X1 U22670 ( .A1(n25394), .A2(n20482), .B1(n25900), .B2(n25386), .ZN(
        n5542) );
  OAI22_X1 U22671 ( .A1(n25394), .A2(n20481), .B1(n25903), .B2(n25386), .ZN(
        n5543) );
  OAI22_X1 U22672 ( .A1(n25394), .A2(n20480), .B1(n25906), .B2(n25386), .ZN(
        n5544) );
  OAI22_X1 U22673 ( .A1(n25394), .A2(n20479), .B1(n25909), .B2(n25386), .ZN(
        n5545) );
  OAI22_X1 U22674 ( .A1(n25394), .A2(n20478), .B1(n25912), .B2(n25386), .ZN(
        n5546) );
  OAI22_X1 U22675 ( .A1(n25394), .A2(n20477), .B1(n25915), .B2(n25386), .ZN(
        n5547) );
  OAI22_X1 U22676 ( .A1(n25394), .A2(n20476), .B1(n25918), .B2(n25386), .ZN(
        n5548) );
  OAI22_X1 U22677 ( .A1(n25394), .A2(n20475), .B1(n25921), .B2(n25386), .ZN(
        n5549) );
  OAI22_X1 U22678 ( .A1(n25394), .A2(n20474), .B1(n25924), .B2(n25386), .ZN(
        n5550) );
  OAI22_X1 U22679 ( .A1(n25394), .A2(n20473), .B1(n25927), .B2(n25387), .ZN(
        n5551) );
  OAI22_X1 U22680 ( .A1(n25394), .A2(n20472), .B1(n25930), .B2(n25387), .ZN(
        n5552) );
  OAI22_X1 U22681 ( .A1(n25394), .A2(n20471), .B1(n25933), .B2(n25387), .ZN(
        n5553) );
  OAI22_X1 U22682 ( .A1(n25395), .A2(n20470), .B1(n25936), .B2(n25387), .ZN(
        n5554) );
  OAI22_X1 U22683 ( .A1(n25395), .A2(n20469), .B1(n25939), .B2(n25387), .ZN(
        n5555) );
  OAI22_X1 U22684 ( .A1(n25395), .A2(n20468), .B1(n25942), .B2(n25387), .ZN(
        n5556) );
  OAI22_X1 U22685 ( .A1(n25395), .A2(n20467), .B1(n25945), .B2(n25387), .ZN(
        n5557) );
  OAI22_X1 U22686 ( .A1(n25395), .A2(n20466), .B1(n25948), .B2(n25387), .ZN(
        n5558) );
  OAI22_X1 U22687 ( .A1(n25395), .A2(n20465), .B1(n25951), .B2(n25387), .ZN(
        n5559) );
  OAI22_X1 U22688 ( .A1(n25395), .A2(n20464), .B1(n25954), .B2(n25387), .ZN(
        n5560) );
  OAI22_X1 U22689 ( .A1(n25395), .A2(n20463), .B1(n25957), .B2(n25387), .ZN(
        n5561) );
  OAI22_X1 U22690 ( .A1(n25395), .A2(n20462), .B1(n25960), .B2(n25387), .ZN(
        n5562) );
  OAI22_X1 U22691 ( .A1(n25469), .A2(n21349), .B1(n25782), .B2(n25461), .ZN(
        n5887) );
  OAI22_X1 U22692 ( .A1(n25469), .A2(n21348), .B1(n25785), .B2(n25461), .ZN(
        n5888) );
  OAI22_X1 U22693 ( .A1(n25469), .A2(n21347), .B1(n25788), .B2(n25461), .ZN(
        n5889) );
  OAI22_X1 U22694 ( .A1(n25469), .A2(n21346), .B1(n25791), .B2(n25461), .ZN(
        n5890) );
  OAI22_X1 U22695 ( .A1(n25469), .A2(n21345), .B1(n25794), .B2(n25461), .ZN(
        n5891) );
  OAI22_X1 U22696 ( .A1(n25469), .A2(n21344), .B1(n25797), .B2(n25461), .ZN(
        n5892) );
  OAI22_X1 U22697 ( .A1(n25469), .A2(n21343), .B1(n25800), .B2(n25461), .ZN(
        n5893) );
  OAI22_X1 U22698 ( .A1(n25469), .A2(n21342), .B1(n25803), .B2(n25461), .ZN(
        n5894) );
  OAI22_X1 U22699 ( .A1(n25469), .A2(n21341), .B1(n25806), .B2(n25461), .ZN(
        n5895) );
  OAI22_X1 U22700 ( .A1(n25469), .A2(n21340), .B1(n25809), .B2(n25461), .ZN(
        n5896) );
  OAI22_X1 U22701 ( .A1(n25469), .A2(n21339), .B1(n25812), .B2(n25461), .ZN(
        n5897) );
  OAI22_X1 U22702 ( .A1(n25469), .A2(n21338), .B1(n25815), .B2(n25461), .ZN(
        n5898) );
  OAI22_X1 U22703 ( .A1(n25470), .A2(n21337), .B1(n25818), .B2(n25462), .ZN(
        n5899) );
  OAI22_X1 U22704 ( .A1(n25470), .A2(n21336), .B1(n25821), .B2(n25462), .ZN(
        n5900) );
  OAI22_X1 U22705 ( .A1(n25470), .A2(n21335), .B1(n25824), .B2(n25462), .ZN(
        n5901) );
  OAI22_X1 U22706 ( .A1(n25470), .A2(n21334), .B1(n25827), .B2(n25462), .ZN(
        n5902) );
  OAI22_X1 U22707 ( .A1(n25470), .A2(n21333), .B1(n25830), .B2(n25462), .ZN(
        n5903) );
  OAI22_X1 U22708 ( .A1(n25470), .A2(n21332), .B1(n25833), .B2(n25462), .ZN(
        n5904) );
  OAI22_X1 U22709 ( .A1(n25470), .A2(n21331), .B1(n25836), .B2(n25462), .ZN(
        n5905) );
  OAI22_X1 U22710 ( .A1(n25470), .A2(n21330), .B1(n25839), .B2(n25462), .ZN(
        n5906) );
  OAI22_X1 U22711 ( .A1(n25470), .A2(n21329), .B1(n25842), .B2(n25462), .ZN(
        n5907) );
  OAI22_X1 U22712 ( .A1(n25470), .A2(n21328), .B1(n25845), .B2(n25462), .ZN(
        n5908) );
  OAI22_X1 U22713 ( .A1(n25470), .A2(n21327), .B1(n25848), .B2(n25462), .ZN(
        n5909) );
  OAI22_X1 U22714 ( .A1(n25470), .A2(n21326), .B1(n25851), .B2(n25462), .ZN(
        n5910) );
  OAI22_X1 U22715 ( .A1(n25470), .A2(n21325), .B1(n25854), .B2(n25463), .ZN(
        n5911) );
  OAI22_X1 U22716 ( .A1(n25471), .A2(n21324), .B1(n25857), .B2(n25463), .ZN(
        n5912) );
  OAI22_X1 U22717 ( .A1(n25471), .A2(n21323), .B1(n25860), .B2(n25463), .ZN(
        n5913) );
  OAI22_X1 U22718 ( .A1(n25471), .A2(n21322), .B1(n25863), .B2(n25463), .ZN(
        n5914) );
  OAI22_X1 U22719 ( .A1(n25471), .A2(n21321), .B1(n25866), .B2(n25463), .ZN(
        n5915) );
  OAI22_X1 U22720 ( .A1(n25471), .A2(n21320), .B1(n25869), .B2(n25463), .ZN(
        n5916) );
  OAI22_X1 U22721 ( .A1(n25471), .A2(n21319), .B1(n25872), .B2(n25463), .ZN(
        n5917) );
  OAI22_X1 U22722 ( .A1(n25471), .A2(n21318), .B1(n25875), .B2(n25463), .ZN(
        n5918) );
  OAI22_X1 U22723 ( .A1(n25471), .A2(n21317), .B1(n25878), .B2(n25463), .ZN(
        n5919) );
  OAI22_X1 U22724 ( .A1(n25471), .A2(n21316), .B1(n25881), .B2(n25463), .ZN(
        n5920) );
  OAI22_X1 U22725 ( .A1(n25471), .A2(n21315), .B1(n25884), .B2(n25463), .ZN(
        n5921) );
  OAI22_X1 U22726 ( .A1(n25471), .A2(n21314), .B1(n25887), .B2(n25463), .ZN(
        n5922) );
  OAI22_X1 U22727 ( .A1(n25471), .A2(n21313), .B1(n25890), .B2(n25464), .ZN(
        n5923) );
  OAI22_X1 U22728 ( .A1(n25471), .A2(n21312), .B1(n25893), .B2(n25464), .ZN(
        n5924) );
  OAI22_X1 U22729 ( .A1(n25472), .A2(n21311), .B1(n25896), .B2(n25464), .ZN(
        n5925) );
  OAI22_X1 U22730 ( .A1(n25472), .A2(n21310), .B1(n25899), .B2(n25464), .ZN(
        n5926) );
  OAI22_X1 U22731 ( .A1(n25472), .A2(n21309), .B1(n25902), .B2(n25464), .ZN(
        n5927) );
  OAI22_X1 U22732 ( .A1(n25472), .A2(n21308), .B1(n25905), .B2(n25464), .ZN(
        n5928) );
  OAI22_X1 U22733 ( .A1(n25472), .A2(n21307), .B1(n25908), .B2(n25464), .ZN(
        n5929) );
  OAI22_X1 U22734 ( .A1(n25472), .A2(n21306), .B1(n25911), .B2(n25464), .ZN(
        n5930) );
  OAI22_X1 U22735 ( .A1(n25472), .A2(n21305), .B1(n25914), .B2(n25464), .ZN(
        n5931) );
  OAI22_X1 U22736 ( .A1(n25472), .A2(n21304), .B1(n25917), .B2(n25464), .ZN(
        n5932) );
  OAI22_X1 U22737 ( .A1(n25472), .A2(n21303), .B1(n25920), .B2(n25464), .ZN(
        n5933) );
  OAI22_X1 U22738 ( .A1(n25472), .A2(n21302), .B1(n25923), .B2(n25464), .ZN(
        n5934) );
  OAI22_X1 U22739 ( .A1(n25472), .A2(n21301), .B1(n25926), .B2(n25465), .ZN(
        n5935) );
  OAI22_X1 U22740 ( .A1(n25472), .A2(n21300), .B1(n25929), .B2(n25465), .ZN(
        n5936) );
  OAI22_X1 U22741 ( .A1(n25472), .A2(n21299), .B1(n25932), .B2(n25465), .ZN(
        n5937) );
  OAI22_X1 U22742 ( .A1(n25473), .A2(n21298), .B1(n25935), .B2(n25465), .ZN(
        n5938) );
  OAI22_X1 U22743 ( .A1(n25473), .A2(n21297), .B1(n25938), .B2(n25465), .ZN(
        n5939) );
  OAI22_X1 U22744 ( .A1(n25473), .A2(n21296), .B1(n25941), .B2(n25465), .ZN(
        n5940) );
  OAI22_X1 U22745 ( .A1(n25473), .A2(n21295), .B1(n25944), .B2(n25465), .ZN(
        n5941) );
  OAI22_X1 U22746 ( .A1(n25473), .A2(n21294), .B1(n25947), .B2(n25465), .ZN(
        n5942) );
  OAI22_X1 U22747 ( .A1(n25473), .A2(n21293), .B1(n25950), .B2(n25465), .ZN(
        n5943) );
  OAI22_X1 U22748 ( .A1(n25473), .A2(n21292), .B1(n25953), .B2(n25465), .ZN(
        n5944) );
  OAI22_X1 U22749 ( .A1(n25473), .A2(n21291), .B1(n25956), .B2(n25465), .ZN(
        n5945) );
  OAI22_X1 U22750 ( .A1(n25473), .A2(n21290), .B1(n25959), .B2(n25465), .ZN(
        n5946) );
  OAI22_X1 U22751 ( .A1(n25649), .A2(n20645), .B1(n25781), .B2(n25641), .ZN(
        n6783) );
  OAI22_X1 U22752 ( .A1(n25649), .A2(n20644), .B1(n25784), .B2(n25641), .ZN(
        n6784) );
  OAI22_X1 U22753 ( .A1(n25649), .A2(n20643), .B1(n25787), .B2(n25641), .ZN(
        n6785) );
  OAI22_X1 U22754 ( .A1(n25649), .A2(n20642), .B1(n25790), .B2(n25641), .ZN(
        n6786) );
  OAI22_X1 U22755 ( .A1(n25649), .A2(n20641), .B1(n25793), .B2(n25641), .ZN(
        n6787) );
  OAI22_X1 U22756 ( .A1(n25649), .A2(n20640), .B1(n25796), .B2(n25641), .ZN(
        n6788) );
  OAI22_X1 U22757 ( .A1(n25649), .A2(n20639), .B1(n25799), .B2(n25641), .ZN(
        n6789) );
  OAI22_X1 U22758 ( .A1(n25649), .A2(n20638), .B1(n25802), .B2(n25641), .ZN(
        n6790) );
  OAI22_X1 U22759 ( .A1(n25649), .A2(n20637), .B1(n25805), .B2(n25641), .ZN(
        n6791) );
  OAI22_X1 U22760 ( .A1(n25649), .A2(n20636), .B1(n25808), .B2(n25641), .ZN(
        n6792) );
  OAI22_X1 U22761 ( .A1(n25649), .A2(n20635), .B1(n25811), .B2(n25641), .ZN(
        n6793) );
  OAI22_X1 U22762 ( .A1(n25649), .A2(n20634), .B1(n25814), .B2(n25641), .ZN(
        n6794) );
  OAI22_X1 U22763 ( .A1(n25650), .A2(n20633), .B1(n25817), .B2(n25642), .ZN(
        n6795) );
  OAI22_X1 U22764 ( .A1(n25650), .A2(n20632), .B1(n25820), .B2(n25642), .ZN(
        n6796) );
  OAI22_X1 U22765 ( .A1(n25650), .A2(n20631), .B1(n25823), .B2(n25642), .ZN(
        n6797) );
  OAI22_X1 U22766 ( .A1(n25650), .A2(n20630), .B1(n25826), .B2(n25642), .ZN(
        n6798) );
  OAI22_X1 U22767 ( .A1(n25650), .A2(n20629), .B1(n25829), .B2(n25642), .ZN(
        n6799) );
  OAI22_X1 U22768 ( .A1(n25650), .A2(n20628), .B1(n25832), .B2(n25642), .ZN(
        n6800) );
  OAI22_X1 U22769 ( .A1(n25650), .A2(n20627), .B1(n25835), .B2(n25642), .ZN(
        n6801) );
  OAI22_X1 U22770 ( .A1(n25650), .A2(n20626), .B1(n25838), .B2(n25642), .ZN(
        n6802) );
  OAI22_X1 U22771 ( .A1(n25650), .A2(n20625), .B1(n25841), .B2(n25642), .ZN(
        n6803) );
  OAI22_X1 U22772 ( .A1(n25650), .A2(n20624), .B1(n25844), .B2(n25642), .ZN(
        n6804) );
  OAI22_X1 U22773 ( .A1(n25650), .A2(n20623), .B1(n25847), .B2(n25642), .ZN(
        n6805) );
  OAI22_X1 U22774 ( .A1(n25650), .A2(n20622), .B1(n25850), .B2(n25642), .ZN(
        n6806) );
  OAI22_X1 U22775 ( .A1(n25650), .A2(n20621), .B1(n25853), .B2(n25643), .ZN(
        n6807) );
  OAI22_X1 U22776 ( .A1(n25651), .A2(n20620), .B1(n25856), .B2(n25643), .ZN(
        n6808) );
  OAI22_X1 U22777 ( .A1(n25651), .A2(n20619), .B1(n25859), .B2(n25643), .ZN(
        n6809) );
  OAI22_X1 U22778 ( .A1(n25651), .A2(n20618), .B1(n25862), .B2(n25643), .ZN(
        n6810) );
  OAI22_X1 U22779 ( .A1(n25651), .A2(n20617), .B1(n25865), .B2(n25643), .ZN(
        n6811) );
  OAI22_X1 U22780 ( .A1(n25651), .A2(n20616), .B1(n25868), .B2(n25643), .ZN(
        n6812) );
  OAI22_X1 U22781 ( .A1(n25651), .A2(n20615), .B1(n25871), .B2(n25643), .ZN(
        n6813) );
  OAI22_X1 U22782 ( .A1(n25651), .A2(n20614), .B1(n25874), .B2(n25643), .ZN(
        n6814) );
  OAI22_X1 U22783 ( .A1(n25651), .A2(n20613), .B1(n25877), .B2(n25643), .ZN(
        n6815) );
  OAI22_X1 U22784 ( .A1(n25651), .A2(n20612), .B1(n25880), .B2(n25643), .ZN(
        n6816) );
  OAI22_X1 U22785 ( .A1(n25651), .A2(n20611), .B1(n25883), .B2(n25643), .ZN(
        n6817) );
  OAI22_X1 U22786 ( .A1(n25651), .A2(n20610), .B1(n25886), .B2(n25643), .ZN(
        n6818) );
  OAI22_X1 U22787 ( .A1(n25651), .A2(n20609), .B1(n25889), .B2(n25644), .ZN(
        n6819) );
  OAI22_X1 U22788 ( .A1(n25651), .A2(n20608), .B1(n25892), .B2(n25644), .ZN(
        n6820) );
  OAI22_X1 U22789 ( .A1(n25652), .A2(n20607), .B1(n25895), .B2(n25644), .ZN(
        n6821) );
  OAI22_X1 U22790 ( .A1(n25652), .A2(n20606), .B1(n25898), .B2(n25644), .ZN(
        n6822) );
  OAI22_X1 U22791 ( .A1(n25652), .A2(n20605), .B1(n25901), .B2(n25644), .ZN(
        n6823) );
  OAI22_X1 U22792 ( .A1(n25652), .A2(n20604), .B1(n25904), .B2(n25644), .ZN(
        n6824) );
  OAI22_X1 U22793 ( .A1(n25652), .A2(n20603), .B1(n25907), .B2(n25644), .ZN(
        n6825) );
  OAI22_X1 U22794 ( .A1(n25652), .A2(n20602), .B1(n25910), .B2(n25644), .ZN(
        n6826) );
  OAI22_X1 U22795 ( .A1(n25652), .A2(n20601), .B1(n25913), .B2(n25644), .ZN(
        n6827) );
  OAI22_X1 U22796 ( .A1(n25652), .A2(n20600), .B1(n25916), .B2(n25644), .ZN(
        n6828) );
  OAI22_X1 U22797 ( .A1(n25652), .A2(n20599), .B1(n25919), .B2(n25644), .ZN(
        n6829) );
  OAI22_X1 U22798 ( .A1(n25652), .A2(n20598), .B1(n25922), .B2(n25644), .ZN(
        n6830) );
  OAI22_X1 U22799 ( .A1(n25652), .A2(n20597), .B1(n25925), .B2(n25645), .ZN(
        n6831) );
  OAI22_X1 U22800 ( .A1(n25652), .A2(n20596), .B1(n25928), .B2(n25645), .ZN(
        n6832) );
  OAI22_X1 U22801 ( .A1(n25652), .A2(n20595), .B1(n25931), .B2(n25645), .ZN(
        n6833) );
  OAI22_X1 U22802 ( .A1(n25653), .A2(n20594), .B1(n25934), .B2(n25645), .ZN(
        n6834) );
  OAI22_X1 U22803 ( .A1(n25653), .A2(n20593), .B1(n25937), .B2(n25645), .ZN(
        n6835) );
  OAI22_X1 U22804 ( .A1(n25653), .A2(n20592), .B1(n25940), .B2(n25645), .ZN(
        n6836) );
  OAI22_X1 U22805 ( .A1(n25653), .A2(n20591), .B1(n25943), .B2(n25645), .ZN(
        n6837) );
  OAI22_X1 U22806 ( .A1(n25653), .A2(n20590), .B1(n25946), .B2(n25645), .ZN(
        n6838) );
  OAI22_X1 U22807 ( .A1(n25653), .A2(n20589), .B1(n25949), .B2(n25645), .ZN(
        n6839) );
  OAI22_X1 U22808 ( .A1(n25653), .A2(n20588), .B1(n25952), .B2(n25645), .ZN(
        n6840) );
  OAI22_X1 U22809 ( .A1(n25653), .A2(n20587), .B1(n25955), .B2(n25645), .ZN(
        n6841) );
  OAI22_X1 U22810 ( .A1(n25653), .A2(n20586), .B1(n25958), .B2(n25645), .ZN(
        n6842) );
  OAI22_X1 U22811 ( .A1(n25739), .A2(n20261), .B1(n25781), .B2(n25731), .ZN(
        n7231) );
  OAI22_X1 U22812 ( .A1(n25739), .A2(n20260), .B1(n25784), .B2(n25731), .ZN(
        n7232) );
  OAI22_X1 U22813 ( .A1(n25739), .A2(n20259), .B1(n25787), .B2(n25731), .ZN(
        n7233) );
  OAI22_X1 U22814 ( .A1(n25739), .A2(n20258), .B1(n25790), .B2(n25731), .ZN(
        n7234) );
  OAI22_X1 U22815 ( .A1(n25739), .A2(n20257), .B1(n25793), .B2(n25731), .ZN(
        n7235) );
  OAI22_X1 U22816 ( .A1(n25739), .A2(n20256), .B1(n25796), .B2(n25731), .ZN(
        n7236) );
  OAI22_X1 U22817 ( .A1(n25739), .A2(n20255), .B1(n25799), .B2(n25731), .ZN(
        n7237) );
  OAI22_X1 U22818 ( .A1(n25739), .A2(n20254), .B1(n25802), .B2(n25731), .ZN(
        n7238) );
  OAI22_X1 U22819 ( .A1(n25739), .A2(n20253), .B1(n25805), .B2(n25731), .ZN(
        n7239) );
  OAI22_X1 U22820 ( .A1(n25739), .A2(n20252), .B1(n25808), .B2(n25731), .ZN(
        n7240) );
  OAI22_X1 U22821 ( .A1(n25739), .A2(n20251), .B1(n25811), .B2(n25731), .ZN(
        n7241) );
  OAI22_X1 U22822 ( .A1(n25739), .A2(n20250), .B1(n25814), .B2(n25731), .ZN(
        n7242) );
  OAI22_X1 U22823 ( .A1(n25740), .A2(n20249), .B1(n25817), .B2(n25732), .ZN(
        n7243) );
  OAI22_X1 U22824 ( .A1(n25740), .A2(n20248), .B1(n25820), .B2(n25732), .ZN(
        n7244) );
  OAI22_X1 U22825 ( .A1(n25740), .A2(n20247), .B1(n25823), .B2(n25732), .ZN(
        n7245) );
  OAI22_X1 U22826 ( .A1(n25740), .A2(n20246), .B1(n25826), .B2(n25732), .ZN(
        n7246) );
  OAI22_X1 U22827 ( .A1(n25740), .A2(n20245), .B1(n25829), .B2(n25732), .ZN(
        n7247) );
  OAI22_X1 U22828 ( .A1(n25740), .A2(n20244), .B1(n25832), .B2(n25732), .ZN(
        n7248) );
  OAI22_X1 U22829 ( .A1(n25740), .A2(n20243), .B1(n25835), .B2(n25732), .ZN(
        n7249) );
  OAI22_X1 U22830 ( .A1(n25740), .A2(n20242), .B1(n25838), .B2(n25732), .ZN(
        n7250) );
  OAI22_X1 U22831 ( .A1(n25740), .A2(n20241), .B1(n25841), .B2(n25732), .ZN(
        n7251) );
  OAI22_X1 U22832 ( .A1(n25740), .A2(n20240), .B1(n25844), .B2(n25732), .ZN(
        n7252) );
  OAI22_X1 U22833 ( .A1(n25740), .A2(n20239), .B1(n25847), .B2(n25732), .ZN(
        n7253) );
  OAI22_X1 U22834 ( .A1(n25740), .A2(n20238), .B1(n25850), .B2(n25732), .ZN(
        n7254) );
  OAI22_X1 U22835 ( .A1(n25740), .A2(n20237), .B1(n25853), .B2(n25733), .ZN(
        n7255) );
  OAI22_X1 U22836 ( .A1(n25741), .A2(n20236), .B1(n25856), .B2(n25733), .ZN(
        n7256) );
  OAI22_X1 U22837 ( .A1(n25741), .A2(n20235), .B1(n25859), .B2(n25733), .ZN(
        n7257) );
  OAI22_X1 U22838 ( .A1(n25741), .A2(n20234), .B1(n25862), .B2(n25733), .ZN(
        n7258) );
  OAI22_X1 U22839 ( .A1(n25741), .A2(n20233), .B1(n25865), .B2(n25733), .ZN(
        n7259) );
  OAI22_X1 U22840 ( .A1(n25741), .A2(n20232), .B1(n25868), .B2(n25733), .ZN(
        n7260) );
  OAI22_X1 U22841 ( .A1(n25741), .A2(n20231), .B1(n25871), .B2(n25733), .ZN(
        n7261) );
  OAI22_X1 U22842 ( .A1(n25741), .A2(n20230), .B1(n25874), .B2(n25733), .ZN(
        n7262) );
  OAI22_X1 U22843 ( .A1(n25741), .A2(n20229), .B1(n25877), .B2(n25733), .ZN(
        n7263) );
  OAI22_X1 U22844 ( .A1(n25741), .A2(n20228), .B1(n25880), .B2(n25733), .ZN(
        n7264) );
  OAI22_X1 U22845 ( .A1(n25741), .A2(n20227), .B1(n25883), .B2(n25733), .ZN(
        n7265) );
  OAI22_X1 U22846 ( .A1(n25741), .A2(n20226), .B1(n25886), .B2(n25733), .ZN(
        n7266) );
  OAI22_X1 U22847 ( .A1(n25741), .A2(n20225), .B1(n25889), .B2(n25734), .ZN(
        n7267) );
  OAI22_X1 U22848 ( .A1(n25741), .A2(n20224), .B1(n25892), .B2(n25734), .ZN(
        n7268) );
  OAI22_X1 U22849 ( .A1(n25742), .A2(n20223), .B1(n25895), .B2(n25734), .ZN(
        n7269) );
  OAI22_X1 U22850 ( .A1(n25742), .A2(n20222), .B1(n25898), .B2(n25734), .ZN(
        n7270) );
  OAI22_X1 U22851 ( .A1(n25742), .A2(n20221), .B1(n25901), .B2(n25734), .ZN(
        n7271) );
  OAI22_X1 U22852 ( .A1(n25742), .A2(n20220), .B1(n25904), .B2(n25734), .ZN(
        n7272) );
  OAI22_X1 U22853 ( .A1(n25742), .A2(n20219), .B1(n25907), .B2(n25734), .ZN(
        n7273) );
  OAI22_X1 U22854 ( .A1(n25742), .A2(n20218), .B1(n25910), .B2(n25734), .ZN(
        n7274) );
  OAI22_X1 U22855 ( .A1(n25742), .A2(n20217), .B1(n25913), .B2(n25734), .ZN(
        n7275) );
  OAI22_X1 U22856 ( .A1(n25742), .A2(n20216), .B1(n25916), .B2(n25734), .ZN(
        n7276) );
  OAI22_X1 U22857 ( .A1(n25742), .A2(n20215), .B1(n25919), .B2(n25734), .ZN(
        n7277) );
  OAI22_X1 U22858 ( .A1(n25742), .A2(n20214), .B1(n25922), .B2(n25734), .ZN(
        n7278) );
  OAI22_X1 U22859 ( .A1(n25742), .A2(n20213), .B1(n25925), .B2(n25735), .ZN(
        n7279) );
  OAI22_X1 U22860 ( .A1(n25742), .A2(n20212), .B1(n25928), .B2(n25735), .ZN(
        n7280) );
  OAI22_X1 U22861 ( .A1(n25742), .A2(n20211), .B1(n25931), .B2(n25735), .ZN(
        n7281) );
  OAI22_X1 U22862 ( .A1(n25743), .A2(n20210), .B1(n25934), .B2(n25735), .ZN(
        n7282) );
  OAI22_X1 U22863 ( .A1(n25743), .A2(n20209), .B1(n25937), .B2(n25735), .ZN(
        n7283) );
  OAI22_X1 U22864 ( .A1(n25743), .A2(n20208), .B1(n25940), .B2(n25735), .ZN(
        n7284) );
  OAI22_X1 U22865 ( .A1(n25743), .A2(n20207), .B1(n25943), .B2(n25735), .ZN(
        n7285) );
  OAI22_X1 U22866 ( .A1(n25743), .A2(n20206), .B1(n25946), .B2(n25735), .ZN(
        n7286) );
  OAI22_X1 U22867 ( .A1(n25743), .A2(n20205), .B1(n25949), .B2(n25735), .ZN(
        n7287) );
  OAI22_X1 U22868 ( .A1(n25743), .A2(n20204), .B1(n25952), .B2(n25735), .ZN(
        n7288) );
  OAI22_X1 U22869 ( .A1(n25743), .A2(n20203), .B1(n25955), .B2(n25735), .ZN(
        n7289) );
  OAI22_X1 U22870 ( .A1(n25743), .A2(n20202), .B1(n25958), .B2(n25735), .ZN(
        n7290) );
  OAI22_X1 U22871 ( .A1(n9286), .A2(n25583), .B1(n25782), .B2(n25577), .ZN(
        n6463) );
  OAI22_X1 U22872 ( .A1(n9285), .A2(n25583), .B1(n25785), .B2(n25577), .ZN(
        n6464) );
  OAI22_X1 U22873 ( .A1(n9284), .A2(n25583), .B1(n25788), .B2(n25577), .ZN(
        n6465) );
  OAI22_X1 U22874 ( .A1(n9283), .A2(n25583), .B1(n25791), .B2(n25577), .ZN(
        n6466) );
  OAI22_X1 U22875 ( .A1(n9282), .A2(n25583), .B1(n25794), .B2(n25577), .ZN(
        n6467) );
  OAI22_X1 U22876 ( .A1(n9281), .A2(n25583), .B1(n25797), .B2(n25577), .ZN(
        n6468) );
  OAI22_X1 U22877 ( .A1(n9280), .A2(n25583), .B1(n25800), .B2(n25577), .ZN(
        n6469) );
  OAI22_X1 U22878 ( .A1(n9279), .A2(n25583), .B1(n25803), .B2(n25577), .ZN(
        n6470) );
  OAI22_X1 U22879 ( .A1(n9278), .A2(n25583), .B1(n25806), .B2(n25577), .ZN(
        n6471) );
  OAI22_X1 U22880 ( .A1(n9277), .A2(n25583), .B1(n25809), .B2(n25577), .ZN(
        n6472) );
  OAI22_X1 U22881 ( .A1(n9276), .A2(n25583), .B1(n25812), .B2(n25577), .ZN(
        n6473) );
  OAI22_X1 U22882 ( .A1(n9275), .A2(n25584), .B1(n25815), .B2(n25577), .ZN(
        n6474) );
  OAI22_X1 U22883 ( .A1(n9274), .A2(n25584), .B1(n25818), .B2(n25578), .ZN(
        n6475) );
  OAI22_X1 U22884 ( .A1(n9273), .A2(n25584), .B1(n25821), .B2(n25578), .ZN(
        n6476) );
  OAI22_X1 U22885 ( .A1(n9272), .A2(n25584), .B1(n25824), .B2(n25578), .ZN(
        n6477) );
  OAI22_X1 U22886 ( .A1(n9271), .A2(n25584), .B1(n25827), .B2(n25578), .ZN(
        n6478) );
  OAI22_X1 U22887 ( .A1(n9270), .A2(n25584), .B1(n25830), .B2(n25578), .ZN(
        n6479) );
  OAI22_X1 U22888 ( .A1(n9269), .A2(n25584), .B1(n25833), .B2(n25578), .ZN(
        n6480) );
  OAI22_X1 U22889 ( .A1(n9268), .A2(n25584), .B1(n25836), .B2(n25578), .ZN(
        n6481) );
  OAI22_X1 U22890 ( .A1(n9267), .A2(n25584), .B1(n25839), .B2(n25578), .ZN(
        n6482) );
  OAI22_X1 U22891 ( .A1(n9266), .A2(n25584), .B1(n25842), .B2(n25578), .ZN(
        n6483) );
  OAI22_X1 U22892 ( .A1(n9265), .A2(n25584), .B1(n25845), .B2(n25578), .ZN(
        n6484) );
  OAI22_X1 U22893 ( .A1(n9264), .A2(n25584), .B1(n25848), .B2(n25578), .ZN(
        n6485) );
  OAI22_X1 U22894 ( .A1(n9263), .A2(n25585), .B1(n25851), .B2(n25578), .ZN(
        n6486) );
  OAI22_X1 U22895 ( .A1(n9262), .A2(n25585), .B1(n25854), .B2(n25579), .ZN(
        n6487) );
  OAI22_X1 U22896 ( .A1(n9261), .A2(n25585), .B1(n25857), .B2(n25579), .ZN(
        n6488) );
  OAI22_X1 U22897 ( .A1(n9260), .A2(n25585), .B1(n25860), .B2(n25579), .ZN(
        n6489) );
  OAI22_X1 U22898 ( .A1(n9259), .A2(n25585), .B1(n25863), .B2(n25579), .ZN(
        n6490) );
  OAI22_X1 U22899 ( .A1(n9258), .A2(n25585), .B1(n25866), .B2(n25579), .ZN(
        n6491) );
  OAI22_X1 U22900 ( .A1(n9257), .A2(n25585), .B1(n25869), .B2(n25579), .ZN(
        n6492) );
  OAI22_X1 U22901 ( .A1(n9256), .A2(n25585), .B1(n25872), .B2(n25579), .ZN(
        n6493) );
  OAI22_X1 U22902 ( .A1(n9255), .A2(n25585), .B1(n25875), .B2(n25579), .ZN(
        n6494) );
  OAI22_X1 U22903 ( .A1(n9254), .A2(n25585), .B1(n25878), .B2(n25579), .ZN(
        n6495) );
  OAI22_X1 U22904 ( .A1(n9253), .A2(n25585), .B1(n25881), .B2(n25579), .ZN(
        n6496) );
  OAI22_X1 U22905 ( .A1(n9252), .A2(n25585), .B1(n25884), .B2(n25579), .ZN(
        n6497) );
  OAI22_X1 U22906 ( .A1(n9251), .A2(n25586), .B1(n25887), .B2(n25579), .ZN(
        n6498) );
  OAI22_X1 U22907 ( .A1(n9250), .A2(n25586), .B1(n25890), .B2(n25580), .ZN(
        n6499) );
  OAI22_X1 U22908 ( .A1(n9249), .A2(n25586), .B1(n25893), .B2(n25580), .ZN(
        n6500) );
  OAI22_X1 U22909 ( .A1(n9248), .A2(n25586), .B1(n25896), .B2(n25580), .ZN(
        n6501) );
  OAI22_X1 U22910 ( .A1(n9247), .A2(n25586), .B1(n25899), .B2(n25580), .ZN(
        n6502) );
  OAI22_X1 U22911 ( .A1(n9246), .A2(n25586), .B1(n25902), .B2(n25580), .ZN(
        n6503) );
  OAI22_X1 U22912 ( .A1(n9245), .A2(n25586), .B1(n25905), .B2(n25580), .ZN(
        n6504) );
  OAI22_X1 U22913 ( .A1(n9244), .A2(n25586), .B1(n25908), .B2(n25580), .ZN(
        n6505) );
  OAI22_X1 U22914 ( .A1(n9243), .A2(n25586), .B1(n25911), .B2(n25580), .ZN(
        n6506) );
  OAI22_X1 U22915 ( .A1(n9242), .A2(n25586), .B1(n25914), .B2(n25580), .ZN(
        n6507) );
  OAI22_X1 U22916 ( .A1(n9241), .A2(n25586), .B1(n25917), .B2(n25580), .ZN(
        n6508) );
  OAI22_X1 U22917 ( .A1(n9240), .A2(n25586), .B1(n25920), .B2(n25580), .ZN(
        n6509) );
  OAI22_X1 U22918 ( .A1(n9239), .A2(n25587), .B1(n25923), .B2(n25580), .ZN(
        n6510) );
  OAI22_X1 U22919 ( .A1(n9238), .A2(n25587), .B1(n25926), .B2(n25581), .ZN(
        n6511) );
  OAI22_X1 U22920 ( .A1(n9237), .A2(n25587), .B1(n25929), .B2(n25581), .ZN(
        n6512) );
  OAI22_X1 U22921 ( .A1(n9236), .A2(n25587), .B1(n25932), .B2(n25581), .ZN(
        n6513) );
  OAI22_X1 U22922 ( .A1(n9235), .A2(n25587), .B1(n25935), .B2(n25581), .ZN(
        n6514) );
  OAI22_X1 U22923 ( .A1(n9234), .A2(n25587), .B1(n25938), .B2(n25581), .ZN(
        n6515) );
  OAI22_X1 U22924 ( .A1(n9233), .A2(n25587), .B1(n25941), .B2(n25581), .ZN(
        n6516) );
  OAI22_X1 U22925 ( .A1(n9232), .A2(n25587), .B1(n25944), .B2(n25581), .ZN(
        n6517) );
  OAI22_X1 U22926 ( .A1(n9231), .A2(n25587), .B1(n25947), .B2(n25581), .ZN(
        n6518) );
  OAI22_X1 U22927 ( .A1(n9230), .A2(n25587), .B1(n25950), .B2(n25581), .ZN(
        n6519) );
  OAI22_X1 U22928 ( .A1(n9229), .A2(n25587), .B1(n25953), .B2(n25581), .ZN(
        n6520) );
  OAI22_X1 U22929 ( .A1(n9228), .A2(n25587), .B1(n25956), .B2(n25581), .ZN(
        n6521) );
  OAI22_X1 U22930 ( .A1(n9227), .A2(n25588), .B1(n25959), .B2(n25581), .ZN(
        n6522) );
  OAI22_X1 U22931 ( .A1(n9030), .A2(n25506), .B1(n25782), .B2(n25500), .ZN(
        n6079) );
  OAI22_X1 U22932 ( .A1(n9029), .A2(n25506), .B1(n25785), .B2(n25500), .ZN(
        n6080) );
  OAI22_X1 U22933 ( .A1(n9028), .A2(n25506), .B1(n25788), .B2(n25500), .ZN(
        n6081) );
  OAI22_X1 U22934 ( .A1(n9027), .A2(n25506), .B1(n25791), .B2(n25500), .ZN(
        n6082) );
  OAI22_X1 U22935 ( .A1(n9026), .A2(n25506), .B1(n25794), .B2(n25500), .ZN(
        n6083) );
  OAI22_X1 U22936 ( .A1(n9025), .A2(n25506), .B1(n25797), .B2(n25500), .ZN(
        n6084) );
  OAI22_X1 U22937 ( .A1(n9024), .A2(n25506), .B1(n25800), .B2(n25500), .ZN(
        n6085) );
  OAI22_X1 U22938 ( .A1(n9023), .A2(n25506), .B1(n25803), .B2(n25500), .ZN(
        n6086) );
  OAI22_X1 U22939 ( .A1(n9022), .A2(n25506), .B1(n25806), .B2(n25500), .ZN(
        n6087) );
  OAI22_X1 U22940 ( .A1(n9021), .A2(n25506), .B1(n25809), .B2(n25500), .ZN(
        n6088) );
  OAI22_X1 U22941 ( .A1(n9020), .A2(n25506), .B1(n25812), .B2(n25500), .ZN(
        n6089) );
  OAI22_X1 U22942 ( .A1(n9019), .A2(n25507), .B1(n25815), .B2(n25500), .ZN(
        n6090) );
  OAI22_X1 U22943 ( .A1(n9018), .A2(n25507), .B1(n25818), .B2(n25501), .ZN(
        n6091) );
  OAI22_X1 U22944 ( .A1(n9017), .A2(n25507), .B1(n25821), .B2(n25501), .ZN(
        n6092) );
  OAI22_X1 U22945 ( .A1(n9016), .A2(n25507), .B1(n25824), .B2(n25501), .ZN(
        n6093) );
  OAI22_X1 U22946 ( .A1(n9015), .A2(n25507), .B1(n25827), .B2(n25501), .ZN(
        n6094) );
  OAI22_X1 U22947 ( .A1(n9014), .A2(n25507), .B1(n25830), .B2(n25501), .ZN(
        n6095) );
  OAI22_X1 U22948 ( .A1(n9013), .A2(n25507), .B1(n25833), .B2(n25501), .ZN(
        n6096) );
  OAI22_X1 U22949 ( .A1(n9012), .A2(n25507), .B1(n25836), .B2(n25501), .ZN(
        n6097) );
  OAI22_X1 U22950 ( .A1(n9011), .A2(n25507), .B1(n25839), .B2(n25501), .ZN(
        n6098) );
  OAI22_X1 U22951 ( .A1(n9010), .A2(n25507), .B1(n25842), .B2(n25501), .ZN(
        n6099) );
  OAI22_X1 U22952 ( .A1(n9009), .A2(n25507), .B1(n25845), .B2(n25501), .ZN(
        n6100) );
  OAI22_X1 U22953 ( .A1(n9008), .A2(n25507), .B1(n25848), .B2(n25501), .ZN(
        n6101) );
  OAI22_X1 U22954 ( .A1(n9007), .A2(n25508), .B1(n25851), .B2(n25501), .ZN(
        n6102) );
  OAI22_X1 U22955 ( .A1(n9006), .A2(n25508), .B1(n25854), .B2(n25502), .ZN(
        n6103) );
  OAI22_X1 U22956 ( .A1(n9005), .A2(n25508), .B1(n25857), .B2(n25502), .ZN(
        n6104) );
  OAI22_X1 U22957 ( .A1(n9004), .A2(n25508), .B1(n25860), .B2(n25502), .ZN(
        n6105) );
  OAI22_X1 U22958 ( .A1(n9003), .A2(n25508), .B1(n25863), .B2(n25502), .ZN(
        n6106) );
  OAI22_X1 U22959 ( .A1(n9002), .A2(n25508), .B1(n25866), .B2(n25502), .ZN(
        n6107) );
  OAI22_X1 U22960 ( .A1(n9001), .A2(n25508), .B1(n25869), .B2(n25502), .ZN(
        n6108) );
  OAI22_X1 U22961 ( .A1(n9000), .A2(n25508), .B1(n25872), .B2(n25502), .ZN(
        n6109) );
  OAI22_X1 U22962 ( .A1(n8999), .A2(n25508), .B1(n25875), .B2(n25502), .ZN(
        n6110) );
  OAI22_X1 U22963 ( .A1(n8998), .A2(n25508), .B1(n25878), .B2(n25502), .ZN(
        n6111) );
  OAI22_X1 U22964 ( .A1(n8997), .A2(n25508), .B1(n25881), .B2(n25502), .ZN(
        n6112) );
  OAI22_X1 U22965 ( .A1(n8996), .A2(n25508), .B1(n25884), .B2(n25502), .ZN(
        n6113) );
  OAI22_X1 U22966 ( .A1(n8995), .A2(n25509), .B1(n25887), .B2(n25502), .ZN(
        n6114) );
  OAI22_X1 U22967 ( .A1(n8994), .A2(n25509), .B1(n25890), .B2(n25503), .ZN(
        n6115) );
  OAI22_X1 U22968 ( .A1(n8993), .A2(n25509), .B1(n25893), .B2(n25503), .ZN(
        n6116) );
  OAI22_X1 U22969 ( .A1(n8992), .A2(n25509), .B1(n25896), .B2(n25503), .ZN(
        n6117) );
  OAI22_X1 U22970 ( .A1(n8991), .A2(n25509), .B1(n25899), .B2(n25503), .ZN(
        n6118) );
  OAI22_X1 U22971 ( .A1(n8990), .A2(n25509), .B1(n25902), .B2(n25503), .ZN(
        n6119) );
  OAI22_X1 U22972 ( .A1(n8989), .A2(n25509), .B1(n25905), .B2(n25503), .ZN(
        n6120) );
  OAI22_X1 U22973 ( .A1(n8988), .A2(n25509), .B1(n25908), .B2(n25503), .ZN(
        n6121) );
  OAI22_X1 U22974 ( .A1(n8987), .A2(n25509), .B1(n25911), .B2(n25503), .ZN(
        n6122) );
  OAI22_X1 U22975 ( .A1(n8986), .A2(n25509), .B1(n25914), .B2(n25503), .ZN(
        n6123) );
  OAI22_X1 U22976 ( .A1(n8985), .A2(n25509), .B1(n25917), .B2(n25503), .ZN(
        n6124) );
  OAI22_X1 U22977 ( .A1(n8984), .A2(n25509), .B1(n25920), .B2(n25503), .ZN(
        n6125) );
  OAI22_X1 U22978 ( .A1(n8983), .A2(n25510), .B1(n25923), .B2(n25503), .ZN(
        n6126) );
  OAI22_X1 U22979 ( .A1(n8982), .A2(n25510), .B1(n25926), .B2(n25504), .ZN(
        n6127) );
  OAI22_X1 U22980 ( .A1(n8981), .A2(n25510), .B1(n25929), .B2(n25504), .ZN(
        n6128) );
  OAI22_X1 U22981 ( .A1(n8980), .A2(n25510), .B1(n25932), .B2(n25504), .ZN(
        n6129) );
  OAI22_X1 U22982 ( .A1(n8979), .A2(n25510), .B1(n25935), .B2(n25504), .ZN(
        n6130) );
  OAI22_X1 U22983 ( .A1(n8978), .A2(n25510), .B1(n25938), .B2(n25504), .ZN(
        n6131) );
  OAI22_X1 U22984 ( .A1(n8977), .A2(n25510), .B1(n25941), .B2(n25504), .ZN(
        n6132) );
  OAI22_X1 U22985 ( .A1(n8976), .A2(n25510), .B1(n25944), .B2(n25504), .ZN(
        n6133) );
  OAI22_X1 U22986 ( .A1(n8975), .A2(n25510), .B1(n25947), .B2(n25504), .ZN(
        n6134) );
  OAI22_X1 U22987 ( .A1(n8974), .A2(n25510), .B1(n25950), .B2(n25504), .ZN(
        n6135) );
  OAI22_X1 U22988 ( .A1(n8973), .A2(n25510), .B1(n25953), .B2(n25504), .ZN(
        n6136) );
  OAI22_X1 U22989 ( .A1(n8972), .A2(n25510), .B1(n25956), .B2(n25504), .ZN(
        n6137) );
  OAI22_X1 U22990 ( .A1(n8971), .A2(n25511), .B1(n25959), .B2(n25504), .ZN(
        n6138) );
  OAI22_X1 U22991 ( .A1(n9478), .A2(n25775), .B1(n25769), .B2(n25781), .ZN(
        n7423) );
  OAI22_X1 U22992 ( .A1(n9477), .A2(n25775), .B1(n25769), .B2(n25784), .ZN(
        n7424) );
  OAI22_X1 U22993 ( .A1(n9476), .A2(n25775), .B1(n25769), .B2(n25787), .ZN(
        n7425) );
  OAI22_X1 U22994 ( .A1(n9475), .A2(n25775), .B1(n25769), .B2(n25790), .ZN(
        n7426) );
  OAI22_X1 U22995 ( .A1(n9474), .A2(n25775), .B1(n25769), .B2(n25793), .ZN(
        n7427) );
  OAI22_X1 U22996 ( .A1(n9473), .A2(n25775), .B1(n25769), .B2(n25796), .ZN(
        n7428) );
  OAI22_X1 U22997 ( .A1(n9472), .A2(n25775), .B1(n25769), .B2(n25799), .ZN(
        n7429) );
  OAI22_X1 U22998 ( .A1(n9471), .A2(n25775), .B1(n25769), .B2(n25802), .ZN(
        n7430) );
  OAI22_X1 U22999 ( .A1(n9470), .A2(n25775), .B1(n25769), .B2(n25805), .ZN(
        n7431) );
  OAI22_X1 U23000 ( .A1(n9469), .A2(n25775), .B1(n25769), .B2(n25808), .ZN(
        n7432) );
  OAI22_X1 U23001 ( .A1(n9468), .A2(n25775), .B1(n25769), .B2(n25811), .ZN(
        n7433) );
  OAI22_X1 U23002 ( .A1(n9467), .A2(n25776), .B1(n25769), .B2(n25814), .ZN(
        n7434) );
  OAI22_X1 U23003 ( .A1(n9094), .A2(n25750), .B1(n25781), .B2(n25744), .ZN(
        n7295) );
  OAI22_X1 U23004 ( .A1(n9093), .A2(n25750), .B1(n25784), .B2(n25744), .ZN(
        n7296) );
  OAI22_X1 U23005 ( .A1(n9092), .A2(n25750), .B1(n25787), .B2(n25744), .ZN(
        n7297) );
  OAI22_X1 U23006 ( .A1(n9091), .A2(n25750), .B1(n25790), .B2(n25744), .ZN(
        n7298) );
  OAI22_X1 U23007 ( .A1(n9090), .A2(n25750), .B1(n25793), .B2(n25744), .ZN(
        n7299) );
  OAI22_X1 U23008 ( .A1(n9089), .A2(n25750), .B1(n25796), .B2(n25744), .ZN(
        n7300) );
  OAI22_X1 U23009 ( .A1(n9088), .A2(n25750), .B1(n25799), .B2(n25744), .ZN(
        n7301) );
  OAI22_X1 U23010 ( .A1(n9087), .A2(n25750), .B1(n25802), .B2(n25744), .ZN(
        n7302) );
  OAI22_X1 U23011 ( .A1(n9086), .A2(n25750), .B1(n25805), .B2(n25744), .ZN(
        n7303) );
  OAI22_X1 U23012 ( .A1(n9085), .A2(n25750), .B1(n25808), .B2(n25744), .ZN(
        n7304) );
  OAI22_X1 U23013 ( .A1(n9084), .A2(n25750), .B1(n25811), .B2(n25744), .ZN(
        n7305) );
  OAI22_X1 U23014 ( .A1(n9083), .A2(n25751), .B1(n25814), .B2(n25744), .ZN(
        n7306) );
  OAI22_X1 U23015 ( .A1(n9082), .A2(n25751), .B1(n25817), .B2(n25745), .ZN(
        n7307) );
  OAI22_X1 U23016 ( .A1(n9081), .A2(n25751), .B1(n25820), .B2(n25745), .ZN(
        n7308) );
  OAI22_X1 U23017 ( .A1(n9080), .A2(n25751), .B1(n25823), .B2(n25745), .ZN(
        n7309) );
  OAI22_X1 U23018 ( .A1(n9079), .A2(n25751), .B1(n25826), .B2(n25745), .ZN(
        n7310) );
  OAI22_X1 U23019 ( .A1(n9078), .A2(n25751), .B1(n25829), .B2(n25745), .ZN(
        n7311) );
  OAI22_X1 U23020 ( .A1(n9077), .A2(n25751), .B1(n25832), .B2(n25745), .ZN(
        n7312) );
  OAI22_X1 U23021 ( .A1(n9076), .A2(n25751), .B1(n25835), .B2(n25745), .ZN(
        n7313) );
  OAI22_X1 U23022 ( .A1(n9075), .A2(n25751), .B1(n25838), .B2(n25745), .ZN(
        n7314) );
  OAI22_X1 U23023 ( .A1(n9074), .A2(n25751), .B1(n25841), .B2(n25745), .ZN(
        n7315) );
  OAI22_X1 U23024 ( .A1(n9073), .A2(n25751), .B1(n25844), .B2(n25745), .ZN(
        n7316) );
  OAI22_X1 U23025 ( .A1(n9072), .A2(n25751), .B1(n25847), .B2(n25745), .ZN(
        n7317) );
  OAI22_X1 U23026 ( .A1(n9071), .A2(n25752), .B1(n25850), .B2(n25745), .ZN(
        n7318) );
  OAI22_X1 U23027 ( .A1(n9070), .A2(n25752), .B1(n25853), .B2(n25746), .ZN(
        n7319) );
  OAI22_X1 U23028 ( .A1(n9069), .A2(n25752), .B1(n25856), .B2(n25746), .ZN(
        n7320) );
  OAI22_X1 U23029 ( .A1(n9068), .A2(n25752), .B1(n25859), .B2(n25746), .ZN(
        n7321) );
  OAI22_X1 U23030 ( .A1(n9067), .A2(n25752), .B1(n25862), .B2(n25746), .ZN(
        n7322) );
  OAI22_X1 U23031 ( .A1(n9066), .A2(n25752), .B1(n25865), .B2(n25746), .ZN(
        n7323) );
  OAI22_X1 U23032 ( .A1(n9065), .A2(n25752), .B1(n25868), .B2(n25746), .ZN(
        n7324) );
  OAI22_X1 U23033 ( .A1(n9064), .A2(n25752), .B1(n25871), .B2(n25746), .ZN(
        n7325) );
  OAI22_X1 U23034 ( .A1(n9063), .A2(n25752), .B1(n25874), .B2(n25746), .ZN(
        n7326) );
  OAI22_X1 U23035 ( .A1(n9062), .A2(n25752), .B1(n25877), .B2(n25746), .ZN(
        n7327) );
  OAI22_X1 U23036 ( .A1(n9061), .A2(n25752), .B1(n25880), .B2(n25746), .ZN(
        n7328) );
  OAI22_X1 U23037 ( .A1(n9060), .A2(n25752), .B1(n25883), .B2(n25746), .ZN(
        n7329) );
  OAI22_X1 U23038 ( .A1(n9059), .A2(n25753), .B1(n25886), .B2(n25746), .ZN(
        n7330) );
  OAI22_X1 U23039 ( .A1(n9058), .A2(n25753), .B1(n25889), .B2(n25747), .ZN(
        n7331) );
  OAI22_X1 U23040 ( .A1(n9057), .A2(n25753), .B1(n25892), .B2(n25747), .ZN(
        n7332) );
  OAI22_X1 U23041 ( .A1(n9056), .A2(n25753), .B1(n25895), .B2(n25747), .ZN(
        n7333) );
  OAI22_X1 U23042 ( .A1(n9055), .A2(n25753), .B1(n25898), .B2(n25747), .ZN(
        n7334) );
  OAI22_X1 U23043 ( .A1(n9054), .A2(n25753), .B1(n25901), .B2(n25747), .ZN(
        n7335) );
  OAI22_X1 U23044 ( .A1(n9053), .A2(n25753), .B1(n25904), .B2(n25747), .ZN(
        n7336) );
  OAI22_X1 U23045 ( .A1(n9052), .A2(n25753), .B1(n25907), .B2(n25747), .ZN(
        n7337) );
  OAI22_X1 U23046 ( .A1(n9051), .A2(n25753), .B1(n25910), .B2(n25747), .ZN(
        n7338) );
  OAI22_X1 U23047 ( .A1(n9050), .A2(n25753), .B1(n25913), .B2(n25747), .ZN(
        n7339) );
  OAI22_X1 U23048 ( .A1(n9049), .A2(n25753), .B1(n25916), .B2(n25747), .ZN(
        n7340) );
  OAI22_X1 U23049 ( .A1(n9048), .A2(n25753), .B1(n25919), .B2(n25747), .ZN(
        n7341) );
  OAI22_X1 U23050 ( .A1(n9047), .A2(n25754), .B1(n25922), .B2(n25747), .ZN(
        n7342) );
  OAI22_X1 U23051 ( .A1(n9046), .A2(n25754), .B1(n25925), .B2(n25748), .ZN(
        n7343) );
  OAI22_X1 U23052 ( .A1(n9045), .A2(n25754), .B1(n25928), .B2(n25748), .ZN(
        n7344) );
  OAI22_X1 U23053 ( .A1(n9044), .A2(n25754), .B1(n25931), .B2(n25748), .ZN(
        n7345) );
  OAI22_X1 U23054 ( .A1(n9043), .A2(n25754), .B1(n25934), .B2(n25748), .ZN(
        n7346) );
  OAI22_X1 U23055 ( .A1(n9042), .A2(n25754), .B1(n25937), .B2(n25748), .ZN(
        n7347) );
  OAI22_X1 U23056 ( .A1(n9041), .A2(n25754), .B1(n25940), .B2(n25748), .ZN(
        n7348) );
  OAI22_X1 U23057 ( .A1(n9040), .A2(n25754), .B1(n25943), .B2(n25748), .ZN(
        n7349) );
  OAI22_X1 U23058 ( .A1(n9039), .A2(n25754), .B1(n25946), .B2(n25748), .ZN(
        n7350) );
  OAI22_X1 U23059 ( .A1(n9038), .A2(n25754), .B1(n25949), .B2(n25748), .ZN(
        n7351) );
  OAI22_X1 U23060 ( .A1(n9037), .A2(n25754), .B1(n25952), .B2(n25748), .ZN(
        n7352) );
  OAI22_X1 U23061 ( .A1(n9036), .A2(n25754), .B1(n25955), .B2(n25748), .ZN(
        n7353) );
  OAI22_X1 U23062 ( .A1(n9035), .A2(n25755), .B1(n25958), .B2(n25748), .ZN(
        n7354) );
  OAI22_X1 U23063 ( .A1(n9350), .A2(n25686), .B1(n25781), .B2(n25680), .ZN(
        n6975) );
  OAI22_X1 U23064 ( .A1(n9349), .A2(n25686), .B1(n25784), .B2(n25680), .ZN(
        n6976) );
  OAI22_X1 U23065 ( .A1(n9348), .A2(n25686), .B1(n25787), .B2(n25680), .ZN(
        n6977) );
  OAI22_X1 U23066 ( .A1(n9347), .A2(n25686), .B1(n25790), .B2(n25680), .ZN(
        n6978) );
  OAI22_X1 U23067 ( .A1(n9346), .A2(n25686), .B1(n25793), .B2(n25680), .ZN(
        n6979) );
  OAI22_X1 U23068 ( .A1(n9345), .A2(n25686), .B1(n25796), .B2(n25680), .ZN(
        n6980) );
  OAI22_X1 U23069 ( .A1(n9344), .A2(n25686), .B1(n25799), .B2(n25680), .ZN(
        n6981) );
  OAI22_X1 U23070 ( .A1(n9343), .A2(n25686), .B1(n25802), .B2(n25680), .ZN(
        n6982) );
  OAI22_X1 U23071 ( .A1(n9342), .A2(n25686), .B1(n25805), .B2(n25680), .ZN(
        n6983) );
  OAI22_X1 U23072 ( .A1(n9341), .A2(n25686), .B1(n25808), .B2(n25680), .ZN(
        n6984) );
  OAI22_X1 U23073 ( .A1(n9340), .A2(n25686), .B1(n25811), .B2(n25680), .ZN(
        n6985) );
  OAI22_X1 U23074 ( .A1(n9339), .A2(n25687), .B1(n25814), .B2(n25680), .ZN(
        n6986) );
  OAI22_X1 U23075 ( .A1(n9338), .A2(n25687), .B1(n25817), .B2(n25681), .ZN(
        n6987) );
  OAI22_X1 U23076 ( .A1(n9337), .A2(n25687), .B1(n25820), .B2(n25681), .ZN(
        n6988) );
  OAI22_X1 U23077 ( .A1(n9336), .A2(n25687), .B1(n25823), .B2(n25681), .ZN(
        n6989) );
  OAI22_X1 U23078 ( .A1(n9335), .A2(n25687), .B1(n25826), .B2(n25681), .ZN(
        n6990) );
  OAI22_X1 U23079 ( .A1(n9334), .A2(n25687), .B1(n25829), .B2(n25681), .ZN(
        n6991) );
  OAI22_X1 U23080 ( .A1(n9333), .A2(n25687), .B1(n25832), .B2(n25681), .ZN(
        n6992) );
  OAI22_X1 U23081 ( .A1(n9332), .A2(n25687), .B1(n25835), .B2(n25681), .ZN(
        n6993) );
  OAI22_X1 U23082 ( .A1(n9331), .A2(n25687), .B1(n25838), .B2(n25681), .ZN(
        n6994) );
  OAI22_X1 U23083 ( .A1(n9330), .A2(n25687), .B1(n25841), .B2(n25681), .ZN(
        n6995) );
  OAI22_X1 U23084 ( .A1(n9329), .A2(n25687), .B1(n25844), .B2(n25681), .ZN(
        n6996) );
  OAI22_X1 U23085 ( .A1(n9328), .A2(n25687), .B1(n25847), .B2(n25681), .ZN(
        n6997) );
  OAI22_X1 U23086 ( .A1(n9327), .A2(n25688), .B1(n25850), .B2(n25681), .ZN(
        n6998) );
  OAI22_X1 U23087 ( .A1(n9326), .A2(n25688), .B1(n25853), .B2(n25682), .ZN(
        n6999) );
  OAI22_X1 U23088 ( .A1(n9325), .A2(n25688), .B1(n25856), .B2(n25682), .ZN(
        n7000) );
  OAI22_X1 U23089 ( .A1(n9324), .A2(n25688), .B1(n25859), .B2(n25682), .ZN(
        n7001) );
  OAI22_X1 U23090 ( .A1(n9323), .A2(n25688), .B1(n25862), .B2(n25682), .ZN(
        n7002) );
  OAI22_X1 U23091 ( .A1(n9322), .A2(n25688), .B1(n25865), .B2(n25682), .ZN(
        n7003) );
  OAI22_X1 U23092 ( .A1(n9321), .A2(n25688), .B1(n25868), .B2(n25682), .ZN(
        n7004) );
  OAI22_X1 U23093 ( .A1(n9320), .A2(n25688), .B1(n25871), .B2(n25682), .ZN(
        n7005) );
  OAI22_X1 U23094 ( .A1(n9319), .A2(n25688), .B1(n25874), .B2(n25682), .ZN(
        n7006) );
  OAI22_X1 U23095 ( .A1(n9318), .A2(n25688), .B1(n25877), .B2(n25682), .ZN(
        n7007) );
  OAI22_X1 U23096 ( .A1(n9317), .A2(n25688), .B1(n25880), .B2(n25682), .ZN(
        n7008) );
  OAI22_X1 U23097 ( .A1(n9316), .A2(n25688), .B1(n25883), .B2(n25682), .ZN(
        n7009) );
  OAI22_X1 U23098 ( .A1(n9315), .A2(n25689), .B1(n25886), .B2(n25682), .ZN(
        n7010) );
  OAI22_X1 U23099 ( .A1(n9314), .A2(n25689), .B1(n25889), .B2(n25683), .ZN(
        n7011) );
  OAI22_X1 U23100 ( .A1(n9313), .A2(n25689), .B1(n25892), .B2(n25683), .ZN(
        n7012) );
  OAI22_X1 U23101 ( .A1(n9312), .A2(n25689), .B1(n25895), .B2(n25683), .ZN(
        n7013) );
  OAI22_X1 U23102 ( .A1(n9311), .A2(n25689), .B1(n25898), .B2(n25683), .ZN(
        n7014) );
  OAI22_X1 U23103 ( .A1(n9310), .A2(n25689), .B1(n25901), .B2(n25683), .ZN(
        n7015) );
  OAI22_X1 U23104 ( .A1(n9309), .A2(n25689), .B1(n25904), .B2(n25683), .ZN(
        n7016) );
  OAI22_X1 U23105 ( .A1(n9308), .A2(n25689), .B1(n25907), .B2(n25683), .ZN(
        n7017) );
  OAI22_X1 U23106 ( .A1(n9307), .A2(n25689), .B1(n25910), .B2(n25683), .ZN(
        n7018) );
  OAI22_X1 U23107 ( .A1(n9306), .A2(n25689), .B1(n25913), .B2(n25683), .ZN(
        n7019) );
  OAI22_X1 U23108 ( .A1(n9305), .A2(n25689), .B1(n25916), .B2(n25683), .ZN(
        n7020) );
  OAI22_X1 U23109 ( .A1(n9304), .A2(n25689), .B1(n25919), .B2(n25683), .ZN(
        n7021) );
  OAI22_X1 U23110 ( .A1(n9303), .A2(n25690), .B1(n25922), .B2(n25683), .ZN(
        n7022) );
  OAI22_X1 U23111 ( .A1(n9302), .A2(n25690), .B1(n25925), .B2(n25684), .ZN(
        n7023) );
  OAI22_X1 U23112 ( .A1(n9301), .A2(n25690), .B1(n25928), .B2(n25684), .ZN(
        n7024) );
  OAI22_X1 U23113 ( .A1(n9300), .A2(n25690), .B1(n25931), .B2(n25684), .ZN(
        n7025) );
  OAI22_X1 U23114 ( .A1(n9299), .A2(n25690), .B1(n25934), .B2(n25684), .ZN(
        n7026) );
  OAI22_X1 U23115 ( .A1(n9298), .A2(n25690), .B1(n25937), .B2(n25684), .ZN(
        n7027) );
  OAI22_X1 U23116 ( .A1(n9297), .A2(n25690), .B1(n25940), .B2(n25684), .ZN(
        n7028) );
  OAI22_X1 U23117 ( .A1(n9296), .A2(n25690), .B1(n25943), .B2(n25684), .ZN(
        n7029) );
  OAI22_X1 U23118 ( .A1(n9295), .A2(n25690), .B1(n25946), .B2(n25684), .ZN(
        n7030) );
  OAI22_X1 U23119 ( .A1(n9294), .A2(n25690), .B1(n25949), .B2(n25684), .ZN(
        n7031) );
  OAI22_X1 U23120 ( .A1(n9293), .A2(n25690), .B1(n25952), .B2(n25684), .ZN(
        n7032) );
  OAI22_X1 U23121 ( .A1(n9292), .A2(n25690), .B1(n25955), .B2(n25684), .ZN(
        n7033) );
  OAI22_X1 U23122 ( .A1(n9291), .A2(n25691), .B1(n25958), .B2(n25684), .ZN(
        n7034) );
  OAI22_X1 U23123 ( .A1(n25495), .A2(n19940), .B1(n25782), .B2(n25487), .ZN(
        n6015) );
  OAI22_X1 U23124 ( .A1(n25495), .A2(n19939), .B1(n25785), .B2(n25487), .ZN(
        n6016) );
  OAI22_X1 U23125 ( .A1(n25495), .A2(n19938), .B1(n25788), .B2(n25487), .ZN(
        n6017) );
  OAI22_X1 U23126 ( .A1(n25495), .A2(n19937), .B1(n25791), .B2(n25487), .ZN(
        n6018) );
  OAI22_X1 U23127 ( .A1(n25495), .A2(n19936), .B1(n25794), .B2(n25487), .ZN(
        n6019) );
  OAI22_X1 U23128 ( .A1(n25495), .A2(n19935), .B1(n25797), .B2(n25487), .ZN(
        n6020) );
  OAI22_X1 U23129 ( .A1(n25495), .A2(n19934), .B1(n25800), .B2(n25487), .ZN(
        n6021) );
  OAI22_X1 U23130 ( .A1(n25495), .A2(n19933), .B1(n25803), .B2(n25487), .ZN(
        n6022) );
  OAI22_X1 U23131 ( .A1(n25495), .A2(n19932), .B1(n25806), .B2(n25487), .ZN(
        n6023) );
  OAI22_X1 U23132 ( .A1(n25495), .A2(n19931), .B1(n25809), .B2(n25487), .ZN(
        n6024) );
  OAI22_X1 U23133 ( .A1(n25495), .A2(n19930), .B1(n25812), .B2(n25487), .ZN(
        n6025) );
  OAI22_X1 U23134 ( .A1(n25495), .A2(n19929), .B1(n25815), .B2(n25487), .ZN(
        n6026) );
  OAI22_X1 U23135 ( .A1(n25496), .A2(n19928), .B1(n25818), .B2(n25488), .ZN(
        n6027) );
  OAI22_X1 U23136 ( .A1(n25496), .A2(n19927), .B1(n25821), .B2(n25488), .ZN(
        n6028) );
  OAI22_X1 U23137 ( .A1(n25496), .A2(n19926), .B1(n25824), .B2(n25488), .ZN(
        n6029) );
  OAI22_X1 U23138 ( .A1(n25496), .A2(n19925), .B1(n25827), .B2(n25488), .ZN(
        n6030) );
  OAI22_X1 U23139 ( .A1(n25496), .A2(n19924), .B1(n25830), .B2(n25488), .ZN(
        n6031) );
  OAI22_X1 U23140 ( .A1(n25496), .A2(n19923), .B1(n25833), .B2(n25488), .ZN(
        n6032) );
  OAI22_X1 U23141 ( .A1(n25496), .A2(n19922), .B1(n25836), .B2(n25488), .ZN(
        n6033) );
  OAI22_X1 U23142 ( .A1(n25496), .A2(n19921), .B1(n25839), .B2(n25488), .ZN(
        n6034) );
  OAI22_X1 U23143 ( .A1(n25496), .A2(n19920), .B1(n25842), .B2(n25488), .ZN(
        n6035) );
  OAI22_X1 U23144 ( .A1(n25496), .A2(n19919), .B1(n25845), .B2(n25488), .ZN(
        n6036) );
  OAI22_X1 U23145 ( .A1(n25496), .A2(n19918), .B1(n25848), .B2(n25488), .ZN(
        n6037) );
  OAI22_X1 U23146 ( .A1(n25496), .A2(n19917), .B1(n25851), .B2(n25488), .ZN(
        n6038) );
  OAI22_X1 U23147 ( .A1(n25496), .A2(n19916), .B1(n25854), .B2(n25489), .ZN(
        n6039) );
  OAI22_X1 U23148 ( .A1(n25497), .A2(n19915), .B1(n25857), .B2(n25489), .ZN(
        n6040) );
  OAI22_X1 U23149 ( .A1(n25497), .A2(n19914), .B1(n25860), .B2(n25489), .ZN(
        n6041) );
  OAI22_X1 U23150 ( .A1(n25497), .A2(n19913), .B1(n25863), .B2(n25489), .ZN(
        n6042) );
  OAI22_X1 U23151 ( .A1(n25497), .A2(n19912), .B1(n25866), .B2(n25489), .ZN(
        n6043) );
  OAI22_X1 U23152 ( .A1(n25497), .A2(n19911), .B1(n25869), .B2(n25489), .ZN(
        n6044) );
  OAI22_X1 U23153 ( .A1(n25497), .A2(n19910), .B1(n25872), .B2(n25489), .ZN(
        n6045) );
  OAI22_X1 U23154 ( .A1(n25497), .A2(n19909), .B1(n25875), .B2(n25489), .ZN(
        n6046) );
  OAI22_X1 U23155 ( .A1(n25497), .A2(n19908), .B1(n25878), .B2(n25489), .ZN(
        n6047) );
  OAI22_X1 U23156 ( .A1(n25497), .A2(n19907), .B1(n25881), .B2(n25489), .ZN(
        n6048) );
  OAI22_X1 U23157 ( .A1(n25497), .A2(n19906), .B1(n25884), .B2(n25489), .ZN(
        n6049) );
  OAI22_X1 U23158 ( .A1(n25497), .A2(n19905), .B1(n25887), .B2(n25489), .ZN(
        n6050) );
  OAI22_X1 U23159 ( .A1(n25497), .A2(n19904), .B1(n25890), .B2(n25490), .ZN(
        n6051) );
  OAI22_X1 U23160 ( .A1(n25497), .A2(n19903), .B1(n25893), .B2(n25490), .ZN(
        n6052) );
  OAI22_X1 U23161 ( .A1(n25498), .A2(n19902), .B1(n25896), .B2(n25490), .ZN(
        n6053) );
  OAI22_X1 U23162 ( .A1(n25498), .A2(n19901), .B1(n25899), .B2(n25490), .ZN(
        n6054) );
  OAI22_X1 U23163 ( .A1(n25498), .A2(n19900), .B1(n25902), .B2(n25490), .ZN(
        n6055) );
  OAI22_X1 U23164 ( .A1(n25498), .A2(n19899), .B1(n25905), .B2(n25490), .ZN(
        n6056) );
  OAI22_X1 U23165 ( .A1(n25498), .A2(n19898), .B1(n25908), .B2(n25490), .ZN(
        n6057) );
  OAI22_X1 U23166 ( .A1(n25498), .A2(n19897), .B1(n25911), .B2(n25490), .ZN(
        n6058) );
  OAI22_X1 U23167 ( .A1(n25498), .A2(n19896), .B1(n25914), .B2(n25490), .ZN(
        n6059) );
  OAI22_X1 U23168 ( .A1(n25498), .A2(n19895), .B1(n25917), .B2(n25490), .ZN(
        n6060) );
  OAI22_X1 U23169 ( .A1(n25498), .A2(n19894), .B1(n25920), .B2(n25490), .ZN(
        n6061) );
  OAI22_X1 U23170 ( .A1(n25498), .A2(n19893), .B1(n25923), .B2(n25490), .ZN(
        n6062) );
  OAI22_X1 U23171 ( .A1(n25498), .A2(n19892), .B1(n25926), .B2(n25491), .ZN(
        n6063) );
  OAI22_X1 U23172 ( .A1(n25498), .A2(n19891), .B1(n25929), .B2(n25491), .ZN(
        n6064) );
  OAI22_X1 U23173 ( .A1(n25498), .A2(n19890), .B1(n25932), .B2(n25491), .ZN(
        n6065) );
  OAI22_X1 U23174 ( .A1(n25499), .A2(n19889), .B1(n25935), .B2(n25491), .ZN(
        n6066) );
  OAI22_X1 U23175 ( .A1(n25499), .A2(n19888), .B1(n25938), .B2(n25491), .ZN(
        n6067) );
  OAI22_X1 U23176 ( .A1(n25499), .A2(n19887), .B1(n25941), .B2(n25491), .ZN(
        n6068) );
  OAI22_X1 U23177 ( .A1(n25499), .A2(n19886), .B1(n25944), .B2(n25491), .ZN(
        n6069) );
  OAI22_X1 U23178 ( .A1(n25499), .A2(n19885), .B1(n25947), .B2(n25491), .ZN(
        n6070) );
  OAI22_X1 U23179 ( .A1(n25499), .A2(n19884), .B1(n25950), .B2(n25491), .ZN(
        n6071) );
  OAI22_X1 U23180 ( .A1(n25499), .A2(n19883), .B1(n25953), .B2(n25491), .ZN(
        n6072) );
  OAI22_X1 U23181 ( .A1(n25499), .A2(n19882), .B1(n25956), .B2(n25491), .ZN(
        n6073) );
  OAI22_X1 U23182 ( .A1(n25499), .A2(n19881), .B1(n25959), .B2(n25491), .ZN(
        n6074) );
  OAI22_X1 U23183 ( .A1(n25700), .A2(n19685), .B1(n25781), .B2(n25692), .ZN(
        n7039) );
  OAI22_X1 U23184 ( .A1(n25700), .A2(n19684), .B1(n25784), .B2(n25692), .ZN(
        n7040) );
  OAI22_X1 U23185 ( .A1(n25700), .A2(n19683), .B1(n25787), .B2(n25692), .ZN(
        n7041) );
  OAI22_X1 U23186 ( .A1(n25700), .A2(n19682), .B1(n25790), .B2(n25692), .ZN(
        n7042) );
  OAI22_X1 U23187 ( .A1(n25700), .A2(n19681), .B1(n25793), .B2(n25692), .ZN(
        n7043) );
  OAI22_X1 U23188 ( .A1(n25700), .A2(n19680), .B1(n25796), .B2(n25692), .ZN(
        n7044) );
  OAI22_X1 U23189 ( .A1(n25700), .A2(n19679), .B1(n25799), .B2(n25692), .ZN(
        n7045) );
  OAI22_X1 U23190 ( .A1(n25700), .A2(n19678), .B1(n25802), .B2(n25692), .ZN(
        n7046) );
  OAI22_X1 U23191 ( .A1(n25700), .A2(n19677), .B1(n25805), .B2(n25692), .ZN(
        n7047) );
  OAI22_X1 U23192 ( .A1(n25700), .A2(n19676), .B1(n25808), .B2(n25692), .ZN(
        n7048) );
  OAI22_X1 U23193 ( .A1(n25700), .A2(n19675), .B1(n25811), .B2(n25692), .ZN(
        n7049) );
  OAI22_X1 U23194 ( .A1(n25700), .A2(n19674), .B1(n25814), .B2(n25692), .ZN(
        n7050) );
  OAI22_X1 U23195 ( .A1(n25701), .A2(n19673), .B1(n25817), .B2(n25693), .ZN(
        n7051) );
  OAI22_X1 U23196 ( .A1(n25701), .A2(n19672), .B1(n25820), .B2(n25693), .ZN(
        n7052) );
  OAI22_X1 U23197 ( .A1(n25701), .A2(n19671), .B1(n25823), .B2(n25693), .ZN(
        n7053) );
  OAI22_X1 U23198 ( .A1(n25701), .A2(n19670), .B1(n25826), .B2(n25693), .ZN(
        n7054) );
  OAI22_X1 U23199 ( .A1(n25701), .A2(n19669), .B1(n25829), .B2(n25693), .ZN(
        n7055) );
  OAI22_X1 U23200 ( .A1(n25701), .A2(n19668), .B1(n25832), .B2(n25693), .ZN(
        n7056) );
  OAI22_X1 U23201 ( .A1(n25701), .A2(n19667), .B1(n25835), .B2(n25693), .ZN(
        n7057) );
  OAI22_X1 U23202 ( .A1(n25701), .A2(n19666), .B1(n25838), .B2(n25693), .ZN(
        n7058) );
  OAI22_X1 U23203 ( .A1(n25701), .A2(n19665), .B1(n25841), .B2(n25693), .ZN(
        n7059) );
  OAI22_X1 U23204 ( .A1(n25701), .A2(n19664), .B1(n25844), .B2(n25693), .ZN(
        n7060) );
  OAI22_X1 U23205 ( .A1(n25701), .A2(n19663), .B1(n25847), .B2(n25693), .ZN(
        n7061) );
  OAI22_X1 U23206 ( .A1(n25701), .A2(n19662), .B1(n25850), .B2(n25693), .ZN(
        n7062) );
  OAI22_X1 U23207 ( .A1(n25701), .A2(n19661), .B1(n25853), .B2(n25694), .ZN(
        n7063) );
  OAI22_X1 U23208 ( .A1(n25702), .A2(n19660), .B1(n25856), .B2(n25694), .ZN(
        n7064) );
  OAI22_X1 U23209 ( .A1(n25702), .A2(n19659), .B1(n25859), .B2(n25694), .ZN(
        n7065) );
  OAI22_X1 U23210 ( .A1(n25702), .A2(n19658), .B1(n25862), .B2(n25694), .ZN(
        n7066) );
  OAI22_X1 U23211 ( .A1(n25702), .A2(n19657), .B1(n25865), .B2(n25694), .ZN(
        n7067) );
  OAI22_X1 U23212 ( .A1(n25702), .A2(n19656), .B1(n25868), .B2(n25694), .ZN(
        n7068) );
  OAI22_X1 U23213 ( .A1(n25702), .A2(n19655), .B1(n25871), .B2(n25694), .ZN(
        n7069) );
  OAI22_X1 U23214 ( .A1(n25702), .A2(n19654), .B1(n25874), .B2(n25694), .ZN(
        n7070) );
  OAI22_X1 U23215 ( .A1(n25702), .A2(n19653), .B1(n25877), .B2(n25694), .ZN(
        n7071) );
  OAI22_X1 U23216 ( .A1(n25702), .A2(n19652), .B1(n25880), .B2(n25694), .ZN(
        n7072) );
  OAI22_X1 U23217 ( .A1(n25702), .A2(n19651), .B1(n25883), .B2(n25694), .ZN(
        n7073) );
  OAI22_X1 U23218 ( .A1(n25702), .A2(n19650), .B1(n25886), .B2(n25694), .ZN(
        n7074) );
  OAI22_X1 U23219 ( .A1(n25702), .A2(n19649), .B1(n25889), .B2(n25695), .ZN(
        n7075) );
  OAI22_X1 U23220 ( .A1(n25702), .A2(n19648), .B1(n25892), .B2(n25695), .ZN(
        n7076) );
  OAI22_X1 U23221 ( .A1(n25703), .A2(n19647), .B1(n25895), .B2(n25695), .ZN(
        n7077) );
  OAI22_X1 U23222 ( .A1(n25703), .A2(n19646), .B1(n25898), .B2(n25695), .ZN(
        n7078) );
  OAI22_X1 U23223 ( .A1(n25703), .A2(n19645), .B1(n25901), .B2(n25695), .ZN(
        n7079) );
  OAI22_X1 U23224 ( .A1(n25703), .A2(n19644), .B1(n25904), .B2(n25695), .ZN(
        n7080) );
  OAI22_X1 U23225 ( .A1(n25703), .A2(n19643), .B1(n25907), .B2(n25695), .ZN(
        n7081) );
  OAI22_X1 U23226 ( .A1(n25703), .A2(n19642), .B1(n25910), .B2(n25695), .ZN(
        n7082) );
  OAI22_X1 U23227 ( .A1(n25703), .A2(n19641), .B1(n25913), .B2(n25695), .ZN(
        n7083) );
  OAI22_X1 U23228 ( .A1(n25703), .A2(n19640), .B1(n25916), .B2(n25695), .ZN(
        n7084) );
  OAI22_X1 U23229 ( .A1(n25703), .A2(n19639), .B1(n25919), .B2(n25695), .ZN(
        n7085) );
  OAI22_X1 U23230 ( .A1(n25703), .A2(n19638), .B1(n25922), .B2(n25695), .ZN(
        n7086) );
  OAI22_X1 U23231 ( .A1(n25703), .A2(n19637), .B1(n25925), .B2(n25696), .ZN(
        n7087) );
  OAI22_X1 U23232 ( .A1(n25703), .A2(n19636), .B1(n25928), .B2(n25696), .ZN(
        n7088) );
  OAI22_X1 U23233 ( .A1(n25703), .A2(n19635), .B1(n25931), .B2(n25696), .ZN(
        n7089) );
  OAI22_X1 U23234 ( .A1(n25704), .A2(n19634), .B1(n25934), .B2(n25696), .ZN(
        n7090) );
  OAI22_X1 U23235 ( .A1(n25704), .A2(n19633), .B1(n25937), .B2(n25696), .ZN(
        n7091) );
  OAI22_X1 U23236 ( .A1(n25704), .A2(n19632), .B1(n25940), .B2(n25696), .ZN(
        n7092) );
  OAI22_X1 U23237 ( .A1(n25704), .A2(n19631), .B1(n25943), .B2(n25696), .ZN(
        n7093) );
  OAI22_X1 U23238 ( .A1(n25704), .A2(n19630), .B1(n25946), .B2(n25696), .ZN(
        n7094) );
  OAI22_X1 U23239 ( .A1(n25704), .A2(n19629), .B1(n25949), .B2(n25696), .ZN(
        n7095) );
  OAI22_X1 U23240 ( .A1(n25704), .A2(n19628), .B1(n25952), .B2(n25696), .ZN(
        n7096) );
  OAI22_X1 U23241 ( .A1(n25704), .A2(n19627), .B1(n25955), .B2(n25696), .ZN(
        n7097) );
  OAI22_X1 U23242 ( .A1(n25704), .A2(n19626), .B1(n25958), .B2(n25696), .ZN(
        n7098) );
  NAND2_X1 U23243 ( .A1(n22753), .A2(n22754), .ZN(n5374) );
  NOR4_X1 U23244 ( .A1(n22780), .A2(n22781), .A3(n22782), .A4(n22783), .ZN(
        n22753) );
  NOR4_X1 U23245 ( .A1(n22755), .A2(n22756), .A3(n22757), .A4(n22758), .ZN(
        n22754) );
  OAI221_X1 U23246 ( .B1(n20710), .B2(n24997), .C1(n8967), .C2(n24991), .A(
        n22801), .ZN(n22780) );
  NAND2_X1 U23247 ( .A1(n22840), .A2(n22841), .ZN(n5371) );
  NOR4_X1 U23248 ( .A1(n22850), .A2(n22851), .A3(n22852), .A4(n22853), .ZN(
        n22840) );
  NOR4_X1 U23249 ( .A1(n22842), .A2(n22843), .A3(n22844), .A4(n22845), .ZN(
        n22841) );
  OAI221_X1 U23250 ( .B1(n20713), .B2(n24997), .C1(n8970), .C2(n24991), .A(
        n22857), .ZN(n22850) );
  NAND2_X1 U23251 ( .A1(n22822), .A2(n22823), .ZN(n5372) );
  NOR4_X1 U23252 ( .A1(n22832), .A2(n22833), .A3(n22834), .A4(n22835), .ZN(
        n22822) );
  NOR4_X1 U23253 ( .A1(n22824), .A2(n22825), .A3(n22826), .A4(n22827), .ZN(
        n22823) );
  OAI221_X1 U23254 ( .B1(n20712), .B2(n24997), .C1(n8969), .C2(n24991), .A(
        n22839), .ZN(n22832) );
  NAND2_X1 U23255 ( .A1(n22804), .A2(n22805), .ZN(n5373) );
  NOR4_X1 U23256 ( .A1(n22814), .A2(n22815), .A3(n22816), .A4(n22817), .ZN(
        n22804) );
  NOR4_X1 U23257 ( .A1(n22806), .A2(n22807), .A3(n22808), .A4(n22809), .ZN(
        n22805) );
  OAI221_X1 U23258 ( .B1(n20711), .B2(n24997), .C1(n8968), .C2(n24991), .A(
        n22821), .ZN(n22814) );
  NAND2_X1 U23259 ( .A1(n21643), .A2(n21644), .ZN(n5435) );
  NOR4_X1 U23260 ( .A1(n21653), .A2(n21654), .A3(n21655), .A4(n21656), .ZN(
        n21643) );
  NOR4_X1 U23261 ( .A1(n21645), .A2(n21646), .A3(n21647), .A4(n21648), .ZN(
        n21644) );
  OAI221_X1 U23262 ( .B1(n20713), .B2(n25195), .C1(n8970), .C2(n25189), .A(
        n21660), .ZN(n21653) );
  NAND2_X1 U23263 ( .A1(n21625), .A2(n21626), .ZN(n5436) );
  NOR4_X1 U23264 ( .A1(n21635), .A2(n21636), .A3(n21637), .A4(n21638), .ZN(
        n21625) );
  NOR4_X1 U23265 ( .A1(n21627), .A2(n21628), .A3(n21629), .A4(n21630), .ZN(
        n21626) );
  OAI221_X1 U23266 ( .B1(n20712), .B2(n25195), .C1(n8969), .C2(n25189), .A(
        n21642), .ZN(n21635) );
  NAND2_X1 U23267 ( .A1(n21607), .A2(n21608), .ZN(n5437) );
  NOR4_X1 U23268 ( .A1(n21617), .A2(n21618), .A3(n21619), .A4(n21620), .ZN(
        n21607) );
  NOR4_X1 U23269 ( .A1(n21609), .A2(n21610), .A3(n21611), .A4(n21612), .ZN(
        n21608) );
  OAI221_X1 U23270 ( .B1(n20711), .B2(n25195), .C1(n8968), .C2(n25189), .A(
        n21624), .ZN(n21617) );
  NAND2_X1 U23271 ( .A1(n21556), .A2(n21557), .ZN(n5438) );
  NOR4_X1 U23272 ( .A1(n21583), .A2(n21584), .A3(n21585), .A4(n21586), .ZN(
        n21556) );
  NOR4_X1 U23273 ( .A1(n21558), .A2(n21559), .A3(n21560), .A4(n21561), .ZN(
        n21557) );
  OAI221_X1 U23274 ( .B1(n20710), .B2(n25195), .C1(n8967), .C2(n25189), .A(
        n21604), .ZN(n21583) );
  NAND2_X1 U23275 ( .A1(n23920), .A2(n23921), .ZN(n5311) );
  NOR4_X1 U23276 ( .A1(n23941), .A2(n23942), .A3(n23943), .A4(n23944), .ZN(
        n23920) );
  NOR4_X1 U23277 ( .A1(n23922), .A2(n23923), .A3(n23924), .A4(n23925), .ZN(
        n23921) );
  OAI221_X1 U23278 ( .B1(n20773), .B2(n24992), .C1(n9030), .C2(n24986), .A(
        n23949), .ZN(n23941) );
  NAND2_X1 U23279 ( .A1(n23902), .A2(n23903), .ZN(n5312) );
  NOR4_X1 U23280 ( .A1(n23912), .A2(n23913), .A3(n23914), .A4(n23915), .ZN(
        n23902) );
  NOR4_X1 U23281 ( .A1(n23904), .A2(n23905), .A3(n23906), .A4(n23907), .ZN(
        n23903) );
  OAI221_X1 U23282 ( .B1(n20772), .B2(n24992), .C1(n9029), .C2(n24986), .A(
        n23919), .ZN(n23912) );
  NAND2_X1 U23283 ( .A1(n23884), .A2(n23885), .ZN(n5313) );
  NOR4_X1 U23284 ( .A1(n23894), .A2(n23895), .A3(n23896), .A4(n23897), .ZN(
        n23884) );
  NOR4_X1 U23285 ( .A1(n23886), .A2(n23887), .A3(n23888), .A4(n23889), .ZN(
        n23885) );
  OAI221_X1 U23286 ( .B1(n20771), .B2(n24992), .C1(n9028), .C2(n24986), .A(
        n23901), .ZN(n23894) );
  NAND2_X1 U23287 ( .A1(n23866), .A2(n23867), .ZN(n5314) );
  NOR4_X1 U23288 ( .A1(n23876), .A2(n23877), .A3(n23878), .A4(n23879), .ZN(
        n23866) );
  NOR4_X1 U23289 ( .A1(n23868), .A2(n23869), .A3(n23870), .A4(n23871), .ZN(
        n23867) );
  OAI221_X1 U23290 ( .B1(n20770), .B2(n24992), .C1(n9027), .C2(n24986), .A(
        n23883), .ZN(n23876) );
  NAND2_X1 U23291 ( .A1(n23848), .A2(n23849), .ZN(n5315) );
  NOR4_X1 U23292 ( .A1(n23858), .A2(n23859), .A3(n23860), .A4(n23861), .ZN(
        n23848) );
  NOR4_X1 U23293 ( .A1(n23850), .A2(n23851), .A3(n23852), .A4(n23853), .ZN(
        n23849) );
  OAI221_X1 U23294 ( .B1(n20769), .B2(n24992), .C1(n9026), .C2(n24986), .A(
        n23865), .ZN(n23858) );
  NAND2_X1 U23295 ( .A1(n23830), .A2(n23831), .ZN(n5316) );
  NOR4_X1 U23296 ( .A1(n23840), .A2(n23841), .A3(n23842), .A4(n23843), .ZN(
        n23830) );
  NOR4_X1 U23297 ( .A1(n23832), .A2(n23833), .A3(n23834), .A4(n23835), .ZN(
        n23831) );
  OAI221_X1 U23298 ( .B1(n20768), .B2(n24992), .C1(n9025), .C2(n24986), .A(
        n23847), .ZN(n23840) );
  NAND2_X1 U23299 ( .A1(n23812), .A2(n23813), .ZN(n5317) );
  NOR4_X1 U23300 ( .A1(n23822), .A2(n23823), .A3(n23824), .A4(n23825), .ZN(
        n23812) );
  NOR4_X1 U23301 ( .A1(n23814), .A2(n23815), .A3(n23816), .A4(n23817), .ZN(
        n23813) );
  OAI221_X1 U23302 ( .B1(n20767), .B2(n24992), .C1(n9024), .C2(n24986), .A(
        n23829), .ZN(n23822) );
  NAND2_X1 U23303 ( .A1(n23794), .A2(n23795), .ZN(n5318) );
  NOR4_X1 U23304 ( .A1(n23804), .A2(n23805), .A3(n23806), .A4(n23807), .ZN(
        n23794) );
  NOR4_X1 U23305 ( .A1(n23796), .A2(n23797), .A3(n23798), .A4(n23799), .ZN(
        n23795) );
  OAI221_X1 U23306 ( .B1(n20766), .B2(n24992), .C1(n9023), .C2(n24986), .A(
        n23811), .ZN(n23804) );
  NAND2_X1 U23307 ( .A1(n23776), .A2(n23777), .ZN(n5319) );
  NOR4_X1 U23308 ( .A1(n23786), .A2(n23787), .A3(n23788), .A4(n23789), .ZN(
        n23776) );
  NOR4_X1 U23309 ( .A1(n23778), .A2(n23779), .A3(n23780), .A4(n23781), .ZN(
        n23777) );
  OAI221_X1 U23310 ( .B1(n20765), .B2(n24992), .C1(n9022), .C2(n24986), .A(
        n23793), .ZN(n23786) );
  NAND2_X1 U23311 ( .A1(n23758), .A2(n23759), .ZN(n5320) );
  NOR4_X1 U23312 ( .A1(n23768), .A2(n23769), .A3(n23770), .A4(n23771), .ZN(
        n23758) );
  NOR4_X1 U23313 ( .A1(n23760), .A2(n23761), .A3(n23762), .A4(n23763), .ZN(
        n23759) );
  OAI221_X1 U23314 ( .B1(n20764), .B2(n24992), .C1(n9021), .C2(n24986), .A(
        n23775), .ZN(n23768) );
  NAND2_X1 U23315 ( .A1(n23740), .A2(n23741), .ZN(n5321) );
  NOR4_X1 U23316 ( .A1(n23750), .A2(n23751), .A3(n23752), .A4(n23753), .ZN(
        n23740) );
  NOR4_X1 U23317 ( .A1(n23742), .A2(n23743), .A3(n23744), .A4(n23745), .ZN(
        n23741) );
  OAI221_X1 U23318 ( .B1(n20763), .B2(n24992), .C1(n9020), .C2(n24986), .A(
        n23757), .ZN(n23750) );
  NAND2_X1 U23319 ( .A1(n23722), .A2(n23723), .ZN(n5322) );
  NOR4_X1 U23320 ( .A1(n23732), .A2(n23733), .A3(n23734), .A4(n23735), .ZN(
        n23722) );
  NOR4_X1 U23321 ( .A1(n23724), .A2(n23725), .A3(n23726), .A4(n23727), .ZN(
        n23723) );
  OAI221_X1 U23322 ( .B1(n20762), .B2(n24992), .C1(n9019), .C2(n24986), .A(
        n23739), .ZN(n23732) );
  NAND2_X1 U23323 ( .A1(n23704), .A2(n23705), .ZN(n5323) );
  NOR4_X1 U23324 ( .A1(n23714), .A2(n23715), .A3(n23716), .A4(n23717), .ZN(
        n23704) );
  NOR4_X1 U23325 ( .A1(n23706), .A2(n23707), .A3(n23708), .A4(n23709), .ZN(
        n23705) );
  OAI221_X1 U23326 ( .B1(n20761), .B2(n24993), .C1(n9018), .C2(n24987), .A(
        n23721), .ZN(n23714) );
  NAND2_X1 U23327 ( .A1(n23686), .A2(n23687), .ZN(n5324) );
  NOR4_X1 U23328 ( .A1(n23696), .A2(n23697), .A3(n23698), .A4(n23699), .ZN(
        n23686) );
  NOR4_X1 U23329 ( .A1(n23688), .A2(n23689), .A3(n23690), .A4(n23691), .ZN(
        n23687) );
  OAI221_X1 U23330 ( .B1(n20760), .B2(n24993), .C1(n9017), .C2(n24987), .A(
        n23703), .ZN(n23696) );
  NAND2_X1 U23331 ( .A1(n23668), .A2(n23669), .ZN(n5325) );
  NOR4_X1 U23332 ( .A1(n23678), .A2(n23679), .A3(n23680), .A4(n23681), .ZN(
        n23668) );
  NOR4_X1 U23333 ( .A1(n23670), .A2(n23671), .A3(n23672), .A4(n23673), .ZN(
        n23669) );
  OAI221_X1 U23334 ( .B1(n20759), .B2(n24993), .C1(n9016), .C2(n24987), .A(
        n23685), .ZN(n23678) );
  NAND2_X1 U23335 ( .A1(n23650), .A2(n23651), .ZN(n5326) );
  NOR4_X1 U23336 ( .A1(n23660), .A2(n23661), .A3(n23662), .A4(n23663), .ZN(
        n23650) );
  NOR4_X1 U23337 ( .A1(n23652), .A2(n23653), .A3(n23654), .A4(n23655), .ZN(
        n23651) );
  OAI221_X1 U23338 ( .B1(n20758), .B2(n24993), .C1(n9015), .C2(n24987), .A(
        n23667), .ZN(n23660) );
  NAND2_X1 U23339 ( .A1(n23632), .A2(n23633), .ZN(n5327) );
  NOR4_X1 U23340 ( .A1(n23642), .A2(n23643), .A3(n23644), .A4(n23645), .ZN(
        n23632) );
  NOR4_X1 U23341 ( .A1(n23634), .A2(n23635), .A3(n23636), .A4(n23637), .ZN(
        n23633) );
  OAI221_X1 U23342 ( .B1(n20757), .B2(n24993), .C1(n9014), .C2(n24987), .A(
        n23649), .ZN(n23642) );
  NAND2_X1 U23343 ( .A1(n23614), .A2(n23615), .ZN(n5328) );
  NOR4_X1 U23344 ( .A1(n23624), .A2(n23625), .A3(n23626), .A4(n23627), .ZN(
        n23614) );
  NOR4_X1 U23345 ( .A1(n23616), .A2(n23617), .A3(n23618), .A4(n23619), .ZN(
        n23615) );
  OAI221_X1 U23346 ( .B1(n20756), .B2(n24993), .C1(n9013), .C2(n24987), .A(
        n23631), .ZN(n23624) );
  NAND2_X1 U23347 ( .A1(n23596), .A2(n23597), .ZN(n5329) );
  NOR4_X1 U23348 ( .A1(n23606), .A2(n23607), .A3(n23608), .A4(n23609), .ZN(
        n23596) );
  NOR4_X1 U23349 ( .A1(n23598), .A2(n23599), .A3(n23600), .A4(n23601), .ZN(
        n23597) );
  OAI221_X1 U23350 ( .B1(n20755), .B2(n24993), .C1(n9012), .C2(n24987), .A(
        n23613), .ZN(n23606) );
  NAND2_X1 U23351 ( .A1(n23578), .A2(n23579), .ZN(n5330) );
  NOR4_X1 U23352 ( .A1(n23588), .A2(n23589), .A3(n23590), .A4(n23591), .ZN(
        n23578) );
  NOR4_X1 U23353 ( .A1(n23580), .A2(n23581), .A3(n23582), .A4(n23583), .ZN(
        n23579) );
  OAI221_X1 U23354 ( .B1(n20754), .B2(n24993), .C1(n9011), .C2(n24987), .A(
        n23595), .ZN(n23588) );
  NAND2_X1 U23355 ( .A1(n23560), .A2(n23561), .ZN(n5331) );
  NOR4_X1 U23356 ( .A1(n23570), .A2(n23571), .A3(n23572), .A4(n23573), .ZN(
        n23560) );
  NOR4_X1 U23357 ( .A1(n23562), .A2(n23563), .A3(n23564), .A4(n23565), .ZN(
        n23561) );
  OAI221_X1 U23358 ( .B1(n20753), .B2(n24993), .C1(n9010), .C2(n24987), .A(
        n23577), .ZN(n23570) );
  NAND2_X1 U23359 ( .A1(n23542), .A2(n23543), .ZN(n5332) );
  NOR4_X1 U23360 ( .A1(n23552), .A2(n23553), .A3(n23554), .A4(n23555), .ZN(
        n23542) );
  NOR4_X1 U23361 ( .A1(n23544), .A2(n23545), .A3(n23546), .A4(n23547), .ZN(
        n23543) );
  OAI221_X1 U23362 ( .B1(n20752), .B2(n24993), .C1(n9009), .C2(n24987), .A(
        n23559), .ZN(n23552) );
  NAND2_X1 U23363 ( .A1(n23524), .A2(n23525), .ZN(n5333) );
  NOR4_X1 U23364 ( .A1(n23534), .A2(n23535), .A3(n23536), .A4(n23537), .ZN(
        n23524) );
  NOR4_X1 U23365 ( .A1(n23526), .A2(n23527), .A3(n23528), .A4(n23529), .ZN(
        n23525) );
  OAI221_X1 U23366 ( .B1(n20751), .B2(n24993), .C1(n9008), .C2(n24987), .A(
        n23541), .ZN(n23534) );
  NAND2_X1 U23367 ( .A1(n23506), .A2(n23507), .ZN(n5334) );
  NOR4_X1 U23368 ( .A1(n23516), .A2(n23517), .A3(n23518), .A4(n23519), .ZN(
        n23506) );
  NOR4_X1 U23369 ( .A1(n23508), .A2(n23509), .A3(n23510), .A4(n23511), .ZN(
        n23507) );
  OAI221_X1 U23370 ( .B1(n20750), .B2(n24993), .C1(n9007), .C2(n24987), .A(
        n23523), .ZN(n23516) );
  NAND2_X1 U23371 ( .A1(n23488), .A2(n23489), .ZN(n5335) );
  NOR4_X1 U23372 ( .A1(n23498), .A2(n23499), .A3(n23500), .A4(n23501), .ZN(
        n23488) );
  NOR4_X1 U23373 ( .A1(n23490), .A2(n23491), .A3(n23492), .A4(n23493), .ZN(
        n23489) );
  OAI221_X1 U23374 ( .B1(n20749), .B2(n24994), .C1(n9006), .C2(n24988), .A(
        n23505), .ZN(n23498) );
  NAND2_X1 U23375 ( .A1(n23470), .A2(n23471), .ZN(n5336) );
  NOR4_X1 U23376 ( .A1(n23480), .A2(n23481), .A3(n23482), .A4(n23483), .ZN(
        n23470) );
  NOR4_X1 U23377 ( .A1(n23472), .A2(n23473), .A3(n23474), .A4(n23475), .ZN(
        n23471) );
  OAI221_X1 U23378 ( .B1(n20748), .B2(n24994), .C1(n9005), .C2(n24988), .A(
        n23487), .ZN(n23480) );
  NAND2_X1 U23379 ( .A1(n23452), .A2(n23453), .ZN(n5337) );
  NOR4_X1 U23380 ( .A1(n23462), .A2(n23463), .A3(n23464), .A4(n23465), .ZN(
        n23452) );
  NOR4_X1 U23381 ( .A1(n23454), .A2(n23455), .A3(n23456), .A4(n23457), .ZN(
        n23453) );
  OAI221_X1 U23382 ( .B1(n20747), .B2(n24994), .C1(n9004), .C2(n24988), .A(
        n23469), .ZN(n23462) );
  NAND2_X1 U23383 ( .A1(n23434), .A2(n23435), .ZN(n5338) );
  NOR4_X1 U23384 ( .A1(n23444), .A2(n23445), .A3(n23446), .A4(n23447), .ZN(
        n23434) );
  NOR4_X1 U23385 ( .A1(n23436), .A2(n23437), .A3(n23438), .A4(n23439), .ZN(
        n23435) );
  OAI221_X1 U23386 ( .B1(n20746), .B2(n24994), .C1(n9003), .C2(n24988), .A(
        n23451), .ZN(n23444) );
  NAND2_X1 U23387 ( .A1(n23416), .A2(n23417), .ZN(n5339) );
  NOR4_X1 U23388 ( .A1(n23426), .A2(n23427), .A3(n23428), .A4(n23429), .ZN(
        n23416) );
  NOR4_X1 U23389 ( .A1(n23418), .A2(n23419), .A3(n23420), .A4(n23421), .ZN(
        n23417) );
  OAI221_X1 U23390 ( .B1(n20745), .B2(n24994), .C1(n9002), .C2(n24988), .A(
        n23433), .ZN(n23426) );
  NAND2_X1 U23391 ( .A1(n23398), .A2(n23399), .ZN(n5340) );
  NOR4_X1 U23392 ( .A1(n23408), .A2(n23409), .A3(n23410), .A4(n23411), .ZN(
        n23398) );
  NOR4_X1 U23393 ( .A1(n23400), .A2(n23401), .A3(n23402), .A4(n23403), .ZN(
        n23399) );
  OAI221_X1 U23394 ( .B1(n20744), .B2(n24994), .C1(n9001), .C2(n24988), .A(
        n23415), .ZN(n23408) );
  NAND2_X1 U23395 ( .A1(n23380), .A2(n23381), .ZN(n5341) );
  NOR4_X1 U23396 ( .A1(n23390), .A2(n23391), .A3(n23392), .A4(n23393), .ZN(
        n23380) );
  NOR4_X1 U23397 ( .A1(n23382), .A2(n23383), .A3(n23384), .A4(n23385), .ZN(
        n23381) );
  OAI221_X1 U23398 ( .B1(n20743), .B2(n24994), .C1(n9000), .C2(n24988), .A(
        n23397), .ZN(n23390) );
  NAND2_X1 U23399 ( .A1(n23362), .A2(n23363), .ZN(n5342) );
  NOR4_X1 U23400 ( .A1(n23372), .A2(n23373), .A3(n23374), .A4(n23375), .ZN(
        n23362) );
  NOR4_X1 U23401 ( .A1(n23364), .A2(n23365), .A3(n23366), .A4(n23367), .ZN(
        n23363) );
  OAI221_X1 U23402 ( .B1(n20742), .B2(n24994), .C1(n8999), .C2(n24988), .A(
        n23379), .ZN(n23372) );
  NAND2_X1 U23403 ( .A1(n23344), .A2(n23345), .ZN(n5343) );
  NOR4_X1 U23404 ( .A1(n23354), .A2(n23355), .A3(n23356), .A4(n23357), .ZN(
        n23344) );
  NOR4_X1 U23405 ( .A1(n23346), .A2(n23347), .A3(n23348), .A4(n23349), .ZN(
        n23345) );
  OAI221_X1 U23406 ( .B1(n20741), .B2(n24994), .C1(n8998), .C2(n24988), .A(
        n23361), .ZN(n23354) );
  NAND2_X1 U23407 ( .A1(n23326), .A2(n23327), .ZN(n5344) );
  NOR4_X1 U23408 ( .A1(n23336), .A2(n23337), .A3(n23338), .A4(n23339), .ZN(
        n23326) );
  NOR4_X1 U23409 ( .A1(n23328), .A2(n23329), .A3(n23330), .A4(n23331), .ZN(
        n23327) );
  OAI221_X1 U23410 ( .B1(n20740), .B2(n24994), .C1(n8997), .C2(n24988), .A(
        n23343), .ZN(n23336) );
  NAND2_X1 U23411 ( .A1(n23308), .A2(n23309), .ZN(n5345) );
  NOR4_X1 U23412 ( .A1(n23318), .A2(n23319), .A3(n23320), .A4(n23321), .ZN(
        n23308) );
  NOR4_X1 U23413 ( .A1(n23310), .A2(n23311), .A3(n23312), .A4(n23313), .ZN(
        n23309) );
  OAI221_X1 U23414 ( .B1(n20739), .B2(n24994), .C1(n8996), .C2(n24988), .A(
        n23325), .ZN(n23318) );
  NAND2_X1 U23415 ( .A1(n23290), .A2(n23291), .ZN(n5346) );
  NOR4_X1 U23416 ( .A1(n23300), .A2(n23301), .A3(n23302), .A4(n23303), .ZN(
        n23290) );
  NOR4_X1 U23417 ( .A1(n23292), .A2(n23293), .A3(n23294), .A4(n23295), .ZN(
        n23291) );
  OAI221_X1 U23418 ( .B1(n20738), .B2(n24994), .C1(n8995), .C2(n24988), .A(
        n23307), .ZN(n23300) );
  NAND2_X1 U23419 ( .A1(n23272), .A2(n23273), .ZN(n5347) );
  NOR4_X1 U23420 ( .A1(n23282), .A2(n23283), .A3(n23284), .A4(n23285), .ZN(
        n23272) );
  NOR4_X1 U23421 ( .A1(n23274), .A2(n23275), .A3(n23276), .A4(n23277), .ZN(
        n23273) );
  OAI221_X1 U23422 ( .B1(n20737), .B2(n24995), .C1(n8994), .C2(n24989), .A(
        n23289), .ZN(n23282) );
  NAND2_X1 U23423 ( .A1(n23254), .A2(n23255), .ZN(n5348) );
  NOR4_X1 U23424 ( .A1(n23264), .A2(n23265), .A3(n23266), .A4(n23267), .ZN(
        n23254) );
  NOR4_X1 U23425 ( .A1(n23256), .A2(n23257), .A3(n23258), .A4(n23259), .ZN(
        n23255) );
  OAI221_X1 U23426 ( .B1(n20736), .B2(n24995), .C1(n8993), .C2(n24989), .A(
        n23271), .ZN(n23264) );
  NAND2_X1 U23427 ( .A1(n23236), .A2(n23237), .ZN(n5349) );
  NOR4_X1 U23428 ( .A1(n23246), .A2(n23247), .A3(n23248), .A4(n23249), .ZN(
        n23236) );
  NOR4_X1 U23429 ( .A1(n23238), .A2(n23239), .A3(n23240), .A4(n23241), .ZN(
        n23237) );
  OAI221_X1 U23430 ( .B1(n20735), .B2(n24995), .C1(n8992), .C2(n24989), .A(
        n23253), .ZN(n23246) );
  NAND2_X1 U23431 ( .A1(n23218), .A2(n23219), .ZN(n5350) );
  NOR4_X1 U23432 ( .A1(n23228), .A2(n23229), .A3(n23230), .A4(n23231), .ZN(
        n23218) );
  NOR4_X1 U23433 ( .A1(n23220), .A2(n23221), .A3(n23222), .A4(n23223), .ZN(
        n23219) );
  OAI221_X1 U23434 ( .B1(n20734), .B2(n24995), .C1(n8991), .C2(n24989), .A(
        n23235), .ZN(n23228) );
  NAND2_X1 U23435 ( .A1(n23200), .A2(n23201), .ZN(n5351) );
  NOR4_X1 U23436 ( .A1(n23210), .A2(n23211), .A3(n23212), .A4(n23213), .ZN(
        n23200) );
  NOR4_X1 U23437 ( .A1(n23202), .A2(n23203), .A3(n23204), .A4(n23205), .ZN(
        n23201) );
  OAI221_X1 U23438 ( .B1(n20733), .B2(n24995), .C1(n8990), .C2(n24989), .A(
        n23217), .ZN(n23210) );
  NAND2_X1 U23439 ( .A1(n23182), .A2(n23183), .ZN(n5352) );
  NOR4_X1 U23440 ( .A1(n23192), .A2(n23193), .A3(n23194), .A4(n23195), .ZN(
        n23182) );
  NOR4_X1 U23441 ( .A1(n23184), .A2(n23185), .A3(n23186), .A4(n23187), .ZN(
        n23183) );
  OAI221_X1 U23442 ( .B1(n20732), .B2(n24995), .C1(n8989), .C2(n24989), .A(
        n23199), .ZN(n23192) );
  NAND2_X1 U23443 ( .A1(n23164), .A2(n23165), .ZN(n5353) );
  NOR4_X1 U23444 ( .A1(n23174), .A2(n23175), .A3(n23176), .A4(n23177), .ZN(
        n23164) );
  NOR4_X1 U23445 ( .A1(n23166), .A2(n23167), .A3(n23168), .A4(n23169), .ZN(
        n23165) );
  OAI221_X1 U23446 ( .B1(n20731), .B2(n24995), .C1(n8988), .C2(n24989), .A(
        n23181), .ZN(n23174) );
  NAND2_X1 U23447 ( .A1(n23146), .A2(n23147), .ZN(n5354) );
  NOR4_X1 U23448 ( .A1(n23156), .A2(n23157), .A3(n23158), .A4(n23159), .ZN(
        n23146) );
  NOR4_X1 U23449 ( .A1(n23148), .A2(n23149), .A3(n23150), .A4(n23151), .ZN(
        n23147) );
  OAI221_X1 U23450 ( .B1(n20730), .B2(n24995), .C1(n8987), .C2(n24989), .A(
        n23163), .ZN(n23156) );
  NAND2_X1 U23451 ( .A1(n23128), .A2(n23129), .ZN(n5355) );
  NOR4_X1 U23452 ( .A1(n23138), .A2(n23139), .A3(n23140), .A4(n23141), .ZN(
        n23128) );
  NOR4_X1 U23453 ( .A1(n23130), .A2(n23131), .A3(n23132), .A4(n23133), .ZN(
        n23129) );
  OAI221_X1 U23454 ( .B1(n20729), .B2(n24995), .C1(n8986), .C2(n24989), .A(
        n23145), .ZN(n23138) );
  NAND2_X1 U23455 ( .A1(n23110), .A2(n23111), .ZN(n5356) );
  NOR4_X1 U23456 ( .A1(n23120), .A2(n23121), .A3(n23122), .A4(n23123), .ZN(
        n23110) );
  NOR4_X1 U23457 ( .A1(n23112), .A2(n23113), .A3(n23114), .A4(n23115), .ZN(
        n23111) );
  OAI221_X1 U23458 ( .B1(n20728), .B2(n24995), .C1(n8985), .C2(n24989), .A(
        n23127), .ZN(n23120) );
  NAND2_X1 U23459 ( .A1(n23092), .A2(n23093), .ZN(n5357) );
  NOR4_X1 U23460 ( .A1(n23102), .A2(n23103), .A3(n23104), .A4(n23105), .ZN(
        n23092) );
  NOR4_X1 U23461 ( .A1(n23094), .A2(n23095), .A3(n23096), .A4(n23097), .ZN(
        n23093) );
  OAI221_X1 U23462 ( .B1(n20727), .B2(n24995), .C1(n8984), .C2(n24989), .A(
        n23109), .ZN(n23102) );
  NAND2_X1 U23463 ( .A1(n23074), .A2(n23075), .ZN(n5358) );
  NOR4_X1 U23464 ( .A1(n23084), .A2(n23085), .A3(n23086), .A4(n23087), .ZN(
        n23074) );
  NOR4_X1 U23465 ( .A1(n23076), .A2(n23077), .A3(n23078), .A4(n23079), .ZN(
        n23075) );
  OAI221_X1 U23466 ( .B1(n20726), .B2(n24995), .C1(n8983), .C2(n24989), .A(
        n23091), .ZN(n23084) );
  NAND2_X1 U23467 ( .A1(n23056), .A2(n23057), .ZN(n5359) );
  NOR4_X1 U23468 ( .A1(n23066), .A2(n23067), .A3(n23068), .A4(n23069), .ZN(
        n23056) );
  NOR4_X1 U23469 ( .A1(n23058), .A2(n23059), .A3(n23060), .A4(n23061), .ZN(
        n23057) );
  OAI221_X1 U23470 ( .B1(n20725), .B2(n24996), .C1(n8982), .C2(n24990), .A(
        n23073), .ZN(n23066) );
  NAND2_X1 U23471 ( .A1(n23038), .A2(n23039), .ZN(n5360) );
  NOR4_X1 U23472 ( .A1(n23048), .A2(n23049), .A3(n23050), .A4(n23051), .ZN(
        n23038) );
  NOR4_X1 U23473 ( .A1(n23040), .A2(n23041), .A3(n23042), .A4(n23043), .ZN(
        n23039) );
  OAI221_X1 U23474 ( .B1(n20724), .B2(n24996), .C1(n8981), .C2(n24990), .A(
        n23055), .ZN(n23048) );
  NAND2_X1 U23475 ( .A1(n23020), .A2(n23021), .ZN(n5361) );
  NOR4_X1 U23476 ( .A1(n23030), .A2(n23031), .A3(n23032), .A4(n23033), .ZN(
        n23020) );
  NOR4_X1 U23477 ( .A1(n23022), .A2(n23023), .A3(n23024), .A4(n23025), .ZN(
        n23021) );
  OAI221_X1 U23478 ( .B1(n20723), .B2(n24996), .C1(n8980), .C2(n24990), .A(
        n23037), .ZN(n23030) );
  NAND2_X1 U23479 ( .A1(n23002), .A2(n23003), .ZN(n5362) );
  NOR4_X1 U23480 ( .A1(n23012), .A2(n23013), .A3(n23014), .A4(n23015), .ZN(
        n23002) );
  NOR4_X1 U23481 ( .A1(n23004), .A2(n23005), .A3(n23006), .A4(n23007), .ZN(
        n23003) );
  OAI221_X1 U23482 ( .B1(n20722), .B2(n24996), .C1(n8979), .C2(n24990), .A(
        n23019), .ZN(n23012) );
  NAND2_X1 U23483 ( .A1(n22984), .A2(n22985), .ZN(n5363) );
  NOR4_X1 U23484 ( .A1(n22994), .A2(n22995), .A3(n22996), .A4(n22997), .ZN(
        n22984) );
  NOR4_X1 U23485 ( .A1(n22986), .A2(n22987), .A3(n22988), .A4(n22989), .ZN(
        n22985) );
  OAI221_X1 U23486 ( .B1(n20721), .B2(n24996), .C1(n8978), .C2(n24990), .A(
        n23001), .ZN(n22994) );
  NAND2_X1 U23487 ( .A1(n22966), .A2(n22967), .ZN(n5364) );
  NOR4_X1 U23488 ( .A1(n22976), .A2(n22977), .A3(n22978), .A4(n22979), .ZN(
        n22966) );
  NOR4_X1 U23489 ( .A1(n22968), .A2(n22969), .A3(n22970), .A4(n22971), .ZN(
        n22967) );
  OAI221_X1 U23490 ( .B1(n20720), .B2(n24996), .C1(n8977), .C2(n24990), .A(
        n22983), .ZN(n22976) );
  NAND2_X1 U23491 ( .A1(n22948), .A2(n22949), .ZN(n5365) );
  NOR4_X1 U23492 ( .A1(n22958), .A2(n22959), .A3(n22960), .A4(n22961), .ZN(
        n22948) );
  NOR4_X1 U23493 ( .A1(n22950), .A2(n22951), .A3(n22952), .A4(n22953), .ZN(
        n22949) );
  OAI221_X1 U23494 ( .B1(n20719), .B2(n24996), .C1(n8976), .C2(n24990), .A(
        n22965), .ZN(n22958) );
  NAND2_X1 U23495 ( .A1(n22930), .A2(n22931), .ZN(n5366) );
  NOR4_X1 U23496 ( .A1(n22940), .A2(n22941), .A3(n22942), .A4(n22943), .ZN(
        n22930) );
  NOR4_X1 U23497 ( .A1(n22932), .A2(n22933), .A3(n22934), .A4(n22935), .ZN(
        n22931) );
  OAI221_X1 U23498 ( .B1(n20718), .B2(n24996), .C1(n8975), .C2(n24990), .A(
        n22947), .ZN(n22940) );
  NAND2_X1 U23499 ( .A1(n22912), .A2(n22913), .ZN(n5367) );
  NOR4_X1 U23500 ( .A1(n22922), .A2(n22923), .A3(n22924), .A4(n22925), .ZN(
        n22912) );
  NOR4_X1 U23501 ( .A1(n22914), .A2(n22915), .A3(n22916), .A4(n22917), .ZN(
        n22913) );
  OAI221_X1 U23502 ( .B1(n20717), .B2(n24996), .C1(n8974), .C2(n24990), .A(
        n22929), .ZN(n22922) );
  NAND2_X1 U23503 ( .A1(n22894), .A2(n22895), .ZN(n5368) );
  NOR4_X1 U23504 ( .A1(n22904), .A2(n22905), .A3(n22906), .A4(n22907), .ZN(
        n22894) );
  NOR4_X1 U23505 ( .A1(n22896), .A2(n22897), .A3(n22898), .A4(n22899), .ZN(
        n22895) );
  OAI221_X1 U23506 ( .B1(n20716), .B2(n24996), .C1(n8973), .C2(n24990), .A(
        n22911), .ZN(n22904) );
  NAND2_X1 U23507 ( .A1(n22876), .A2(n22877), .ZN(n5369) );
  NOR4_X1 U23508 ( .A1(n22886), .A2(n22887), .A3(n22888), .A4(n22889), .ZN(
        n22876) );
  NOR4_X1 U23509 ( .A1(n22878), .A2(n22879), .A3(n22880), .A4(n22881), .ZN(
        n22877) );
  OAI221_X1 U23510 ( .B1(n20715), .B2(n24996), .C1(n8972), .C2(n24990), .A(
        n22893), .ZN(n22886) );
  NAND2_X1 U23511 ( .A1(n22858), .A2(n22859), .ZN(n5370) );
  NOR4_X1 U23512 ( .A1(n22868), .A2(n22869), .A3(n22870), .A4(n22871), .ZN(
        n22858) );
  NOR4_X1 U23513 ( .A1(n22860), .A2(n22861), .A3(n22862), .A4(n22863), .ZN(
        n22859) );
  OAI221_X1 U23514 ( .B1(n20714), .B2(n24996), .C1(n8971), .C2(n24990), .A(
        n22875), .ZN(n22868) );
  NAND2_X1 U23515 ( .A1(n22723), .A2(n22724), .ZN(n5375) );
  NOR4_X1 U23516 ( .A1(n22744), .A2(n22745), .A3(n22746), .A4(n22747), .ZN(
        n22723) );
  NOR4_X1 U23517 ( .A1(n22725), .A2(n22726), .A3(n22727), .A4(n22728), .ZN(
        n22724) );
  OAI221_X1 U23518 ( .B1(n20773), .B2(n25190), .C1(n9030), .C2(n25184), .A(
        n22752), .ZN(n22744) );
  NAND2_X1 U23519 ( .A1(n22705), .A2(n22706), .ZN(n5376) );
  NOR4_X1 U23520 ( .A1(n22715), .A2(n22716), .A3(n22717), .A4(n22718), .ZN(
        n22705) );
  NOR4_X1 U23521 ( .A1(n22707), .A2(n22708), .A3(n22709), .A4(n22710), .ZN(
        n22706) );
  OAI221_X1 U23522 ( .B1(n20772), .B2(n25190), .C1(n9029), .C2(n25184), .A(
        n22722), .ZN(n22715) );
  NAND2_X1 U23523 ( .A1(n22687), .A2(n22688), .ZN(n5377) );
  NOR4_X1 U23524 ( .A1(n22697), .A2(n22698), .A3(n22699), .A4(n22700), .ZN(
        n22687) );
  NOR4_X1 U23525 ( .A1(n22689), .A2(n22690), .A3(n22691), .A4(n22692), .ZN(
        n22688) );
  OAI221_X1 U23526 ( .B1(n20771), .B2(n25190), .C1(n9028), .C2(n25184), .A(
        n22704), .ZN(n22697) );
  NAND2_X1 U23527 ( .A1(n22669), .A2(n22670), .ZN(n5378) );
  NOR4_X1 U23528 ( .A1(n22679), .A2(n22680), .A3(n22681), .A4(n22682), .ZN(
        n22669) );
  NOR4_X1 U23529 ( .A1(n22671), .A2(n22672), .A3(n22673), .A4(n22674), .ZN(
        n22670) );
  OAI221_X1 U23530 ( .B1(n20770), .B2(n25190), .C1(n9027), .C2(n25184), .A(
        n22686), .ZN(n22679) );
  NAND2_X1 U23531 ( .A1(n22651), .A2(n22652), .ZN(n5379) );
  NOR4_X1 U23532 ( .A1(n22661), .A2(n22662), .A3(n22663), .A4(n22664), .ZN(
        n22651) );
  NOR4_X1 U23533 ( .A1(n22653), .A2(n22654), .A3(n22655), .A4(n22656), .ZN(
        n22652) );
  OAI221_X1 U23534 ( .B1(n20769), .B2(n25190), .C1(n9026), .C2(n25184), .A(
        n22668), .ZN(n22661) );
  NAND2_X1 U23535 ( .A1(n22633), .A2(n22634), .ZN(n5380) );
  NOR4_X1 U23536 ( .A1(n22643), .A2(n22644), .A3(n22645), .A4(n22646), .ZN(
        n22633) );
  NOR4_X1 U23537 ( .A1(n22635), .A2(n22636), .A3(n22637), .A4(n22638), .ZN(
        n22634) );
  OAI221_X1 U23538 ( .B1(n20768), .B2(n25190), .C1(n9025), .C2(n25184), .A(
        n22650), .ZN(n22643) );
  NAND2_X1 U23539 ( .A1(n22615), .A2(n22616), .ZN(n5381) );
  NOR4_X1 U23540 ( .A1(n22625), .A2(n22626), .A3(n22627), .A4(n22628), .ZN(
        n22615) );
  NOR4_X1 U23541 ( .A1(n22617), .A2(n22618), .A3(n22619), .A4(n22620), .ZN(
        n22616) );
  OAI221_X1 U23542 ( .B1(n20767), .B2(n25190), .C1(n9024), .C2(n25184), .A(
        n22632), .ZN(n22625) );
  NAND2_X1 U23543 ( .A1(n22597), .A2(n22598), .ZN(n5382) );
  NOR4_X1 U23544 ( .A1(n22607), .A2(n22608), .A3(n22609), .A4(n22610), .ZN(
        n22597) );
  NOR4_X1 U23545 ( .A1(n22599), .A2(n22600), .A3(n22601), .A4(n22602), .ZN(
        n22598) );
  OAI221_X1 U23546 ( .B1(n20766), .B2(n25190), .C1(n9023), .C2(n25184), .A(
        n22614), .ZN(n22607) );
  NAND2_X1 U23547 ( .A1(n22579), .A2(n22580), .ZN(n5383) );
  NOR4_X1 U23548 ( .A1(n22589), .A2(n22590), .A3(n22591), .A4(n22592), .ZN(
        n22579) );
  NOR4_X1 U23549 ( .A1(n22581), .A2(n22582), .A3(n22583), .A4(n22584), .ZN(
        n22580) );
  OAI221_X1 U23550 ( .B1(n20765), .B2(n25190), .C1(n9022), .C2(n25184), .A(
        n22596), .ZN(n22589) );
  NAND2_X1 U23551 ( .A1(n22561), .A2(n22562), .ZN(n5384) );
  NOR4_X1 U23552 ( .A1(n22571), .A2(n22572), .A3(n22573), .A4(n22574), .ZN(
        n22561) );
  NOR4_X1 U23553 ( .A1(n22563), .A2(n22564), .A3(n22565), .A4(n22566), .ZN(
        n22562) );
  OAI221_X1 U23554 ( .B1(n20764), .B2(n25190), .C1(n9021), .C2(n25184), .A(
        n22578), .ZN(n22571) );
  NAND2_X1 U23555 ( .A1(n22543), .A2(n22544), .ZN(n5385) );
  NOR4_X1 U23556 ( .A1(n22553), .A2(n22554), .A3(n22555), .A4(n22556), .ZN(
        n22543) );
  NOR4_X1 U23557 ( .A1(n22545), .A2(n22546), .A3(n22547), .A4(n22548), .ZN(
        n22544) );
  OAI221_X1 U23558 ( .B1(n20763), .B2(n25190), .C1(n9020), .C2(n25184), .A(
        n22560), .ZN(n22553) );
  NAND2_X1 U23559 ( .A1(n22525), .A2(n22526), .ZN(n5386) );
  NOR4_X1 U23560 ( .A1(n22535), .A2(n22536), .A3(n22537), .A4(n22538), .ZN(
        n22525) );
  NOR4_X1 U23561 ( .A1(n22527), .A2(n22528), .A3(n22529), .A4(n22530), .ZN(
        n22526) );
  OAI221_X1 U23562 ( .B1(n20762), .B2(n25190), .C1(n9019), .C2(n25184), .A(
        n22542), .ZN(n22535) );
  NAND2_X1 U23563 ( .A1(n22507), .A2(n22508), .ZN(n5387) );
  NOR4_X1 U23564 ( .A1(n22517), .A2(n22518), .A3(n22519), .A4(n22520), .ZN(
        n22507) );
  NOR4_X1 U23565 ( .A1(n22509), .A2(n22510), .A3(n22511), .A4(n22512), .ZN(
        n22508) );
  OAI221_X1 U23566 ( .B1(n20761), .B2(n25191), .C1(n9018), .C2(n25185), .A(
        n22524), .ZN(n22517) );
  NAND2_X1 U23567 ( .A1(n22489), .A2(n22490), .ZN(n5388) );
  NOR4_X1 U23568 ( .A1(n22499), .A2(n22500), .A3(n22501), .A4(n22502), .ZN(
        n22489) );
  NOR4_X1 U23569 ( .A1(n22491), .A2(n22492), .A3(n22493), .A4(n22494), .ZN(
        n22490) );
  OAI221_X1 U23570 ( .B1(n20760), .B2(n25191), .C1(n9017), .C2(n25185), .A(
        n22506), .ZN(n22499) );
  NAND2_X1 U23571 ( .A1(n22471), .A2(n22472), .ZN(n5389) );
  NOR4_X1 U23572 ( .A1(n22481), .A2(n22482), .A3(n22483), .A4(n22484), .ZN(
        n22471) );
  NOR4_X1 U23573 ( .A1(n22473), .A2(n22474), .A3(n22475), .A4(n22476), .ZN(
        n22472) );
  OAI221_X1 U23574 ( .B1(n20759), .B2(n25191), .C1(n9016), .C2(n25185), .A(
        n22488), .ZN(n22481) );
  NAND2_X1 U23575 ( .A1(n22453), .A2(n22454), .ZN(n5390) );
  NOR4_X1 U23576 ( .A1(n22463), .A2(n22464), .A3(n22465), .A4(n22466), .ZN(
        n22453) );
  NOR4_X1 U23577 ( .A1(n22455), .A2(n22456), .A3(n22457), .A4(n22458), .ZN(
        n22454) );
  OAI221_X1 U23578 ( .B1(n20758), .B2(n25191), .C1(n9015), .C2(n25185), .A(
        n22470), .ZN(n22463) );
  NAND2_X1 U23579 ( .A1(n22435), .A2(n22436), .ZN(n5391) );
  NOR4_X1 U23580 ( .A1(n22445), .A2(n22446), .A3(n22447), .A4(n22448), .ZN(
        n22435) );
  NOR4_X1 U23581 ( .A1(n22437), .A2(n22438), .A3(n22439), .A4(n22440), .ZN(
        n22436) );
  OAI221_X1 U23582 ( .B1(n20757), .B2(n25191), .C1(n9014), .C2(n25185), .A(
        n22452), .ZN(n22445) );
  NAND2_X1 U23583 ( .A1(n22417), .A2(n22418), .ZN(n5392) );
  NOR4_X1 U23584 ( .A1(n22427), .A2(n22428), .A3(n22429), .A4(n22430), .ZN(
        n22417) );
  NOR4_X1 U23585 ( .A1(n22419), .A2(n22420), .A3(n22421), .A4(n22422), .ZN(
        n22418) );
  OAI221_X1 U23586 ( .B1(n20756), .B2(n25191), .C1(n9013), .C2(n25185), .A(
        n22434), .ZN(n22427) );
  NAND2_X1 U23587 ( .A1(n22399), .A2(n22400), .ZN(n5393) );
  NOR4_X1 U23588 ( .A1(n22409), .A2(n22410), .A3(n22411), .A4(n22412), .ZN(
        n22399) );
  NOR4_X1 U23589 ( .A1(n22401), .A2(n22402), .A3(n22403), .A4(n22404), .ZN(
        n22400) );
  OAI221_X1 U23590 ( .B1(n20755), .B2(n25191), .C1(n9012), .C2(n25185), .A(
        n22416), .ZN(n22409) );
  NAND2_X1 U23591 ( .A1(n22381), .A2(n22382), .ZN(n5394) );
  NOR4_X1 U23592 ( .A1(n22391), .A2(n22392), .A3(n22393), .A4(n22394), .ZN(
        n22381) );
  NOR4_X1 U23593 ( .A1(n22383), .A2(n22384), .A3(n22385), .A4(n22386), .ZN(
        n22382) );
  OAI221_X1 U23594 ( .B1(n20754), .B2(n25191), .C1(n9011), .C2(n25185), .A(
        n22398), .ZN(n22391) );
  NAND2_X1 U23595 ( .A1(n22363), .A2(n22364), .ZN(n5395) );
  NOR4_X1 U23596 ( .A1(n22373), .A2(n22374), .A3(n22375), .A4(n22376), .ZN(
        n22363) );
  NOR4_X1 U23597 ( .A1(n22365), .A2(n22366), .A3(n22367), .A4(n22368), .ZN(
        n22364) );
  OAI221_X1 U23598 ( .B1(n20753), .B2(n25191), .C1(n9010), .C2(n25185), .A(
        n22380), .ZN(n22373) );
  NAND2_X1 U23599 ( .A1(n22345), .A2(n22346), .ZN(n5396) );
  NOR4_X1 U23600 ( .A1(n22355), .A2(n22356), .A3(n22357), .A4(n22358), .ZN(
        n22345) );
  NOR4_X1 U23601 ( .A1(n22347), .A2(n22348), .A3(n22349), .A4(n22350), .ZN(
        n22346) );
  OAI221_X1 U23602 ( .B1(n20752), .B2(n25191), .C1(n9009), .C2(n25185), .A(
        n22362), .ZN(n22355) );
  NAND2_X1 U23603 ( .A1(n22327), .A2(n22328), .ZN(n5397) );
  NOR4_X1 U23604 ( .A1(n22337), .A2(n22338), .A3(n22339), .A4(n22340), .ZN(
        n22327) );
  NOR4_X1 U23605 ( .A1(n22329), .A2(n22330), .A3(n22331), .A4(n22332), .ZN(
        n22328) );
  OAI221_X1 U23606 ( .B1(n20751), .B2(n25191), .C1(n9008), .C2(n25185), .A(
        n22344), .ZN(n22337) );
  NAND2_X1 U23607 ( .A1(n22309), .A2(n22310), .ZN(n5398) );
  NOR4_X1 U23608 ( .A1(n22319), .A2(n22320), .A3(n22321), .A4(n22322), .ZN(
        n22309) );
  NOR4_X1 U23609 ( .A1(n22311), .A2(n22312), .A3(n22313), .A4(n22314), .ZN(
        n22310) );
  OAI221_X1 U23610 ( .B1(n20750), .B2(n25191), .C1(n9007), .C2(n25185), .A(
        n22326), .ZN(n22319) );
  NAND2_X1 U23611 ( .A1(n22291), .A2(n22292), .ZN(n5399) );
  NOR4_X1 U23612 ( .A1(n22301), .A2(n22302), .A3(n22303), .A4(n22304), .ZN(
        n22291) );
  NOR4_X1 U23613 ( .A1(n22293), .A2(n22294), .A3(n22295), .A4(n22296), .ZN(
        n22292) );
  OAI221_X1 U23614 ( .B1(n20749), .B2(n25192), .C1(n9006), .C2(n25186), .A(
        n22308), .ZN(n22301) );
  NAND2_X1 U23615 ( .A1(n22273), .A2(n22274), .ZN(n5400) );
  NOR4_X1 U23616 ( .A1(n22283), .A2(n22284), .A3(n22285), .A4(n22286), .ZN(
        n22273) );
  NOR4_X1 U23617 ( .A1(n22275), .A2(n22276), .A3(n22277), .A4(n22278), .ZN(
        n22274) );
  OAI221_X1 U23618 ( .B1(n20748), .B2(n25192), .C1(n9005), .C2(n25186), .A(
        n22290), .ZN(n22283) );
  NAND2_X1 U23619 ( .A1(n22255), .A2(n22256), .ZN(n5401) );
  NOR4_X1 U23620 ( .A1(n22265), .A2(n22266), .A3(n22267), .A4(n22268), .ZN(
        n22255) );
  NOR4_X1 U23621 ( .A1(n22257), .A2(n22258), .A3(n22259), .A4(n22260), .ZN(
        n22256) );
  OAI221_X1 U23622 ( .B1(n20747), .B2(n25192), .C1(n9004), .C2(n25186), .A(
        n22272), .ZN(n22265) );
  NAND2_X1 U23623 ( .A1(n22237), .A2(n22238), .ZN(n5402) );
  NOR4_X1 U23624 ( .A1(n22247), .A2(n22248), .A3(n22249), .A4(n22250), .ZN(
        n22237) );
  NOR4_X1 U23625 ( .A1(n22239), .A2(n22240), .A3(n22241), .A4(n22242), .ZN(
        n22238) );
  OAI221_X1 U23626 ( .B1(n20746), .B2(n25192), .C1(n9003), .C2(n25186), .A(
        n22254), .ZN(n22247) );
  NAND2_X1 U23627 ( .A1(n22219), .A2(n22220), .ZN(n5403) );
  NOR4_X1 U23628 ( .A1(n22229), .A2(n22230), .A3(n22231), .A4(n22232), .ZN(
        n22219) );
  NOR4_X1 U23629 ( .A1(n22221), .A2(n22222), .A3(n22223), .A4(n22224), .ZN(
        n22220) );
  OAI221_X1 U23630 ( .B1(n20745), .B2(n25192), .C1(n9002), .C2(n25186), .A(
        n22236), .ZN(n22229) );
  NAND2_X1 U23631 ( .A1(n22201), .A2(n22202), .ZN(n5404) );
  NOR4_X1 U23632 ( .A1(n22211), .A2(n22212), .A3(n22213), .A4(n22214), .ZN(
        n22201) );
  NOR4_X1 U23633 ( .A1(n22203), .A2(n22204), .A3(n22205), .A4(n22206), .ZN(
        n22202) );
  OAI221_X1 U23634 ( .B1(n20744), .B2(n25192), .C1(n9001), .C2(n25186), .A(
        n22218), .ZN(n22211) );
  NAND2_X1 U23635 ( .A1(n22183), .A2(n22184), .ZN(n5405) );
  NOR4_X1 U23636 ( .A1(n22193), .A2(n22194), .A3(n22195), .A4(n22196), .ZN(
        n22183) );
  NOR4_X1 U23637 ( .A1(n22185), .A2(n22186), .A3(n22187), .A4(n22188), .ZN(
        n22184) );
  OAI221_X1 U23638 ( .B1(n20743), .B2(n25192), .C1(n9000), .C2(n25186), .A(
        n22200), .ZN(n22193) );
  NAND2_X1 U23639 ( .A1(n22165), .A2(n22166), .ZN(n5406) );
  NOR4_X1 U23640 ( .A1(n22175), .A2(n22176), .A3(n22177), .A4(n22178), .ZN(
        n22165) );
  NOR4_X1 U23641 ( .A1(n22167), .A2(n22168), .A3(n22169), .A4(n22170), .ZN(
        n22166) );
  OAI221_X1 U23642 ( .B1(n20742), .B2(n25192), .C1(n8999), .C2(n25186), .A(
        n22182), .ZN(n22175) );
  NAND2_X1 U23643 ( .A1(n22147), .A2(n22148), .ZN(n5407) );
  NOR4_X1 U23644 ( .A1(n22157), .A2(n22158), .A3(n22159), .A4(n22160), .ZN(
        n22147) );
  NOR4_X1 U23645 ( .A1(n22149), .A2(n22150), .A3(n22151), .A4(n22152), .ZN(
        n22148) );
  OAI221_X1 U23646 ( .B1(n20741), .B2(n25192), .C1(n8998), .C2(n25186), .A(
        n22164), .ZN(n22157) );
  NAND2_X1 U23647 ( .A1(n22129), .A2(n22130), .ZN(n5408) );
  NOR4_X1 U23648 ( .A1(n22139), .A2(n22140), .A3(n22141), .A4(n22142), .ZN(
        n22129) );
  NOR4_X1 U23649 ( .A1(n22131), .A2(n22132), .A3(n22133), .A4(n22134), .ZN(
        n22130) );
  OAI221_X1 U23650 ( .B1(n20740), .B2(n25192), .C1(n8997), .C2(n25186), .A(
        n22146), .ZN(n22139) );
  NAND2_X1 U23651 ( .A1(n22111), .A2(n22112), .ZN(n5409) );
  NOR4_X1 U23652 ( .A1(n22121), .A2(n22122), .A3(n22123), .A4(n22124), .ZN(
        n22111) );
  NOR4_X1 U23653 ( .A1(n22113), .A2(n22114), .A3(n22115), .A4(n22116), .ZN(
        n22112) );
  OAI221_X1 U23654 ( .B1(n20739), .B2(n25192), .C1(n8996), .C2(n25186), .A(
        n22128), .ZN(n22121) );
  NAND2_X1 U23655 ( .A1(n22093), .A2(n22094), .ZN(n5410) );
  NOR4_X1 U23656 ( .A1(n22103), .A2(n22104), .A3(n22105), .A4(n22106), .ZN(
        n22093) );
  NOR4_X1 U23657 ( .A1(n22095), .A2(n22096), .A3(n22097), .A4(n22098), .ZN(
        n22094) );
  OAI221_X1 U23658 ( .B1(n20738), .B2(n25192), .C1(n8995), .C2(n25186), .A(
        n22110), .ZN(n22103) );
  NAND2_X1 U23659 ( .A1(n22075), .A2(n22076), .ZN(n5411) );
  NOR4_X1 U23660 ( .A1(n22085), .A2(n22086), .A3(n22087), .A4(n22088), .ZN(
        n22075) );
  NOR4_X1 U23661 ( .A1(n22077), .A2(n22078), .A3(n22079), .A4(n22080), .ZN(
        n22076) );
  OAI221_X1 U23662 ( .B1(n20737), .B2(n25193), .C1(n8994), .C2(n25187), .A(
        n22092), .ZN(n22085) );
  NAND2_X1 U23663 ( .A1(n22057), .A2(n22058), .ZN(n5412) );
  NOR4_X1 U23664 ( .A1(n22067), .A2(n22068), .A3(n22069), .A4(n22070), .ZN(
        n22057) );
  NOR4_X1 U23665 ( .A1(n22059), .A2(n22060), .A3(n22061), .A4(n22062), .ZN(
        n22058) );
  OAI221_X1 U23666 ( .B1(n20736), .B2(n25193), .C1(n8993), .C2(n25187), .A(
        n22074), .ZN(n22067) );
  NAND2_X1 U23667 ( .A1(n22039), .A2(n22040), .ZN(n5413) );
  NOR4_X1 U23668 ( .A1(n22049), .A2(n22050), .A3(n22051), .A4(n22052), .ZN(
        n22039) );
  NOR4_X1 U23669 ( .A1(n22041), .A2(n22042), .A3(n22043), .A4(n22044), .ZN(
        n22040) );
  OAI221_X1 U23670 ( .B1(n20735), .B2(n25193), .C1(n8992), .C2(n25187), .A(
        n22056), .ZN(n22049) );
  NAND2_X1 U23671 ( .A1(n22021), .A2(n22022), .ZN(n5414) );
  NOR4_X1 U23672 ( .A1(n22031), .A2(n22032), .A3(n22033), .A4(n22034), .ZN(
        n22021) );
  NOR4_X1 U23673 ( .A1(n22023), .A2(n22024), .A3(n22025), .A4(n22026), .ZN(
        n22022) );
  OAI221_X1 U23674 ( .B1(n20734), .B2(n25193), .C1(n8991), .C2(n25187), .A(
        n22038), .ZN(n22031) );
  NAND2_X1 U23675 ( .A1(n22003), .A2(n22004), .ZN(n5415) );
  NOR4_X1 U23676 ( .A1(n22013), .A2(n22014), .A3(n22015), .A4(n22016), .ZN(
        n22003) );
  NOR4_X1 U23677 ( .A1(n22005), .A2(n22006), .A3(n22007), .A4(n22008), .ZN(
        n22004) );
  OAI221_X1 U23678 ( .B1(n20733), .B2(n25193), .C1(n8990), .C2(n25187), .A(
        n22020), .ZN(n22013) );
  NAND2_X1 U23679 ( .A1(n21985), .A2(n21986), .ZN(n5416) );
  NOR4_X1 U23680 ( .A1(n21995), .A2(n21996), .A3(n21997), .A4(n21998), .ZN(
        n21985) );
  NOR4_X1 U23681 ( .A1(n21987), .A2(n21988), .A3(n21989), .A4(n21990), .ZN(
        n21986) );
  OAI221_X1 U23682 ( .B1(n20732), .B2(n25193), .C1(n8989), .C2(n25187), .A(
        n22002), .ZN(n21995) );
  NAND2_X1 U23683 ( .A1(n21967), .A2(n21968), .ZN(n5417) );
  NOR4_X1 U23684 ( .A1(n21977), .A2(n21978), .A3(n21979), .A4(n21980), .ZN(
        n21967) );
  NOR4_X1 U23685 ( .A1(n21969), .A2(n21970), .A3(n21971), .A4(n21972), .ZN(
        n21968) );
  OAI221_X1 U23686 ( .B1(n20731), .B2(n25193), .C1(n8988), .C2(n25187), .A(
        n21984), .ZN(n21977) );
  NAND2_X1 U23687 ( .A1(n21949), .A2(n21950), .ZN(n5418) );
  NOR4_X1 U23688 ( .A1(n21959), .A2(n21960), .A3(n21961), .A4(n21962), .ZN(
        n21949) );
  NOR4_X1 U23689 ( .A1(n21951), .A2(n21952), .A3(n21953), .A4(n21954), .ZN(
        n21950) );
  OAI221_X1 U23690 ( .B1(n20730), .B2(n25193), .C1(n8987), .C2(n25187), .A(
        n21966), .ZN(n21959) );
  NAND2_X1 U23691 ( .A1(n21931), .A2(n21932), .ZN(n5419) );
  NOR4_X1 U23692 ( .A1(n21941), .A2(n21942), .A3(n21943), .A4(n21944), .ZN(
        n21931) );
  NOR4_X1 U23693 ( .A1(n21933), .A2(n21934), .A3(n21935), .A4(n21936), .ZN(
        n21932) );
  OAI221_X1 U23694 ( .B1(n20729), .B2(n25193), .C1(n8986), .C2(n25187), .A(
        n21948), .ZN(n21941) );
  NAND2_X1 U23695 ( .A1(n21913), .A2(n21914), .ZN(n5420) );
  NOR4_X1 U23696 ( .A1(n21923), .A2(n21924), .A3(n21925), .A4(n21926), .ZN(
        n21913) );
  NOR4_X1 U23697 ( .A1(n21915), .A2(n21916), .A3(n21917), .A4(n21918), .ZN(
        n21914) );
  OAI221_X1 U23698 ( .B1(n20728), .B2(n25193), .C1(n8985), .C2(n25187), .A(
        n21930), .ZN(n21923) );
  NAND2_X1 U23699 ( .A1(n21895), .A2(n21896), .ZN(n5421) );
  NOR4_X1 U23700 ( .A1(n21905), .A2(n21906), .A3(n21907), .A4(n21908), .ZN(
        n21895) );
  NOR4_X1 U23701 ( .A1(n21897), .A2(n21898), .A3(n21899), .A4(n21900), .ZN(
        n21896) );
  OAI221_X1 U23702 ( .B1(n20727), .B2(n25193), .C1(n8984), .C2(n25187), .A(
        n21912), .ZN(n21905) );
  NAND2_X1 U23703 ( .A1(n21877), .A2(n21878), .ZN(n5422) );
  NOR4_X1 U23704 ( .A1(n21887), .A2(n21888), .A3(n21889), .A4(n21890), .ZN(
        n21877) );
  NOR4_X1 U23705 ( .A1(n21879), .A2(n21880), .A3(n21881), .A4(n21882), .ZN(
        n21878) );
  OAI221_X1 U23706 ( .B1(n20726), .B2(n25193), .C1(n8983), .C2(n25187), .A(
        n21894), .ZN(n21887) );
  NAND2_X1 U23707 ( .A1(n21859), .A2(n21860), .ZN(n5423) );
  NOR4_X1 U23708 ( .A1(n21869), .A2(n21870), .A3(n21871), .A4(n21872), .ZN(
        n21859) );
  NOR4_X1 U23709 ( .A1(n21861), .A2(n21862), .A3(n21863), .A4(n21864), .ZN(
        n21860) );
  OAI221_X1 U23710 ( .B1(n20725), .B2(n25194), .C1(n8982), .C2(n25188), .A(
        n21876), .ZN(n21869) );
  NAND2_X1 U23711 ( .A1(n21841), .A2(n21842), .ZN(n5424) );
  NOR4_X1 U23712 ( .A1(n21851), .A2(n21852), .A3(n21853), .A4(n21854), .ZN(
        n21841) );
  NOR4_X1 U23713 ( .A1(n21843), .A2(n21844), .A3(n21845), .A4(n21846), .ZN(
        n21842) );
  OAI221_X1 U23714 ( .B1(n20724), .B2(n25194), .C1(n8981), .C2(n25188), .A(
        n21858), .ZN(n21851) );
  NAND2_X1 U23715 ( .A1(n21823), .A2(n21824), .ZN(n5425) );
  NOR4_X1 U23716 ( .A1(n21833), .A2(n21834), .A3(n21835), .A4(n21836), .ZN(
        n21823) );
  NOR4_X1 U23717 ( .A1(n21825), .A2(n21826), .A3(n21827), .A4(n21828), .ZN(
        n21824) );
  OAI221_X1 U23718 ( .B1(n20723), .B2(n25194), .C1(n8980), .C2(n25188), .A(
        n21840), .ZN(n21833) );
  NAND2_X1 U23719 ( .A1(n21805), .A2(n21806), .ZN(n5426) );
  NOR4_X1 U23720 ( .A1(n21815), .A2(n21816), .A3(n21817), .A4(n21818), .ZN(
        n21805) );
  NOR4_X1 U23721 ( .A1(n21807), .A2(n21808), .A3(n21809), .A4(n21810), .ZN(
        n21806) );
  OAI221_X1 U23722 ( .B1(n20722), .B2(n25194), .C1(n8979), .C2(n25188), .A(
        n21822), .ZN(n21815) );
  NAND2_X1 U23723 ( .A1(n21787), .A2(n21788), .ZN(n5427) );
  NOR4_X1 U23724 ( .A1(n21797), .A2(n21798), .A3(n21799), .A4(n21800), .ZN(
        n21787) );
  NOR4_X1 U23725 ( .A1(n21789), .A2(n21790), .A3(n21791), .A4(n21792), .ZN(
        n21788) );
  OAI221_X1 U23726 ( .B1(n20721), .B2(n25194), .C1(n8978), .C2(n25188), .A(
        n21804), .ZN(n21797) );
  NAND2_X1 U23727 ( .A1(n21769), .A2(n21770), .ZN(n5428) );
  NOR4_X1 U23728 ( .A1(n21779), .A2(n21780), .A3(n21781), .A4(n21782), .ZN(
        n21769) );
  NOR4_X1 U23729 ( .A1(n21771), .A2(n21772), .A3(n21773), .A4(n21774), .ZN(
        n21770) );
  OAI221_X1 U23730 ( .B1(n20720), .B2(n25194), .C1(n8977), .C2(n25188), .A(
        n21786), .ZN(n21779) );
  NAND2_X1 U23731 ( .A1(n21751), .A2(n21752), .ZN(n5429) );
  NOR4_X1 U23732 ( .A1(n21761), .A2(n21762), .A3(n21763), .A4(n21764), .ZN(
        n21751) );
  NOR4_X1 U23733 ( .A1(n21753), .A2(n21754), .A3(n21755), .A4(n21756), .ZN(
        n21752) );
  OAI221_X1 U23734 ( .B1(n20719), .B2(n25194), .C1(n8976), .C2(n25188), .A(
        n21768), .ZN(n21761) );
  NAND2_X1 U23735 ( .A1(n21733), .A2(n21734), .ZN(n5430) );
  NOR4_X1 U23736 ( .A1(n21743), .A2(n21744), .A3(n21745), .A4(n21746), .ZN(
        n21733) );
  NOR4_X1 U23737 ( .A1(n21735), .A2(n21736), .A3(n21737), .A4(n21738), .ZN(
        n21734) );
  OAI221_X1 U23738 ( .B1(n20718), .B2(n25194), .C1(n8975), .C2(n25188), .A(
        n21750), .ZN(n21743) );
  NAND2_X1 U23739 ( .A1(n21715), .A2(n21716), .ZN(n5431) );
  NOR4_X1 U23740 ( .A1(n21725), .A2(n21726), .A3(n21727), .A4(n21728), .ZN(
        n21715) );
  NOR4_X1 U23741 ( .A1(n21717), .A2(n21718), .A3(n21719), .A4(n21720), .ZN(
        n21716) );
  OAI221_X1 U23742 ( .B1(n20717), .B2(n25194), .C1(n8974), .C2(n25188), .A(
        n21732), .ZN(n21725) );
  NAND2_X1 U23743 ( .A1(n21697), .A2(n21698), .ZN(n5432) );
  NOR4_X1 U23744 ( .A1(n21707), .A2(n21708), .A3(n21709), .A4(n21710), .ZN(
        n21697) );
  NOR4_X1 U23745 ( .A1(n21699), .A2(n21700), .A3(n21701), .A4(n21702), .ZN(
        n21698) );
  OAI221_X1 U23746 ( .B1(n20716), .B2(n25194), .C1(n8973), .C2(n25188), .A(
        n21714), .ZN(n21707) );
  NAND2_X1 U23747 ( .A1(n21679), .A2(n21680), .ZN(n5433) );
  NOR4_X1 U23748 ( .A1(n21689), .A2(n21690), .A3(n21691), .A4(n21692), .ZN(
        n21679) );
  NOR4_X1 U23749 ( .A1(n21681), .A2(n21682), .A3(n21683), .A4(n21684), .ZN(
        n21680) );
  OAI221_X1 U23750 ( .B1(n20715), .B2(n25194), .C1(n8972), .C2(n25188), .A(
        n21696), .ZN(n21689) );
  NAND2_X1 U23751 ( .A1(n21661), .A2(n21662), .ZN(n5434) );
  NOR4_X1 U23752 ( .A1(n21671), .A2(n21672), .A3(n21673), .A4(n21674), .ZN(
        n21661) );
  NOR4_X1 U23753 ( .A1(n21663), .A2(n21664), .A3(n21665), .A4(n21666), .ZN(
        n21662) );
  OAI221_X1 U23754 ( .B1(n20714), .B2(n25194), .C1(n8971), .C2(n25188), .A(
        n21678), .ZN(n21671) );
  OAI22_X1 U23755 ( .A1(n25597), .A2(n21477), .B1(n25782), .B2(n25589), .ZN(
        n6527) );
  OAI22_X1 U23756 ( .A1(n25597), .A2(n21476), .B1(n25785), .B2(n25589), .ZN(
        n6528) );
  OAI22_X1 U23757 ( .A1(n25597), .A2(n21475), .B1(n25788), .B2(n25589), .ZN(
        n6529) );
  OAI22_X1 U23758 ( .A1(n25597), .A2(n21474), .B1(n25791), .B2(n25589), .ZN(
        n6530) );
  OAI22_X1 U23759 ( .A1(n25597), .A2(n21473), .B1(n25794), .B2(n25589), .ZN(
        n6531) );
  OAI22_X1 U23760 ( .A1(n25597), .A2(n21472), .B1(n25797), .B2(n25589), .ZN(
        n6532) );
  OAI22_X1 U23761 ( .A1(n25597), .A2(n21471), .B1(n25800), .B2(n25589), .ZN(
        n6533) );
  OAI22_X1 U23762 ( .A1(n25597), .A2(n21470), .B1(n25803), .B2(n25589), .ZN(
        n6534) );
  OAI22_X1 U23763 ( .A1(n25597), .A2(n21469), .B1(n25806), .B2(n25589), .ZN(
        n6535) );
  OAI22_X1 U23764 ( .A1(n25597), .A2(n21468), .B1(n25809), .B2(n25589), .ZN(
        n6536) );
  OAI22_X1 U23765 ( .A1(n25597), .A2(n21467), .B1(n25812), .B2(n25589), .ZN(
        n6537) );
  OAI22_X1 U23766 ( .A1(n25597), .A2(n21466), .B1(n25815), .B2(n25589), .ZN(
        n6538) );
  OAI22_X1 U23767 ( .A1(n25598), .A2(n21465), .B1(n25818), .B2(n25590), .ZN(
        n6539) );
  OAI22_X1 U23768 ( .A1(n25598), .A2(n21464), .B1(n25821), .B2(n25590), .ZN(
        n6540) );
  OAI22_X1 U23769 ( .A1(n25598), .A2(n21463), .B1(n25824), .B2(n25590), .ZN(
        n6541) );
  OAI22_X1 U23770 ( .A1(n25598), .A2(n21462), .B1(n25827), .B2(n25590), .ZN(
        n6542) );
  OAI22_X1 U23771 ( .A1(n25598), .A2(n21461), .B1(n25830), .B2(n25590), .ZN(
        n6543) );
  OAI22_X1 U23772 ( .A1(n25598), .A2(n21460), .B1(n25833), .B2(n25590), .ZN(
        n6544) );
  OAI22_X1 U23773 ( .A1(n25598), .A2(n21459), .B1(n25836), .B2(n25590), .ZN(
        n6545) );
  OAI22_X1 U23774 ( .A1(n25598), .A2(n21458), .B1(n25839), .B2(n25590), .ZN(
        n6546) );
  OAI22_X1 U23775 ( .A1(n25598), .A2(n21457), .B1(n25842), .B2(n25590), .ZN(
        n6547) );
  OAI22_X1 U23776 ( .A1(n25598), .A2(n21456), .B1(n25845), .B2(n25590), .ZN(
        n6548) );
  OAI22_X1 U23777 ( .A1(n25598), .A2(n21455), .B1(n25848), .B2(n25590), .ZN(
        n6549) );
  OAI22_X1 U23778 ( .A1(n25598), .A2(n21454), .B1(n25851), .B2(n25590), .ZN(
        n6550) );
  OAI22_X1 U23779 ( .A1(n25598), .A2(n21453), .B1(n25854), .B2(n25591), .ZN(
        n6551) );
  OAI22_X1 U23780 ( .A1(n25599), .A2(n21452), .B1(n25857), .B2(n25591), .ZN(
        n6552) );
  OAI22_X1 U23781 ( .A1(n25599), .A2(n21451), .B1(n25860), .B2(n25591), .ZN(
        n6553) );
  OAI22_X1 U23782 ( .A1(n25599), .A2(n21450), .B1(n25863), .B2(n25591), .ZN(
        n6554) );
  OAI22_X1 U23783 ( .A1(n25599), .A2(n21449), .B1(n25866), .B2(n25591), .ZN(
        n6555) );
  OAI22_X1 U23784 ( .A1(n25599), .A2(n21448), .B1(n25869), .B2(n25591), .ZN(
        n6556) );
  OAI22_X1 U23785 ( .A1(n25599), .A2(n21447), .B1(n25872), .B2(n25591), .ZN(
        n6557) );
  OAI22_X1 U23786 ( .A1(n25599), .A2(n21446), .B1(n25875), .B2(n25591), .ZN(
        n6558) );
  OAI22_X1 U23787 ( .A1(n25599), .A2(n21445), .B1(n25878), .B2(n25591), .ZN(
        n6559) );
  OAI22_X1 U23788 ( .A1(n25599), .A2(n21444), .B1(n25881), .B2(n25591), .ZN(
        n6560) );
  OAI22_X1 U23789 ( .A1(n25599), .A2(n21443), .B1(n25884), .B2(n25591), .ZN(
        n6561) );
  OAI22_X1 U23790 ( .A1(n25599), .A2(n21442), .B1(n25887), .B2(n25591), .ZN(
        n6562) );
  OAI22_X1 U23791 ( .A1(n25599), .A2(n21441), .B1(n25890), .B2(n25592), .ZN(
        n6563) );
  OAI22_X1 U23792 ( .A1(n25599), .A2(n21440), .B1(n25893), .B2(n25592), .ZN(
        n6564) );
  OAI22_X1 U23793 ( .A1(n25600), .A2(n21439), .B1(n25896), .B2(n25592), .ZN(
        n6565) );
  OAI22_X1 U23794 ( .A1(n25600), .A2(n21438), .B1(n25899), .B2(n25592), .ZN(
        n6566) );
  OAI22_X1 U23795 ( .A1(n25600), .A2(n21437), .B1(n25902), .B2(n25592), .ZN(
        n6567) );
  OAI22_X1 U23796 ( .A1(n25600), .A2(n21436), .B1(n25905), .B2(n25592), .ZN(
        n6568) );
  OAI22_X1 U23797 ( .A1(n25600), .A2(n21435), .B1(n25908), .B2(n25592), .ZN(
        n6569) );
  OAI22_X1 U23798 ( .A1(n25600), .A2(n21434), .B1(n25911), .B2(n25592), .ZN(
        n6570) );
  OAI22_X1 U23799 ( .A1(n25600), .A2(n21433), .B1(n25914), .B2(n25592), .ZN(
        n6571) );
  OAI22_X1 U23800 ( .A1(n25600), .A2(n21432), .B1(n25917), .B2(n25592), .ZN(
        n6572) );
  OAI22_X1 U23801 ( .A1(n25600), .A2(n21431), .B1(n25920), .B2(n25592), .ZN(
        n6573) );
  OAI22_X1 U23802 ( .A1(n25600), .A2(n21430), .B1(n25923), .B2(n25592), .ZN(
        n6574) );
  OAI22_X1 U23803 ( .A1(n25600), .A2(n21429), .B1(n25926), .B2(n25593), .ZN(
        n6575) );
  OAI22_X1 U23804 ( .A1(n25600), .A2(n21428), .B1(n25929), .B2(n25593), .ZN(
        n6576) );
  OAI22_X1 U23805 ( .A1(n25600), .A2(n21427), .B1(n25932), .B2(n25593), .ZN(
        n6577) );
  OAI22_X1 U23806 ( .A1(n25601), .A2(n21426), .B1(n25935), .B2(n25593), .ZN(
        n6578) );
  OAI22_X1 U23807 ( .A1(n25601), .A2(n21425), .B1(n25938), .B2(n25593), .ZN(
        n6579) );
  OAI22_X1 U23808 ( .A1(n25601), .A2(n21424), .B1(n25941), .B2(n25593), .ZN(
        n6580) );
  OAI22_X1 U23809 ( .A1(n25601), .A2(n21423), .B1(n25944), .B2(n25593), .ZN(
        n6581) );
  OAI22_X1 U23810 ( .A1(n25601), .A2(n21422), .B1(n25947), .B2(n25593), .ZN(
        n6582) );
  OAI22_X1 U23811 ( .A1(n25601), .A2(n21421), .B1(n25950), .B2(n25593), .ZN(
        n6583) );
  OAI22_X1 U23812 ( .A1(n25601), .A2(n21420), .B1(n25953), .B2(n25593), .ZN(
        n6584) );
  OAI22_X1 U23813 ( .A1(n25601), .A2(n21419), .B1(n25956), .B2(n25593), .ZN(
        n6585) );
  OAI22_X1 U23814 ( .A1(n25601), .A2(n21418), .B1(n25959), .B2(n25593), .ZN(
        n6586) );
  OAI22_X1 U23815 ( .A1(n25572), .A2(n20965), .B1(n25782), .B2(n25564), .ZN(
        n6399) );
  OAI22_X1 U23816 ( .A1(n25572), .A2(n20964), .B1(n25785), .B2(n25564), .ZN(
        n6400) );
  OAI22_X1 U23817 ( .A1(n25572), .A2(n20963), .B1(n25788), .B2(n25564), .ZN(
        n6401) );
  OAI22_X1 U23818 ( .A1(n25572), .A2(n20962), .B1(n25791), .B2(n25564), .ZN(
        n6402) );
  OAI22_X1 U23819 ( .A1(n25572), .A2(n20961), .B1(n25794), .B2(n25564), .ZN(
        n6403) );
  OAI22_X1 U23820 ( .A1(n25572), .A2(n20960), .B1(n25797), .B2(n25564), .ZN(
        n6404) );
  OAI22_X1 U23821 ( .A1(n25572), .A2(n20959), .B1(n25800), .B2(n25564), .ZN(
        n6405) );
  OAI22_X1 U23822 ( .A1(n25572), .A2(n20958), .B1(n25803), .B2(n25564), .ZN(
        n6406) );
  OAI22_X1 U23823 ( .A1(n25572), .A2(n20957), .B1(n25806), .B2(n25564), .ZN(
        n6407) );
  OAI22_X1 U23824 ( .A1(n25572), .A2(n20956), .B1(n25809), .B2(n25564), .ZN(
        n6408) );
  OAI22_X1 U23825 ( .A1(n25572), .A2(n20955), .B1(n25812), .B2(n25564), .ZN(
        n6409) );
  OAI22_X1 U23826 ( .A1(n25572), .A2(n20954), .B1(n25815), .B2(n25564), .ZN(
        n6410) );
  OAI22_X1 U23827 ( .A1(n25573), .A2(n20953), .B1(n25818), .B2(n25565), .ZN(
        n6411) );
  OAI22_X1 U23828 ( .A1(n25573), .A2(n20952), .B1(n25821), .B2(n25565), .ZN(
        n6412) );
  OAI22_X1 U23829 ( .A1(n25573), .A2(n20951), .B1(n25824), .B2(n25565), .ZN(
        n6413) );
  OAI22_X1 U23830 ( .A1(n25573), .A2(n20950), .B1(n25827), .B2(n25565), .ZN(
        n6414) );
  OAI22_X1 U23831 ( .A1(n25573), .A2(n20949), .B1(n25830), .B2(n25565), .ZN(
        n6415) );
  OAI22_X1 U23832 ( .A1(n25573), .A2(n20948), .B1(n25833), .B2(n25565), .ZN(
        n6416) );
  OAI22_X1 U23833 ( .A1(n25573), .A2(n20947), .B1(n25836), .B2(n25565), .ZN(
        n6417) );
  OAI22_X1 U23834 ( .A1(n25573), .A2(n20946), .B1(n25839), .B2(n25565), .ZN(
        n6418) );
  OAI22_X1 U23835 ( .A1(n25573), .A2(n20945), .B1(n25842), .B2(n25565), .ZN(
        n6419) );
  OAI22_X1 U23836 ( .A1(n25573), .A2(n20944), .B1(n25845), .B2(n25565), .ZN(
        n6420) );
  OAI22_X1 U23837 ( .A1(n25573), .A2(n20943), .B1(n25848), .B2(n25565), .ZN(
        n6421) );
  OAI22_X1 U23838 ( .A1(n25573), .A2(n20942), .B1(n25851), .B2(n25565), .ZN(
        n6422) );
  OAI22_X1 U23839 ( .A1(n25573), .A2(n20941), .B1(n25854), .B2(n25566), .ZN(
        n6423) );
  OAI22_X1 U23840 ( .A1(n25574), .A2(n20940), .B1(n25857), .B2(n25566), .ZN(
        n6424) );
  OAI22_X1 U23841 ( .A1(n25574), .A2(n20939), .B1(n25860), .B2(n25566), .ZN(
        n6425) );
  OAI22_X1 U23842 ( .A1(n25574), .A2(n20938), .B1(n25863), .B2(n25566), .ZN(
        n6426) );
  OAI22_X1 U23843 ( .A1(n25574), .A2(n20937), .B1(n25866), .B2(n25566), .ZN(
        n6427) );
  OAI22_X1 U23844 ( .A1(n25574), .A2(n20936), .B1(n25869), .B2(n25566), .ZN(
        n6428) );
  OAI22_X1 U23845 ( .A1(n25574), .A2(n20935), .B1(n25872), .B2(n25566), .ZN(
        n6429) );
  OAI22_X1 U23846 ( .A1(n25574), .A2(n20934), .B1(n25875), .B2(n25566), .ZN(
        n6430) );
  OAI22_X1 U23847 ( .A1(n25574), .A2(n20933), .B1(n25878), .B2(n25566), .ZN(
        n6431) );
  OAI22_X1 U23848 ( .A1(n25574), .A2(n20932), .B1(n25881), .B2(n25566), .ZN(
        n6432) );
  OAI22_X1 U23849 ( .A1(n25574), .A2(n20931), .B1(n25884), .B2(n25566), .ZN(
        n6433) );
  OAI22_X1 U23850 ( .A1(n25574), .A2(n20930), .B1(n25887), .B2(n25566), .ZN(
        n6434) );
  OAI22_X1 U23851 ( .A1(n25574), .A2(n20929), .B1(n25890), .B2(n25567), .ZN(
        n6435) );
  OAI22_X1 U23852 ( .A1(n25574), .A2(n20928), .B1(n25893), .B2(n25567), .ZN(
        n6436) );
  OAI22_X1 U23853 ( .A1(n25575), .A2(n20927), .B1(n25896), .B2(n25567), .ZN(
        n6437) );
  OAI22_X1 U23854 ( .A1(n25575), .A2(n20926), .B1(n25899), .B2(n25567), .ZN(
        n6438) );
  OAI22_X1 U23855 ( .A1(n25575), .A2(n20925), .B1(n25902), .B2(n25567), .ZN(
        n6439) );
  OAI22_X1 U23856 ( .A1(n25575), .A2(n20924), .B1(n25905), .B2(n25567), .ZN(
        n6440) );
  OAI22_X1 U23857 ( .A1(n25575), .A2(n20923), .B1(n25908), .B2(n25567), .ZN(
        n6441) );
  OAI22_X1 U23858 ( .A1(n25575), .A2(n20922), .B1(n25911), .B2(n25567), .ZN(
        n6442) );
  OAI22_X1 U23859 ( .A1(n25575), .A2(n20921), .B1(n25914), .B2(n25567), .ZN(
        n6443) );
  OAI22_X1 U23860 ( .A1(n25575), .A2(n20920), .B1(n25917), .B2(n25567), .ZN(
        n6444) );
  OAI22_X1 U23861 ( .A1(n25575), .A2(n20919), .B1(n25920), .B2(n25567), .ZN(
        n6445) );
  OAI22_X1 U23862 ( .A1(n25575), .A2(n20918), .B1(n25923), .B2(n25567), .ZN(
        n6446) );
  OAI22_X1 U23863 ( .A1(n25575), .A2(n20917), .B1(n25926), .B2(n25568), .ZN(
        n6447) );
  OAI22_X1 U23864 ( .A1(n25575), .A2(n20916), .B1(n25929), .B2(n25568), .ZN(
        n6448) );
  OAI22_X1 U23865 ( .A1(n25575), .A2(n20915), .B1(n25932), .B2(n25568), .ZN(
        n6449) );
  OAI22_X1 U23866 ( .A1(n25576), .A2(n20914), .B1(n25935), .B2(n25568), .ZN(
        n6450) );
  OAI22_X1 U23867 ( .A1(n25576), .A2(n20913), .B1(n25938), .B2(n25568), .ZN(
        n6451) );
  OAI22_X1 U23868 ( .A1(n25576), .A2(n20912), .B1(n25941), .B2(n25568), .ZN(
        n6452) );
  OAI22_X1 U23869 ( .A1(n25576), .A2(n20911), .B1(n25944), .B2(n25568), .ZN(
        n6453) );
  OAI22_X1 U23870 ( .A1(n25576), .A2(n20910), .B1(n25947), .B2(n25568), .ZN(
        n6454) );
  OAI22_X1 U23871 ( .A1(n25576), .A2(n20909), .B1(n25950), .B2(n25568), .ZN(
        n6455) );
  OAI22_X1 U23872 ( .A1(n25576), .A2(n20908), .B1(n25953), .B2(n25568), .ZN(
        n6456) );
  OAI22_X1 U23873 ( .A1(n25576), .A2(n20907), .B1(n25956), .B2(n25568), .ZN(
        n6457) );
  OAI22_X1 U23874 ( .A1(n25576), .A2(n20906), .B1(n25959), .B2(n25568), .ZN(
        n6458) );
  OAI22_X1 U23875 ( .A1(n25382), .A2(n20777), .B1(n25963), .B2(n25375), .ZN(
        n5499) );
  OAI22_X1 U23876 ( .A1(n25382), .A2(n20776), .B1(n25966), .B2(n25375), .ZN(
        n5500) );
  OAI22_X1 U23877 ( .A1(n25382), .A2(n20775), .B1(n25969), .B2(n25375), .ZN(
        n5501) );
  OAI22_X1 U23878 ( .A1(n25382), .A2(n20774), .B1(n25972), .B2(n25375), .ZN(
        n5502) );
  OAI22_X1 U23879 ( .A1(n25675), .A2(n19749), .B1(n25781), .B2(n25667), .ZN(
        n6911) );
  OAI22_X1 U23880 ( .A1(n25675), .A2(n19748), .B1(n25784), .B2(n25667), .ZN(
        n6912) );
  OAI22_X1 U23881 ( .A1(n25675), .A2(n19747), .B1(n25787), .B2(n25667), .ZN(
        n6913) );
  OAI22_X1 U23882 ( .A1(n25675), .A2(n19746), .B1(n25790), .B2(n25667), .ZN(
        n6914) );
  OAI22_X1 U23883 ( .A1(n25675), .A2(n19745), .B1(n25793), .B2(n25667), .ZN(
        n6915) );
  OAI22_X1 U23884 ( .A1(n25675), .A2(n19744), .B1(n25796), .B2(n25667), .ZN(
        n6916) );
  OAI22_X1 U23885 ( .A1(n25675), .A2(n19743), .B1(n25799), .B2(n25667), .ZN(
        n6917) );
  OAI22_X1 U23886 ( .A1(n25675), .A2(n19742), .B1(n25802), .B2(n25667), .ZN(
        n6918) );
  OAI22_X1 U23887 ( .A1(n25675), .A2(n19741), .B1(n25805), .B2(n25667), .ZN(
        n6919) );
  OAI22_X1 U23888 ( .A1(n25675), .A2(n19740), .B1(n25808), .B2(n25667), .ZN(
        n6920) );
  OAI22_X1 U23889 ( .A1(n25675), .A2(n19739), .B1(n25811), .B2(n25667), .ZN(
        n6921) );
  OAI22_X1 U23890 ( .A1(n25675), .A2(n19738), .B1(n25814), .B2(n25667), .ZN(
        n6922) );
  OAI22_X1 U23891 ( .A1(n25676), .A2(n19737), .B1(n25817), .B2(n25668), .ZN(
        n6923) );
  OAI22_X1 U23892 ( .A1(n25676), .A2(n19736), .B1(n25820), .B2(n25668), .ZN(
        n6924) );
  OAI22_X1 U23893 ( .A1(n25676), .A2(n19735), .B1(n25823), .B2(n25668), .ZN(
        n6925) );
  OAI22_X1 U23894 ( .A1(n25676), .A2(n19734), .B1(n25826), .B2(n25668), .ZN(
        n6926) );
  OAI22_X1 U23895 ( .A1(n25676), .A2(n19733), .B1(n25829), .B2(n25668), .ZN(
        n6927) );
  OAI22_X1 U23896 ( .A1(n25676), .A2(n19732), .B1(n25832), .B2(n25668), .ZN(
        n6928) );
  OAI22_X1 U23897 ( .A1(n25676), .A2(n19731), .B1(n25835), .B2(n25668), .ZN(
        n6929) );
  OAI22_X1 U23898 ( .A1(n25676), .A2(n19730), .B1(n25838), .B2(n25668), .ZN(
        n6930) );
  OAI22_X1 U23899 ( .A1(n25676), .A2(n19729), .B1(n25841), .B2(n25668), .ZN(
        n6931) );
  OAI22_X1 U23900 ( .A1(n25676), .A2(n19728), .B1(n25844), .B2(n25668), .ZN(
        n6932) );
  OAI22_X1 U23901 ( .A1(n25676), .A2(n19727), .B1(n25847), .B2(n25668), .ZN(
        n6933) );
  OAI22_X1 U23902 ( .A1(n25676), .A2(n19726), .B1(n25850), .B2(n25668), .ZN(
        n6934) );
  OAI22_X1 U23903 ( .A1(n25676), .A2(n19725), .B1(n25853), .B2(n25669), .ZN(
        n6935) );
  OAI22_X1 U23904 ( .A1(n25677), .A2(n19724), .B1(n25856), .B2(n25669), .ZN(
        n6936) );
  OAI22_X1 U23905 ( .A1(n25677), .A2(n19723), .B1(n25859), .B2(n25669), .ZN(
        n6937) );
  OAI22_X1 U23906 ( .A1(n25677), .A2(n19722), .B1(n25862), .B2(n25669), .ZN(
        n6938) );
  OAI22_X1 U23907 ( .A1(n25677), .A2(n19721), .B1(n25865), .B2(n25669), .ZN(
        n6939) );
  OAI22_X1 U23908 ( .A1(n25677), .A2(n19720), .B1(n25868), .B2(n25669), .ZN(
        n6940) );
  OAI22_X1 U23909 ( .A1(n25677), .A2(n19719), .B1(n25871), .B2(n25669), .ZN(
        n6941) );
  OAI22_X1 U23910 ( .A1(n25677), .A2(n19718), .B1(n25874), .B2(n25669), .ZN(
        n6942) );
  OAI22_X1 U23911 ( .A1(n25677), .A2(n19717), .B1(n25877), .B2(n25669), .ZN(
        n6943) );
  OAI22_X1 U23912 ( .A1(n25677), .A2(n19716), .B1(n25880), .B2(n25669), .ZN(
        n6944) );
  OAI22_X1 U23913 ( .A1(n25677), .A2(n19715), .B1(n25883), .B2(n25669), .ZN(
        n6945) );
  OAI22_X1 U23914 ( .A1(n25677), .A2(n19714), .B1(n25886), .B2(n25669), .ZN(
        n6946) );
  OAI22_X1 U23915 ( .A1(n25677), .A2(n19713), .B1(n25889), .B2(n25670), .ZN(
        n6947) );
  OAI22_X1 U23916 ( .A1(n25677), .A2(n19712), .B1(n25892), .B2(n25670), .ZN(
        n6948) );
  OAI22_X1 U23917 ( .A1(n25678), .A2(n19711), .B1(n25895), .B2(n25670), .ZN(
        n6949) );
  OAI22_X1 U23918 ( .A1(n25678), .A2(n19710), .B1(n25898), .B2(n25670), .ZN(
        n6950) );
  OAI22_X1 U23919 ( .A1(n25678), .A2(n19709), .B1(n25901), .B2(n25670), .ZN(
        n6951) );
  OAI22_X1 U23920 ( .A1(n25678), .A2(n19708), .B1(n25904), .B2(n25670), .ZN(
        n6952) );
  OAI22_X1 U23921 ( .A1(n25678), .A2(n19707), .B1(n25907), .B2(n25670), .ZN(
        n6953) );
  OAI22_X1 U23922 ( .A1(n25678), .A2(n19706), .B1(n25910), .B2(n25670), .ZN(
        n6954) );
  OAI22_X1 U23923 ( .A1(n25678), .A2(n19705), .B1(n25913), .B2(n25670), .ZN(
        n6955) );
  OAI22_X1 U23924 ( .A1(n25678), .A2(n19704), .B1(n25916), .B2(n25670), .ZN(
        n6956) );
  OAI22_X1 U23925 ( .A1(n25678), .A2(n19703), .B1(n25919), .B2(n25670), .ZN(
        n6957) );
  OAI22_X1 U23926 ( .A1(n25678), .A2(n19702), .B1(n25922), .B2(n25670), .ZN(
        n6958) );
  OAI22_X1 U23927 ( .A1(n25678), .A2(n19701), .B1(n25925), .B2(n25671), .ZN(
        n6959) );
  OAI22_X1 U23928 ( .A1(n25678), .A2(n19700), .B1(n25928), .B2(n25671), .ZN(
        n6960) );
  OAI22_X1 U23929 ( .A1(n25678), .A2(n19699), .B1(n25931), .B2(n25671), .ZN(
        n6961) );
  OAI22_X1 U23930 ( .A1(n25679), .A2(n19698), .B1(n25934), .B2(n25671), .ZN(
        n6962) );
  OAI22_X1 U23931 ( .A1(n25679), .A2(n19697), .B1(n25937), .B2(n25671), .ZN(
        n6963) );
  OAI22_X1 U23932 ( .A1(n25679), .A2(n19696), .B1(n25940), .B2(n25671), .ZN(
        n6964) );
  OAI22_X1 U23933 ( .A1(n25679), .A2(n19695), .B1(n25943), .B2(n25671), .ZN(
        n6965) );
  OAI22_X1 U23934 ( .A1(n25679), .A2(n19694), .B1(n25946), .B2(n25671), .ZN(
        n6966) );
  OAI22_X1 U23935 ( .A1(n25679), .A2(n19693), .B1(n25949), .B2(n25671), .ZN(
        n6967) );
  OAI22_X1 U23936 ( .A1(n25679), .A2(n19692), .B1(n25952), .B2(n25671), .ZN(
        n6968) );
  OAI22_X1 U23937 ( .A1(n25679), .A2(n19691), .B1(n25955), .B2(n25671), .ZN(
        n6969) );
  OAI22_X1 U23938 ( .A1(n25679), .A2(n19690), .B1(n25958), .B2(n25671), .ZN(
        n6970) );
  OAI22_X1 U23939 ( .A1(n25482), .A2(n21093), .B1(n25782), .B2(n25474), .ZN(
        n5951) );
  OAI22_X1 U23940 ( .A1(n25482), .A2(n21092), .B1(n25785), .B2(n25474), .ZN(
        n5952) );
  OAI22_X1 U23941 ( .A1(n25482), .A2(n21091), .B1(n25788), .B2(n25474), .ZN(
        n5953) );
  OAI22_X1 U23942 ( .A1(n25482), .A2(n21090), .B1(n25791), .B2(n25474), .ZN(
        n5954) );
  OAI22_X1 U23943 ( .A1(n25482), .A2(n21089), .B1(n25794), .B2(n25474), .ZN(
        n5955) );
  OAI22_X1 U23944 ( .A1(n25482), .A2(n21088), .B1(n25797), .B2(n25474), .ZN(
        n5956) );
  OAI22_X1 U23945 ( .A1(n25482), .A2(n21087), .B1(n25800), .B2(n25474), .ZN(
        n5957) );
  OAI22_X1 U23946 ( .A1(n25482), .A2(n21086), .B1(n25803), .B2(n25474), .ZN(
        n5958) );
  OAI22_X1 U23947 ( .A1(n25482), .A2(n21085), .B1(n25806), .B2(n25474), .ZN(
        n5959) );
  OAI22_X1 U23948 ( .A1(n25482), .A2(n21084), .B1(n25809), .B2(n25474), .ZN(
        n5960) );
  OAI22_X1 U23949 ( .A1(n25482), .A2(n21083), .B1(n25812), .B2(n25474), .ZN(
        n5961) );
  OAI22_X1 U23950 ( .A1(n25482), .A2(n21082), .B1(n25815), .B2(n25474), .ZN(
        n5962) );
  OAI22_X1 U23951 ( .A1(n25483), .A2(n21081), .B1(n25818), .B2(n25475), .ZN(
        n5963) );
  OAI22_X1 U23952 ( .A1(n25483), .A2(n21080), .B1(n25821), .B2(n25475), .ZN(
        n5964) );
  OAI22_X1 U23953 ( .A1(n25483), .A2(n21079), .B1(n25824), .B2(n25475), .ZN(
        n5965) );
  OAI22_X1 U23954 ( .A1(n25483), .A2(n21078), .B1(n25827), .B2(n25475), .ZN(
        n5966) );
  OAI22_X1 U23955 ( .A1(n25483), .A2(n21077), .B1(n25830), .B2(n25475), .ZN(
        n5967) );
  OAI22_X1 U23956 ( .A1(n25483), .A2(n21076), .B1(n25833), .B2(n25475), .ZN(
        n5968) );
  OAI22_X1 U23957 ( .A1(n25483), .A2(n21075), .B1(n25836), .B2(n25475), .ZN(
        n5969) );
  OAI22_X1 U23958 ( .A1(n25483), .A2(n21074), .B1(n25839), .B2(n25475), .ZN(
        n5970) );
  OAI22_X1 U23959 ( .A1(n25483), .A2(n21073), .B1(n25842), .B2(n25475), .ZN(
        n5971) );
  OAI22_X1 U23960 ( .A1(n25483), .A2(n21072), .B1(n25845), .B2(n25475), .ZN(
        n5972) );
  OAI22_X1 U23961 ( .A1(n25483), .A2(n21071), .B1(n25848), .B2(n25475), .ZN(
        n5973) );
  OAI22_X1 U23962 ( .A1(n25483), .A2(n21070), .B1(n25851), .B2(n25475), .ZN(
        n5974) );
  OAI22_X1 U23963 ( .A1(n25483), .A2(n21069), .B1(n25854), .B2(n25476), .ZN(
        n5975) );
  OAI22_X1 U23964 ( .A1(n25484), .A2(n21068), .B1(n25857), .B2(n25476), .ZN(
        n5976) );
  OAI22_X1 U23965 ( .A1(n25484), .A2(n21067), .B1(n25860), .B2(n25476), .ZN(
        n5977) );
  OAI22_X1 U23966 ( .A1(n25484), .A2(n21066), .B1(n25863), .B2(n25476), .ZN(
        n5978) );
  OAI22_X1 U23967 ( .A1(n25484), .A2(n21065), .B1(n25866), .B2(n25476), .ZN(
        n5979) );
  OAI22_X1 U23968 ( .A1(n25484), .A2(n21064), .B1(n25869), .B2(n25476), .ZN(
        n5980) );
  OAI22_X1 U23969 ( .A1(n25484), .A2(n21063), .B1(n25872), .B2(n25476), .ZN(
        n5981) );
  OAI22_X1 U23970 ( .A1(n25484), .A2(n21062), .B1(n25875), .B2(n25476), .ZN(
        n5982) );
  OAI22_X1 U23971 ( .A1(n25484), .A2(n21061), .B1(n25878), .B2(n25476), .ZN(
        n5983) );
  OAI22_X1 U23972 ( .A1(n25484), .A2(n21060), .B1(n25881), .B2(n25476), .ZN(
        n5984) );
  OAI22_X1 U23973 ( .A1(n25484), .A2(n21059), .B1(n25884), .B2(n25476), .ZN(
        n5985) );
  OAI22_X1 U23974 ( .A1(n25484), .A2(n21058), .B1(n25887), .B2(n25476), .ZN(
        n5986) );
  OAI22_X1 U23975 ( .A1(n25484), .A2(n21057), .B1(n25890), .B2(n25477), .ZN(
        n5987) );
  OAI22_X1 U23976 ( .A1(n25484), .A2(n21056), .B1(n25893), .B2(n25477), .ZN(
        n5988) );
  OAI22_X1 U23977 ( .A1(n25485), .A2(n21055), .B1(n25896), .B2(n25477), .ZN(
        n5989) );
  OAI22_X1 U23978 ( .A1(n25485), .A2(n21054), .B1(n25899), .B2(n25477), .ZN(
        n5990) );
  OAI22_X1 U23979 ( .A1(n25485), .A2(n21053), .B1(n25902), .B2(n25477), .ZN(
        n5991) );
  OAI22_X1 U23980 ( .A1(n25485), .A2(n21052), .B1(n25905), .B2(n25477), .ZN(
        n5992) );
  OAI22_X1 U23981 ( .A1(n25485), .A2(n21051), .B1(n25908), .B2(n25477), .ZN(
        n5993) );
  OAI22_X1 U23982 ( .A1(n25485), .A2(n21050), .B1(n25911), .B2(n25477), .ZN(
        n5994) );
  OAI22_X1 U23983 ( .A1(n25485), .A2(n21049), .B1(n25914), .B2(n25477), .ZN(
        n5995) );
  OAI22_X1 U23984 ( .A1(n25485), .A2(n21048), .B1(n25917), .B2(n25477), .ZN(
        n5996) );
  OAI22_X1 U23985 ( .A1(n25485), .A2(n21047), .B1(n25920), .B2(n25477), .ZN(
        n5997) );
  OAI22_X1 U23986 ( .A1(n25485), .A2(n21046), .B1(n25923), .B2(n25477), .ZN(
        n5998) );
  OAI22_X1 U23987 ( .A1(n25485), .A2(n21045), .B1(n25926), .B2(n25478), .ZN(
        n5999) );
  OAI22_X1 U23988 ( .A1(n25485), .A2(n21044), .B1(n25929), .B2(n25478), .ZN(
        n6000) );
  OAI22_X1 U23989 ( .A1(n25485), .A2(n21043), .B1(n25932), .B2(n25478), .ZN(
        n6001) );
  OAI22_X1 U23990 ( .A1(n25486), .A2(n21042), .B1(n25935), .B2(n25478), .ZN(
        n6002) );
  OAI22_X1 U23991 ( .A1(n25486), .A2(n21041), .B1(n25938), .B2(n25478), .ZN(
        n6003) );
  OAI22_X1 U23992 ( .A1(n25486), .A2(n21040), .B1(n25941), .B2(n25478), .ZN(
        n6004) );
  OAI22_X1 U23993 ( .A1(n25486), .A2(n21039), .B1(n25944), .B2(n25478), .ZN(
        n6005) );
  OAI22_X1 U23994 ( .A1(n25486), .A2(n21038), .B1(n25947), .B2(n25478), .ZN(
        n6006) );
  OAI22_X1 U23995 ( .A1(n25486), .A2(n21037), .B1(n25950), .B2(n25478), .ZN(
        n6007) );
  OAI22_X1 U23996 ( .A1(n25486), .A2(n21036), .B1(n25953), .B2(n25478), .ZN(
        n6008) );
  OAI22_X1 U23997 ( .A1(n25486), .A2(n21035), .B1(n25956), .B2(n25478), .ZN(
        n6009) );
  OAI22_X1 U23998 ( .A1(n25486), .A2(n21034), .B1(n25959), .B2(n25478), .ZN(
        n6010) );
  NOR3_X1 U23999 ( .A1(n19493), .A2(ADD_RD2[3]), .A3(n19489), .ZN(n23940) );
  NOR3_X1 U24000 ( .A1(n19488), .A2(ADD_RD1[3]), .A3(n19484), .ZN(n22743) );
  NOR3_X1 U24001 ( .A1(n19493), .A2(ADD_RD2[4]), .A3(n19490), .ZN(n23929) );
  NOR3_X1 U24002 ( .A1(n19488), .A2(ADD_RD1[4]), .A3(n19485), .ZN(n22732) );
  NOR3_X1 U24003 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n19493), .ZN(n23937)
         );
  NOR3_X1 U24004 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n19488), .ZN(n22740)
         );
  NOR3_X1 U24005 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(
        n23935) );
  NOR3_X1 U24006 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(
        n22738) );
  NOR3_X1 U24007 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n19489), .ZN(n23933)
         );
  NOR3_X1 U24008 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n19484), .ZN(n22736)
         );
  NOR3_X1 U24009 ( .A1(n19489), .A2(ADD_RD2[0]), .A3(n19490), .ZN(n23939) );
  NOR3_X1 U24010 ( .A1(n19484), .A2(ADD_RD1[0]), .A3(n19485), .ZN(n22742) );
  NOR3_X1 U24011 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n19490), .ZN(n23927)
         );
  NOR3_X1 U24012 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n19485), .ZN(n22730)
         );
  NAND2_X1 U24013 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .ZN(n21490) );
  NAND2_X1 U24014 ( .A1(ADD_WR[1]), .A2(n19483), .ZN(n21487) );
  NAND2_X1 U24015 ( .A1(ADD_WR[0]), .A2(n19482), .ZN(n21484) );
  INV_X1 U24016 ( .A(ADD_RD2[3]), .ZN(n19490) );
  INV_X1 U24017 ( .A(ADD_RD1[3]), .ZN(n19485) );
  INV_X1 U24018 ( .A(ADD_RD2[4]), .ZN(n19489) );
  INV_X1 U24019 ( .A(ADD_RD1[4]), .ZN(n19484) );
  INV_X1 U24020 ( .A(ADD_RD2[0]), .ZN(n19493) );
  INV_X1 U24021 ( .A(ADD_RD1[0]), .ZN(n19488) );
  AND3_X1 U24022 ( .A1(WR), .A2(ENABLE), .A3(ADD_WR[4]), .ZN(n21528) );
  AND3_X1 U24023 ( .A1(ENABLE), .A2(n19479), .A3(WR), .ZN(n21491) );
  INV_X1 U24024 ( .A(ADD_WR[4]), .ZN(n19479) );
  INV_X1 U24025 ( .A(RESET), .ZN(n19478) );
  INV_X1 U24026 ( .A(DATAIN[0]), .ZN(n19557) );
  INV_X1 U24027 ( .A(DATAIN[1]), .ZN(n19556) );
  INV_X1 U24028 ( .A(DATAIN[2]), .ZN(n19555) );
  INV_X1 U24029 ( .A(DATAIN[3]), .ZN(n19554) );
  INV_X1 U24030 ( .A(DATAIN[4]), .ZN(n19553) );
  INV_X1 U24031 ( .A(DATAIN[5]), .ZN(n19552) );
  INV_X1 U24032 ( .A(DATAIN[6]), .ZN(n19551) );
  INV_X1 U24033 ( .A(DATAIN[7]), .ZN(n19550) );
  INV_X1 U24034 ( .A(DATAIN[8]), .ZN(n19549) );
  INV_X1 U24035 ( .A(DATAIN[9]), .ZN(n19548) );
  INV_X1 U24036 ( .A(DATAIN[10]), .ZN(n19547) );
  INV_X1 U24037 ( .A(DATAIN[11]), .ZN(n19546) );
  INV_X1 U24038 ( .A(DATAIN[12]), .ZN(n19545) );
  INV_X1 U24039 ( .A(DATAIN[13]), .ZN(n19544) );
  INV_X1 U24040 ( .A(DATAIN[14]), .ZN(n19543) );
  INV_X1 U24041 ( .A(DATAIN[15]), .ZN(n19542) );
  INV_X1 U24042 ( .A(DATAIN[16]), .ZN(n19541) );
  INV_X1 U24043 ( .A(DATAIN[17]), .ZN(n19540) );
  INV_X1 U24044 ( .A(DATAIN[18]), .ZN(n19539) );
  INV_X1 U24045 ( .A(DATAIN[19]), .ZN(n19538) );
  INV_X1 U24046 ( .A(DATAIN[20]), .ZN(n19537) );
  INV_X1 U24047 ( .A(DATAIN[21]), .ZN(n19536) );
  INV_X1 U24048 ( .A(DATAIN[22]), .ZN(n19535) );
  INV_X1 U24049 ( .A(DATAIN[23]), .ZN(n19534) );
  INV_X1 U24050 ( .A(DATAIN[24]), .ZN(n19533) );
  INV_X1 U24051 ( .A(DATAIN[25]), .ZN(n19532) );
  INV_X1 U24052 ( .A(DATAIN[26]), .ZN(n19531) );
  INV_X1 U24053 ( .A(DATAIN[27]), .ZN(n19530) );
  INV_X1 U24054 ( .A(DATAIN[28]), .ZN(n19529) );
  INV_X1 U24055 ( .A(DATAIN[29]), .ZN(n19528) );
  INV_X1 U24056 ( .A(DATAIN[30]), .ZN(n19527) );
  INV_X1 U24057 ( .A(DATAIN[31]), .ZN(n19526) );
  INV_X1 U24058 ( .A(DATAIN[32]), .ZN(n19525) );
  INV_X1 U24059 ( .A(DATAIN[33]), .ZN(n19524) );
  INV_X1 U24060 ( .A(DATAIN[34]), .ZN(n19523) );
  INV_X1 U24061 ( .A(DATAIN[35]), .ZN(n19522) );
  INV_X1 U24062 ( .A(DATAIN[36]), .ZN(n19521) );
  INV_X1 U24063 ( .A(DATAIN[37]), .ZN(n19520) );
  INV_X1 U24064 ( .A(DATAIN[38]), .ZN(n19519) );
  INV_X1 U24065 ( .A(DATAIN[39]), .ZN(n19518) );
  INV_X1 U24066 ( .A(DATAIN[40]), .ZN(n19517) );
  INV_X1 U24067 ( .A(DATAIN[41]), .ZN(n19516) );
  INV_X1 U24068 ( .A(DATAIN[42]), .ZN(n19515) );
  INV_X1 U24069 ( .A(DATAIN[43]), .ZN(n19514) );
  INV_X1 U24070 ( .A(DATAIN[44]), .ZN(n19513) );
  INV_X1 U24071 ( .A(DATAIN[45]), .ZN(n19512) );
  INV_X1 U24072 ( .A(DATAIN[46]), .ZN(n19511) );
  INV_X1 U24073 ( .A(DATAIN[47]), .ZN(n19510) );
  INV_X1 U24074 ( .A(DATAIN[48]), .ZN(n19509) );
  INV_X1 U24075 ( .A(DATAIN[49]), .ZN(n19508) );
  INV_X1 U24076 ( .A(DATAIN[50]), .ZN(n19507) );
  INV_X1 U24077 ( .A(DATAIN[51]), .ZN(n19506) );
  INV_X1 U24078 ( .A(DATAIN[52]), .ZN(n19505) );
  INV_X1 U24079 ( .A(DATAIN[53]), .ZN(n19504) );
  INV_X1 U24080 ( .A(DATAIN[54]), .ZN(n19503) );
  INV_X1 U24081 ( .A(DATAIN[55]), .ZN(n19502) );
  INV_X1 U24082 ( .A(DATAIN[56]), .ZN(n19501) );
  INV_X1 U24083 ( .A(DATAIN[57]), .ZN(n19500) );
  INV_X1 U24084 ( .A(DATAIN[58]), .ZN(n19499) );
  INV_X1 U24085 ( .A(DATAIN[59]), .ZN(n19498) );
  INV_X1 U24086 ( .A(DATAIN[60]), .ZN(n19497) );
  INV_X1 U24087 ( .A(DATAIN[61]), .ZN(n19496) );
  INV_X1 U24088 ( .A(DATAIN[62]), .ZN(n19495) );
  INV_X1 U24089 ( .A(DATAIN[63]), .ZN(n19494) );
  INV_X1 U24090 ( .A(ADD_WR[3]), .ZN(n19480) );
  INV_X1 U24091 ( .A(ADD_WR[2]), .ZN(n19481) );
  INV_X1 U24092 ( .A(ADD_WR[0]), .ZN(n19483) );
  INV_X1 U24093 ( .A(ADD_RD2[2]), .ZN(n19491) );
  INV_X1 U24094 ( .A(ADD_RD1[2]), .ZN(n19486) );
  INV_X1 U24095 ( .A(ADD_RD2[1]), .ZN(n19492) );
  INV_X1 U24096 ( .A(ADD_RD1[1]), .ZN(n19487) );
  INV_X1 U24097 ( .A(ADD_WR[1]), .ZN(n19482) );
  CLKBUF_X1 U24098 ( .A(n22803), .Z(n24979) );
  CLKBUF_X1 U24099 ( .A(n22802), .Z(n24985) );
  CLKBUF_X1 U24100 ( .A(n22800), .Z(n24991) );
  CLKBUF_X1 U24101 ( .A(n22799), .Z(n24997) );
  CLKBUF_X1 U24102 ( .A(n22798), .Z(n25003) );
  CLKBUF_X1 U24103 ( .A(n22797), .Z(n25009) );
  CLKBUF_X1 U24104 ( .A(n22795), .Z(n25015) );
  CLKBUF_X1 U24105 ( .A(n22794), .Z(n25021) );
  CLKBUF_X1 U24106 ( .A(n22793), .Z(n25027) );
  CLKBUF_X1 U24107 ( .A(n22792), .Z(n25033) );
  CLKBUF_X1 U24108 ( .A(n22790), .Z(n25039) );
  CLKBUF_X1 U24109 ( .A(n22789), .Z(n25045) );
  CLKBUF_X1 U24110 ( .A(n22788), .Z(n25051) );
  CLKBUF_X1 U24111 ( .A(n22787), .Z(n25057) );
  CLKBUF_X1 U24112 ( .A(n22785), .Z(n25063) );
  CLKBUF_X1 U24113 ( .A(n22784), .Z(n25069) );
  CLKBUF_X1 U24114 ( .A(n22779), .Z(n25075) );
  CLKBUF_X1 U24115 ( .A(n22778), .Z(n25081) );
  CLKBUF_X1 U24116 ( .A(n22777), .Z(n25087) );
  CLKBUF_X1 U24117 ( .A(n22775), .Z(n25093) );
  CLKBUF_X1 U24118 ( .A(n22774), .Z(n25099) );
  CLKBUF_X1 U24119 ( .A(n22773), .Z(n25105) );
  CLKBUF_X1 U24120 ( .A(n22772), .Z(n25111) );
  CLKBUF_X1 U24121 ( .A(n22770), .Z(n25117) );
  CLKBUF_X1 U24122 ( .A(n22769), .Z(n25123) );
  CLKBUF_X1 U24123 ( .A(n22768), .Z(n25129) );
  CLKBUF_X1 U24124 ( .A(n22767), .Z(n25135) );
  CLKBUF_X1 U24125 ( .A(n22765), .Z(n25141) );
  CLKBUF_X1 U24126 ( .A(n22764), .Z(n25147) );
  CLKBUF_X1 U24127 ( .A(n22763), .Z(n25153) );
  CLKBUF_X1 U24128 ( .A(n22762), .Z(n25159) );
  CLKBUF_X1 U24129 ( .A(n22760), .Z(n25165) );
  CLKBUF_X1 U24130 ( .A(n22759), .Z(n25171) );
  CLKBUF_X1 U24131 ( .A(n21606), .Z(n25177) );
  CLKBUF_X1 U24132 ( .A(n21605), .Z(n25183) );
  CLKBUF_X1 U24133 ( .A(n21603), .Z(n25189) );
  CLKBUF_X1 U24134 ( .A(n21602), .Z(n25195) );
  CLKBUF_X1 U24135 ( .A(n21601), .Z(n25201) );
  CLKBUF_X1 U24136 ( .A(n21600), .Z(n25207) );
  CLKBUF_X1 U24137 ( .A(n21598), .Z(n25213) );
  CLKBUF_X1 U24138 ( .A(n21597), .Z(n25219) );
  CLKBUF_X1 U24139 ( .A(n21596), .Z(n25225) );
  CLKBUF_X1 U24140 ( .A(n21595), .Z(n25231) );
  CLKBUF_X1 U24141 ( .A(n21593), .Z(n25237) );
  CLKBUF_X1 U24142 ( .A(n21592), .Z(n25243) );
  CLKBUF_X1 U24143 ( .A(n21591), .Z(n25249) );
  CLKBUF_X1 U24144 ( .A(n21590), .Z(n25255) );
  CLKBUF_X1 U24145 ( .A(n21588), .Z(n25261) );
  CLKBUF_X1 U24146 ( .A(n21587), .Z(n25267) );
  CLKBUF_X1 U24147 ( .A(n21582), .Z(n25273) );
  CLKBUF_X1 U24148 ( .A(n21581), .Z(n25279) );
  CLKBUF_X1 U24149 ( .A(n21580), .Z(n25285) );
  CLKBUF_X1 U24150 ( .A(n21578), .Z(n25291) );
  CLKBUF_X1 U24151 ( .A(n21577), .Z(n25297) );
  CLKBUF_X1 U24152 ( .A(n21576), .Z(n25303) );
  CLKBUF_X1 U24153 ( .A(n21575), .Z(n25309) );
  CLKBUF_X1 U24154 ( .A(n21573), .Z(n25315) );
  CLKBUF_X1 U24155 ( .A(n21572), .Z(n25321) );
  CLKBUF_X1 U24156 ( .A(n21571), .Z(n25327) );
  CLKBUF_X1 U24157 ( .A(n21570), .Z(n25333) );
  CLKBUF_X1 U24158 ( .A(n21568), .Z(n25339) );
  CLKBUF_X1 U24159 ( .A(n21567), .Z(n25345) );
  CLKBUF_X1 U24160 ( .A(n21566), .Z(n25351) );
  CLKBUF_X1 U24161 ( .A(n21565), .Z(n25357) );
  CLKBUF_X1 U24162 ( .A(n21563), .Z(n25363) );
  CLKBUF_X1 U24163 ( .A(n21562), .Z(n25369) );
  CLKBUF_X1 U24164 ( .A(n21555), .Z(n25375) );
  CLKBUF_X1 U24165 ( .A(n21553), .Z(n25388) );
  CLKBUF_X1 U24166 ( .A(n21551), .Z(n25401) );
  CLKBUF_X1 U24167 ( .A(n21548), .Z(n25414) );
  CLKBUF_X1 U24168 ( .A(n21546), .Z(n25427) );
  CLKBUF_X1 U24169 ( .A(n21544), .Z(n25440) );
  CLKBUF_X1 U24170 ( .A(n21542), .Z(n25453) );
  CLKBUF_X1 U24171 ( .A(n21539), .Z(n25466) );
  CLKBUF_X1 U24172 ( .A(n21537), .Z(n25479) );
  CLKBUF_X1 U24173 ( .A(n21535), .Z(n25492) );
  CLKBUF_X1 U24174 ( .A(n21533), .Z(n25505) );
  CLKBUF_X1 U24175 ( .A(n21532), .Z(n25511) );
  CLKBUF_X1 U24176 ( .A(n21530), .Z(n25517) );
  CLKBUF_X1 U24177 ( .A(n21527), .Z(n25530) );
  CLKBUF_X1 U24178 ( .A(n21525), .Z(n25543) );
  CLKBUF_X1 U24179 ( .A(n21523), .Z(n25556) );
  CLKBUF_X1 U24180 ( .A(n21520), .Z(n25569) );
  CLKBUF_X1 U24181 ( .A(n21518), .Z(n25582) );
  CLKBUF_X1 U24182 ( .A(n21517), .Z(n25588) );
  CLKBUF_X1 U24183 ( .A(n21516), .Z(n25594) );
  CLKBUF_X1 U24184 ( .A(n21514), .Z(n25607) );
  CLKBUF_X1 U24185 ( .A(n21511), .Z(n25620) );
  CLKBUF_X1 U24186 ( .A(n21509), .Z(n25633) );
  CLKBUF_X1 U24187 ( .A(n21507), .Z(n25646) );
  CLKBUF_X1 U24188 ( .A(n21505), .Z(n25659) );
  CLKBUF_X1 U24189 ( .A(n21502), .Z(n25672) );
  CLKBUF_X1 U24190 ( .A(n21500), .Z(n25685) );
  CLKBUF_X1 U24191 ( .A(n21499), .Z(n25691) );
  CLKBUF_X1 U24192 ( .A(n21498), .Z(n25697) );
  CLKBUF_X1 U24193 ( .A(n21496), .Z(n25710) );
  CLKBUF_X1 U24194 ( .A(n21493), .Z(n25723) );
  CLKBUF_X1 U24195 ( .A(n21489), .Z(n25736) );
  CLKBUF_X1 U24196 ( .A(n21486), .Z(n25749) );
  CLKBUF_X1 U24197 ( .A(n21485), .Z(n25755) );
  CLKBUF_X1 U24198 ( .A(n21483), .Z(n25761) );
  CLKBUF_X1 U24199 ( .A(n21479), .Z(n25774) );
  CLKBUF_X1 U24200 ( .A(n21478), .Z(n25780) );
  CLKBUF_X1 U24201 ( .A(n19478), .Z(n25978) );
endmodule

