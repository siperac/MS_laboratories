
module Booth_Encoder_0 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n2, n3, n4, n5, n6;

  NAND2_X1 U3 ( .A1(i[1]), .A2(i[0]), .ZN(n2) );
  AND3_X1 U4 ( .A1(n5), .A2(n2), .A3(i[2]), .ZN(o[2]) );
  OAI21_X1 U5 ( .B1(i[1]), .B2(i[0]), .A(n2), .ZN(n4) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n2), .ZN(n5) );
  OAI21_X1 U7 ( .B1(i[1]), .B2(i[0]), .A(n2), .ZN(n3) );
  OAI22_X1 U8 ( .A1(n3), .A2(n6), .B1(i[2]), .B2(n2), .ZN(o[1]) );
  INV_X1 U9 ( .A(i[2]), .ZN(n6) );
  AOI21_X1 U10 ( .B1(n4), .B2(n2), .A(i[2]), .ZN(o[0]) );
endmodule


module MUX_booth_N64_0 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n3, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         net70125, net70123, net70121, net70119, net70129, net70127, net70137,
         net70133, net70151, net70149, net70145, net70175, net72882, net72880,
         net72879, net72878, net78774, net83777, net84586, net88405, net91117,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211;

  INV_X1 U1 ( .A(n142), .ZN(n139) );
  BUF_X1 U2 ( .A(n169), .Z(n142) );
  CLKBUF_X2 U3 ( .A(n8), .Z(net72880) );
  BUF_X2 U4 ( .A(net72878), .Z(n181) );
  BUF_X1 U5 ( .A(n182), .Z(net84586) );
  NAND2_X1 U6 ( .A1(n92), .A2(n93), .ZN(Y[29]) );
  NAND2_X1 U7 ( .A1(n98), .A2(n99), .ZN(Y[26]) );
  CLKBUF_X1 U8 ( .A(n193), .Z(n185) );
  BUF_X2 U9 ( .A(n193), .Z(n191) );
  BUF_X1 U10 ( .A(n5), .Z(n183) );
  NAND2_X1 U11 ( .A1(n46), .A2(n47), .ZN(Y[4]) );
  AND2_X2 U12 ( .A1(n176), .A2(n179), .ZN(n5) );
  INV_X1 U13 ( .A(E[4]), .ZN(n166) );
  CLKBUF_X1 U14 ( .A(n168), .Z(n140) );
  BUF_X2 U15 ( .A(net70145), .Z(net70149) );
  BUF_X1 U16 ( .A(sel[1]), .Z(n141) );
  BUF_X1 U17 ( .A(n184), .Z(n143) );
  BUF_X2 U18 ( .A(n183), .Z(net70129) );
  NAND2_X1 U19 ( .A1(D[29]), .A2(net70119), .ZN(n144) );
  NAND2_X1 U20 ( .A1(E[29]), .A2(net70133), .ZN(n145) );
  NAND2_X1 U21 ( .A1(B[29]), .A2(net91117), .ZN(n146) );
  AND3_X1 U22 ( .A1(n144), .A2(n145), .A3(n146), .ZN(n93) );
  NAND2_X1 U23 ( .A1(D[23]), .A2(net70119), .ZN(n147) );
  NAND2_X1 U24 ( .A1(E[23]), .A2(net70133), .ZN(n148) );
  NAND2_X1 U25 ( .A1(B[23]), .A2(net91117), .ZN(n149) );
  AND3_X1 U26 ( .A1(n147), .A2(n148), .A3(n149), .ZN(n105) );
  INV_X2 U27 ( .A(n180), .ZN(net70133) );
  AND2_X1 U28 ( .A1(D[14]), .A2(net70127), .ZN(n150) );
  AND2_X1 U29 ( .A1(E[14]), .A2(n143), .ZN(n151) );
  AND2_X1 U30 ( .A1(B[14]), .A2(net84586), .ZN(n152) );
  NOR3_X1 U31 ( .A1(n150), .A2(n151), .A3(n152), .ZN(n125) );
  BUF_X2 U32 ( .A(n5), .Z(net70127) );
  NOR4_X1 U33 ( .A1(net70145), .A2(n5), .A3(n8), .A4(n9), .ZN(n153) );
  NAND2_X1 U34 ( .A1(D[20]), .A2(net70119), .ZN(n154) );
  NAND2_X1 U35 ( .A1(E[20]), .A2(net70133), .ZN(n155) );
  NAND2_X1 U36 ( .A1(B[20]), .A2(net70151), .ZN(n156) );
  AND3_X1 U37 ( .A1(n154), .A2(n155), .A3(n156), .ZN(n111) );
  AND2_X1 U38 ( .A1(D[8]), .A2(net70125), .ZN(n157) );
  AND2_X1 U39 ( .A1(E[8]), .A2(n153), .ZN(n158) );
  AND2_X1 U40 ( .A1(B[8]), .A2(net70151), .ZN(n159) );
  NOR3_X1 U41 ( .A1(n158), .A2(n157), .A3(n159), .ZN(n11) );
  NAND2_X1 U42 ( .A1(D[22]), .A2(net70119), .ZN(n160) );
  NAND2_X1 U43 ( .A1(E[22]), .A2(net70133), .ZN(n161) );
  NAND2_X1 U44 ( .A1(B[22]), .A2(net91117), .ZN(n162) );
  AND3_X1 U45 ( .A1(n160), .A2(n161), .A3(n162), .ZN(n107) );
  AND2_X1 U46 ( .A1(D[5]), .A2(net70125), .ZN(n163) );
  AND2_X1 U47 ( .A1(net70137), .A2(E[5]), .ZN(n164) );
  AND2_X1 U48 ( .A1(B[5]), .A2(n182), .ZN(n165) );
  NOR3_X1 U49 ( .A1(n164), .A2(n163), .A3(n165), .ZN(n25) );
  NAND2_X1 U50 ( .A1(n175), .A2(n176), .ZN(n168) );
  NAND2_X1 U51 ( .A1(n172), .A2(n178), .ZN(n171) );
  NOR2_X1 U52 ( .A1(sel[0]), .A2(sel[1]), .ZN(n175) );
  NOR2_X1 U53 ( .A1(sel[0]), .A2(sel[2]), .ZN(n174) );
  NAND2_X1 U54 ( .A1(n141), .A2(n174), .ZN(n169) );
  NAND2_X1 U55 ( .A1(n173), .A2(n141), .ZN(n170) );
  NOR2_X1 U56 ( .A1(sel[2]), .A2(sel[1]), .ZN(n172) );
  INV_X1 U57 ( .A(n169), .ZN(n8) );
  INV_X2 U58 ( .A(n177), .ZN(net72882) );
  INV_X1 U59 ( .A(n181), .ZN(n177) );
  INV_X1 U60 ( .A(n171), .ZN(net70151) );
  NAND4_X1 U61 ( .A1(n170), .A2(n142), .A3(n168), .A4(n171), .ZN(n167) );
  INV_X1 U62 ( .A(n167), .ZN(net70137) );
  INV_X1 U63 ( .A(sel[2]), .ZN(n176) );
  AND2_X1 U64 ( .A1(n175), .A2(n176), .ZN(n9) );
  BUF_X1 U65 ( .A(sel[0]), .Z(n178) );
  AND2_X1 U66 ( .A1(n176), .A2(n178), .ZN(n173) );
  AND2_X1 U67 ( .A1(sel[0]), .A2(sel[1]), .ZN(n179) );
  INV_X1 U68 ( .A(n171), .ZN(net70145) );
  INV_X1 U69 ( .A(n171), .ZN(n182) );
  NOR2_X1 U70 ( .A1(n166), .A2(n167), .ZN(net83777) );
  INV_X4 U71 ( .A(n140), .ZN(net70175) );
  CLKBUF_X1 U72 ( .A(n167), .Z(n180) );
  BUF_X1 U73 ( .A(n139), .Z(net72879) );
  CLKBUF_X1 U74 ( .A(net70127), .Z(net70123) );
  CLKBUF_X1 U75 ( .A(net70129), .Z(net70121) );
  BUF_X2 U76 ( .A(n182), .Z(net91117) );
  NOR4_X1 U77 ( .A1(net70145), .A2(n5), .A3(n8), .A4(n9), .ZN(n184) );
  NAND2_X1 U78 ( .A1(n90), .A2(n91), .ZN(Y[2]) );
  CLKBUF_X1 U79 ( .A(net70151), .Z(net88405) );
  AND2_X1 U80 ( .A1(D[19]), .A2(net70125), .ZN(n186) );
  AND2_X1 U81 ( .A1(E[19]), .A2(n185), .ZN(n187) );
  AND2_X1 U82 ( .A1(B[19]), .A2(net84586), .ZN(n188) );
  NOR3_X1 U83 ( .A1(n186), .A2(n187), .A3(n188), .ZN(n115) );
  BUF_X2 U84 ( .A(n5), .Z(net70125) );
  NAND2_X1 U85 ( .A1(n130), .A2(n131), .ZN(Y[11]) );
  AND2_X1 U86 ( .A1(D[4]), .A2(net70127), .ZN(n189) );
  AND2_X1 U87 ( .A1(B[4]), .A2(net70145), .ZN(n190) );
  NOR3_X1 U88 ( .A1(n189), .A2(net83777), .A3(n190), .ZN(n47) );
  NAND2_X1 U89 ( .A1(n104), .A2(n105), .ZN(Y[23]) );
  AND2_X1 U90 ( .A1(n205), .A2(n203), .ZN(n192) );
  AND2_X1 U91 ( .A1(n204), .A2(n192), .ZN(n129) );
  NOR4_X1 U92 ( .A1(net70145), .A2(n5), .A3(n8), .A4(n9), .ZN(n193) );
  AND2_X1 U93 ( .A1(D[32]), .A2(net70121), .ZN(n194) );
  AND2_X1 U94 ( .A1(E[32]), .A2(n185), .ZN(n195) );
  AND2_X1 U95 ( .A1(B[32]), .A2(net70149), .ZN(n196) );
  NOR3_X1 U96 ( .A1(n194), .A2(n195), .A3(n196), .ZN(n85) );
  CLKBUF_X1 U97 ( .A(net70133), .Z(net78774) );
  NAND2_X1 U98 ( .A1(D[30]), .A2(net70119), .ZN(n197) );
  NAND2_X1 U99 ( .A1(E[30]), .A2(net70133), .ZN(n198) );
  NAND2_X1 U100 ( .A1(B[30]), .A2(net70151), .ZN(n199) );
  AND3_X1 U101 ( .A1(n197), .A2(n198), .A3(n199), .ZN(n89) );
  AOI222_X1 U102 ( .A1(D[11]), .A2(net70125), .B1(E[11]), .B2(n193), .C1(B[11]), .C2(net91117), .ZN(n131) );
  NAND2_X1 U103 ( .A1(n68), .A2(n69), .ZN(Y[3]) );
  NAND2_X1 U104 ( .A1(D[33]), .A2(net70121), .ZN(n200) );
  NAND2_X1 U105 ( .A1(E[33]), .A2(n185), .ZN(n201) );
  NAND2_X1 U106 ( .A1(B[33]), .A2(net70149), .ZN(n202) );
  AND3_X1 U107 ( .A1(n200), .A2(n201), .A3(n202), .ZN(n83) );
  NAND2_X1 U108 ( .A1(n96), .A2(n97), .ZN(Y[27]) );
  NAND2_X1 U109 ( .A1(n84), .A2(n85), .ZN(Y[32]) );
  NAND2_X1 U110 ( .A1(D[12]), .A2(net70129), .ZN(n203) );
  NAND2_X1 U111 ( .A1(E[12]), .A2(n153), .ZN(n204) );
  NAND2_X1 U112 ( .A1(B[12]), .A2(net70151), .ZN(n205) );
  AND2_X1 U113 ( .A1(D[31]), .A2(net70119), .ZN(n206) );
  AND2_X1 U114 ( .A1(E[31]), .A2(n185), .ZN(n207) );
  AND2_X1 U115 ( .A1(B[31]), .A2(net91117), .ZN(n208) );
  NOR3_X1 U116 ( .A1(n207), .A2(n206), .A3(n208), .ZN(n87) );
  BUF_X2 U117 ( .A(net70125), .Z(net70119) );
  NAND2_X1 U118 ( .A1(D[28]), .A2(net70119), .ZN(n209) );
  NAND2_X1 U119 ( .A1(E[28]), .A2(net70133), .ZN(n210) );
  NAND2_X1 U120 ( .A1(B[28]), .A2(net91117), .ZN(n211) );
  AND3_X1 U121 ( .A1(n209), .A2(n210), .A3(n211), .ZN(n95) );
  NAND2_X1 U122 ( .A1(n74), .A2(n75), .ZN(Y[37]) );
  AOI22_X1 U123 ( .A1(C[37]), .A2(net72882), .B1(A[37]), .B2(net70175), .ZN(
        n74) );
  AOI222_X1 U124 ( .A1(D[37]), .A2(net70121), .B1(E[37]), .B2(n185), .C1(B[37]), .C2(net88405), .ZN(n75) );
  AOI22_X1 U125 ( .A1(C[36]), .A2(net72879), .B1(A[36]), .B2(net70175), .ZN(
        n76) );
  NAND2_X1 U126 ( .A1(n82), .A2(n83), .ZN(Y[33]) );
  NAND2_X1 U127 ( .A1(n78), .A2(n79), .ZN(Y[35]) );
  AOI222_X1 U128 ( .A1(D[35]), .A2(net70121), .B1(E[35]), .B2(n191), .C1(B[35]), .C2(net88405), .ZN(n79) );
  NAND2_X1 U129 ( .A1(n70), .A2(n71), .ZN(Y[39]) );
  AOI22_X1 U130 ( .A1(C[39]), .A2(net72880), .B1(A[39]), .B2(net70175), .ZN(
        n70) );
  AOI222_X1 U131 ( .A1(D[39]), .A2(net70121), .B1(E[39]), .B2(n185), .C1(B[39]), .C2(net88405), .ZN(n71) );
  NAND2_X1 U132 ( .A1(n108), .A2(n109), .ZN(Y[21]) );
  AOI222_X1 U133 ( .A1(D[21]), .A2(net70119), .B1(E[21]), .B2(net70133), .C1(
        B[21]), .C2(net91117), .ZN(n109) );
  AOI22_X1 U134 ( .A1(C[21]), .A2(net72879), .B1(A[21]), .B2(net70175), .ZN(
        n108) );
  NAND2_X1 U135 ( .A1(n100), .A2(n101), .ZN(Y[25]) );
  AOI222_X1 U136 ( .A1(D[25]), .A2(net70119), .B1(E[25]), .B2(net70133), .C1(
        B[25]), .C2(net91117), .ZN(n101) );
  AOI22_X1 U137 ( .A1(C[25]), .A2(net72880), .B1(A[25]), .B2(net70175), .ZN(
        n100) );
  NAND2_X1 U138 ( .A1(n102), .A2(n103), .ZN(Y[24]) );
  AOI22_X1 U139 ( .A1(C[24]), .A2(net72882), .B1(A[24]), .B2(net70175), .ZN(
        n102) );
  AOI22_X1 U140 ( .A1(C[29]), .A2(net72882), .B1(A[29]), .B2(net70175), .ZN(
        n92) );
  NAND2_X1 U141 ( .A1(n129), .A2(n128), .ZN(Y[12]) );
  AOI22_X1 U142 ( .A1(C[12]), .A2(net72879), .B1(A[12]), .B2(net70175), .ZN(
        n128) );
  NAND2_X1 U143 ( .A1(n56), .A2(n57), .ZN(Y[45]) );
  AOI22_X1 U144 ( .A1(C[45]), .A2(net72879), .B1(A[45]), .B2(net70175), .ZN(
        n56) );
  AOI222_X1 U145 ( .A1(D[45]), .A2(net70123), .B1(E[45]), .B2(net78774), .C1(
        B[45]), .C2(net70151), .ZN(n57) );
  NAND2_X1 U146 ( .A1(n106), .A2(n107), .ZN(Y[22]) );
  AOI22_X1 U147 ( .A1(C[22]), .A2(net72882), .B1(A[22]), .B2(net70175), .ZN(
        n106) );
  NAND2_X1 U148 ( .A1(n72), .A2(n73), .ZN(Y[38]) );
  AOI22_X1 U149 ( .A1(C[38]), .A2(n181), .B1(A[38]), .B2(net70175), .ZN(n72)
         );
  AOI222_X1 U150 ( .A1(D[38]), .A2(net70121), .B1(E[38]), .B2(n185), .C1(B[38]), .C2(net70149), .ZN(n73) );
  NAND2_X1 U151 ( .A1(n58), .A2(n59), .ZN(Y[44]) );
  AOI22_X1 U152 ( .A1(C[44]), .A2(n181), .B1(A[44]), .B2(net70175), .ZN(n58)
         );
  AOI222_X1 U153 ( .A1(D[44]), .A2(net70123), .B1(E[44]), .B2(net78774), .C1(
        B[44]), .C2(net91117), .ZN(n59) );
  NAND2_X1 U154 ( .A1(n62), .A2(n63), .ZN(Y[42]) );
  AOI22_X1 U155 ( .A1(C[42]), .A2(net72879), .B1(A[42]), .B2(net70175), .ZN(
        n62) );
  AOI222_X1 U156 ( .A1(D[42]), .A2(net70121), .B1(E[42]), .B2(net78774), .C1(
        B[42]), .C2(net70149), .ZN(n63) );
  NAND2_X1 U157 ( .A1(n60), .A2(n61), .ZN(Y[43]) );
  AOI22_X1 U158 ( .A1(C[43]), .A2(net72882), .B1(A[43]), .B2(net70175), .ZN(
        n60) );
  AOI222_X1 U159 ( .A1(D[43]), .A2(net70121), .B1(E[43]), .B2(net78774), .C1(
        B[43]), .C2(net88405), .ZN(n61) );
  NAND2_X1 U160 ( .A1(n54), .A2(n55), .ZN(Y[46]) );
  AOI22_X1 U161 ( .A1(C[46]), .A2(net72880), .B1(A[46]), .B2(net70175), .ZN(
        n54) );
  AOI222_X1 U162 ( .A1(D[46]), .A2(net70123), .B1(E[46]), .B2(net78774), .C1(
        B[46]), .C2(net91117), .ZN(n55) );
  NAND2_X1 U163 ( .A1(n132), .A2(n133), .ZN(Y[10]) );
  AOI22_X1 U164 ( .A1(C[10]), .A2(n181), .B1(A[10]), .B2(net70175), .ZN(n132)
         );
  AOI222_X1 U165 ( .A1(D[10]), .A2(net70125), .B1(E[10]), .B2(n143), .C1(B[10]), .C2(net84586), .ZN(n133) );
  NAND2_X1 U166 ( .A1(n116), .A2(n117), .ZN(Y[18]) );
  AOI222_X1 U167 ( .A1(D[18]), .A2(net70127), .B1(E[18]), .B2(n185), .C1(B[18]), .C2(net84586), .ZN(n117) );
  AOI22_X1 U168 ( .A1(C[18]), .A2(n181), .B1(A[18]), .B2(net70175), .ZN(n116)
         );
  AOI22_X1 U169 ( .A1(C[26]), .A2(net72879), .B1(A[26]), .B2(net70175), .ZN(
        n98) );
  AOI222_X1 U170 ( .A1(D[26]), .A2(net70119), .B1(E[26]), .B2(net70133), .C1(
        B[26]), .C2(net91117), .ZN(n99) );
  NAND2_X1 U171 ( .A1(n52), .A2(n53), .ZN(Y[47]) );
  AOI22_X1 U172 ( .A1(C[47]), .A2(net72879), .B1(A[47]), .B2(net70175), .ZN(
        n52) );
  AOI222_X1 U173 ( .A1(D[47]), .A2(net70123), .B1(E[47]), .B2(net78774), .C1(
        B[47]), .C2(net91117), .ZN(n53) );
  NAND2_X1 U174 ( .A1(n66), .A2(n67), .ZN(Y[40]) );
  AOI22_X1 U175 ( .A1(C[40]), .A2(net72880), .B1(A[40]), .B2(net70175), .ZN(
        n66) );
  AOI222_X1 U176 ( .A1(D[40]), .A2(net70121), .B1(E[40]), .B2(n191), .C1(B[40]), .C2(net88405), .ZN(n67) );
  NAND2_X1 U177 ( .A1(n80), .A2(n81), .ZN(Y[34]) );
  AOI222_X1 U178 ( .A1(D[34]), .A2(net70121), .B1(E[34]), .B2(n191), .C1(B[34]), .C2(net88405), .ZN(n81) );
  NAND2_X1 U179 ( .A1(n64), .A2(n65), .ZN(Y[41]) );
  AOI22_X1 U180 ( .A1(C[41]), .A2(net72882), .B1(A[41]), .B2(net70175), .ZN(
        n64) );
  AOI222_X1 U181 ( .A1(D[41]), .A2(net70121), .B1(E[41]), .B2(n191), .C1(B[41]), .C2(net88405), .ZN(n65) );
  NAND2_X1 U182 ( .A1(n12), .A2(n13), .ZN(Y[7]) );
  AOI22_X1 U183 ( .A1(C[7]), .A2(net72878), .B1(A[7]), .B2(net70175), .ZN(n12)
         );
  AOI222_X1 U184 ( .A1(D[7]), .A2(net70129), .B1(n153), .B2(E[7]), .C1(B[7]), 
        .C2(n182), .ZN(n13) );
  AOI22_X1 U185 ( .A1(C[11]), .A2(net72879), .B1(A[11]), .B2(net70175), .ZN(
        n130) );
  NAND2_X1 U186 ( .A1(n122), .A2(n123), .ZN(Y[15]) );
  AOI222_X1 U187 ( .A1(D[15]), .A2(net70127), .B1(E[15]), .B2(n143), .C1(B[15]), .C2(net91117), .ZN(n123) );
  AOI22_X1 U188 ( .A1(C[15]), .A2(n181), .B1(A[15]), .B2(net70175), .ZN(n122)
         );
  NAND2_X1 U189 ( .A1(n114), .A2(n115), .ZN(Y[19]) );
  AOI22_X1 U190 ( .A1(C[19]), .A2(net72882), .B1(A[19]), .B2(net70175), .ZN(
        n114) );
  NAND2_X1 U191 ( .A1(n10), .A2(n11), .ZN(Y[8]) );
  AOI22_X1 U192 ( .A1(C[8]), .A2(net72879), .B1(A[8]), .B2(net70175), .ZN(n10)
         );
  NAND2_X1 U193 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  AOI22_X1 U194 ( .A1(C[9]), .A2(net72880), .B1(A[9]), .B2(net70175), .ZN(n3)
         );
  AOI222_X1 U195 ( .A1(D[9]), .A2(net70129), .B1(E[9]), .B2(n193), .C1(B[9]), 
        .C2(net70149), .ZN(n4) );
  NAND2_X1 U196 ( .A1(n120), .A2(n121), .ZN(Y[16]) );
  AOI22_X1 U197 ( .A1(C[16]), .A2(net72880), .B1(A[16]), .B2(net70175), .ZN(
        n120) );
  AOI222_X1 U198 ( .A1(D[16]), .A2(net70129), .B1(E[16]), .B2(n191), .C1(B[16]), .C2(net84586), .ZN(n121) );
  NAND2_X1 U199 ( .A1(n118), .A2(n119), .ZN(Y[17]) );
  AOI222_X1 U200 ( .A1(D[17]), .A2(net70129), .B1(E[17]), .B2(n185), .C1(B[17]), .C2(net84586), .ZN(n119) );
  AOI22_X1 U201 ( .A1(C[17]), .A2(net72882), .B1(A[17]), .B2(net70175), .ZN(
        n118) );
  NAND2_X1 U202 ( .A1(n24), .A2(n25), .ZN(Y[5]) );
  AOI22_X1 U203 ( .A1(C[5]), .A2(net72878), .B1(A[5]), .B2(net70175), .ZN(n24)
         );
  NAND2_X1 U204 ( .A1(n14), .A2(n15), .ZN(Y[6]) );
  AOI22_X1 U205 ( .A1(C[6]), .A2(net72878), .B1(A[6]), .B2(net70175), .ZN(n14)
         );
  AOI222_X1 U206 ( .A1(D[6]), .A2(net70125), .B1(n143), .B2(E[6]), .C1(B[6]), 
        .C2(net70149), .ZN(n15) );
  NAND2_X1 U207 ( .A1(n124), .A2(n125), .ZN(Y[14]) );
  AOI22_X1 U208 ( .A1(C[14]), .A2(net72879), .B1(A[14]), .B2(net70175), .ZN(
        n124) );
  NAND2_X1 U209 ( .A1(n88), .A2(n89), .ZN(Y[30]) );
  AOI22_X1 U210 ( .A1(C[30]), .A2(net72882), .B1(A[30]), .B2(net70175), .ZN(
        n88) );
  NAND2_X1 U211 ( .A1(n126), .A2(n127), .ZN(Y[13]) );
  AOI222_X1 U212 ( .A1(D[13]), .A2(net70129), .B1(E[13]), .B2(n193), .C1(B[13]), .C2(net70151), .ZN(n127) );
  AOI22_X1 U213 ( .A1(C[13]), .A2(net72879), .B1(A[13]), .B2(net70175), .ZN(
        n126) );
  AOI22_X1 U214 ( .A1(C[2]), .A2(net72878), .B1(A[2]), .B2(net70175), .ZN(n90)
         );
  AOI22_X1 U215 ( .A1(C[3]), .A2(net72880), .B1(A[3]), .B2(net70175), .ZN(n68)
         );
  AOI22_X1 U216 ( .A1(net72878), .A2(C[4]), .B1(A[4]), .B2(net70175), .ZN(n46)
         );
  NAND2_X1 U217 ( .A1(n42), .A2(n43), .ZN(Y[51]) );
  AOI22_X1 U218 ( .A1(C[51]), .A2(net72879), .B1(A[51]), .B2(net70175), .ZN(
        n42) );
  AOI222_X1 U219 ( .A1(D[51]), .A2(net70123), .B1(E[51]), .B2(net78774), .C1(
        B[51]), .C2(net91117), .ZN(n43) );
  NAND2_X1 U220 ( .A1(n36), .A2(n37), .ZN(Y[54]) );
  AOI22_X1 U221 ( .A1(C[54]), .A2(net72882), .B1(A[54]), .B2(net70175), .ZN(
        n36) );
  AOI222_X1 U222 ( .A1(D[54]), .A2(net70123), .B1(E[54]), .B2(net78774), .C1(
        B[54]), .C2(net91117), .ZN(n37) );
  NAND2_X1 U223 ( .A1(n38), .A2(n39), .ZN(Y[53]) );
  AOI22_X1 U224 ( .A1(C[53]), .A2(net72880), .B1(A[53]), .B2(net70175), .ZN(
        n38) );
  AOI222_X1 U225 ( .A1(D[53]), .A2(net70123), .B1(E[53]), .B2(net78774), .C1(
        B[53]), .C2(net91117), .ZN(n39) );
  NAND2_X1 U226 ( .A1(n32), .A2(n33), .ZN(Y[56]) );
  AOI22_X1 U227 ( .A1(C[56]), .A2(n181), .B1(A[56]), .B2(net70175), .ZN(n32)
         );
  AOI222_X1 U228 ( .A1(D[56]), .A2(net70125), .B1(E[56]), .B2(net78774), .C1(
        B[56]), .C2(net70149), .ZN(n33) );
  NAND2_X1 U229 ( .A1(n30), .A2(n31), .ZN(Y[57]) );
  AOI22_X1 U230 ( .A1(C[57]), .A2(net72879), .B1(A[57]), .B2(net70175), .ZN(
        n30) );
  AOI222_X1 U231 ( .A1(D[57]), .A2(net70129), .B1(E[57]), .B2(net78774), .C1(
        B[57]), .C2(net88405), .ZN(n31) );
  NAND2_X1 U232 ( .A1(n28), .A2(n29), .ZN(Y[58]) );
  AOI22_X1 U233 ( .A1(C[58]), .A2(net72880), .B1(A[58]), .B2(net70175), .ZN(
        n28) );
  AOI222_X1 U234 ( .A1(D[58]), .A2(net70125), .B1(E[58]), .B2(net78774), .C1(
        B[58]), .C2(net70149), .ZN(n29) );
  NAND2_X1 U235 ( .A1(n26), .A2(n27), .ZN(Y[59]) );
  AOI22_X1 U236 ( .A1(C[59]), .A2(net72882), .B1(A[59]), .B2(net70175), .ZN(
        n26) );
  AOI222_X1 U237 ( .A1(D[59]), .A2(net70129), .B1(E[59]), .B2(net78774), .C1(
        B[59]), .C2(net88405), .ZN(n27) );
  NAND2_X1 U238 ( .A1(n50), .A2(n51), .ZN(Y[48]) );
  AOI22_X1 U239 ( .A1(C[48]), .A2(net72882), .B1(A[48]), .B2(net70175), .ZN(
        n50) );
  AOI222_X1 U240 ( .A1(D[48]), .A2(net70123), .B1(E[48]), .B2(net78774), .C1(
        B[48]), .C2(net70151), .ZN(n51) );
  NAND2_X1 U241 ( .A1(n48), .A2(n49), .ZN(Y[49]) );
  AOI22_X1 U242 ( .A1(C[49]), .A2(net72880), .B1(A[49]), .B2(net70175), .ZN(
        n48) );
  AOI222_X1 U243 ( .A1(D[49]), .A2(net70123), .B1(E[49]), .B2(net78774), .C1(
        B[49]), .C2(net91117), .ZN(n49) );
  NAND2_X1 U244 ( .A1(n44), .A2(n45), .ZN(Y[50]) );
  AOI22_X1 U245 ( .A1(C[50]), .A2(n181), .B1(A[50]), .B2(net70175), .ZN(n44)
         );
  AOI222_X1 U246 ( .A1(D[50]), .A2(net70123), .B1(E[50]), .B2(net78774), .C1(
        B[50]), .C2(net91117), .ZN(n45) );
  NAND2_X1 U247 ( .A1(n40), .A2(n41), .ZN(Y[52]) );
  AOI22_X1 U248 ( .A1(C[52]), .A2(net72880), .B1(A[52]), .B2(net70175), .ZN(
        n40) );
  AOI222_X1 U249 ( .A1(D[52]), .A2(net70123), .B1(E[52]), .B2(net78774), .C1(
        B[52]), .C2(net70151), .ZN(n41) );
  NAND2_X1 U250 ( .A1(n34), .A2(n35), .ZN(Y[55]) );
  AOI22_X1 U251 ( .A1(C[55]), .A2(n181), .B1(A[55]), .B2(net70175), .ZN(n34)
         );
  AOI222_X1 U252 ( .A1(D[55]), .A2(net70123), .B1(E[55]), .B2(net78774), .C1(
        B[55]), .C2(net70151), .ZN(n35) );
  NAND2_X1 U253 ( .A1(n22), .A2(n23), .ZN(Y[60]) );
  AOI22_X1 U254 ( .A1(C[60]), .A2(net72882), .B1(A[60]), .B2(net70175), .ZN(
        n22) );
  AOI222_X1 U255 ( .A1(D[60]), .A2(net70127), .B1(E[60]), .B2(net78774), .C1(
        B[60]), .C2(net70149), .ZN(n23) );
  NAND2_X1 U256 ( .A1(n20), .A2(n21), .ZN(Y[61]) );
  AOI22_X1 U257 ( .A1(C[61]), .A2(net72882), .B1(A[61]), .B2(net70175), .ZN(
        n20) );
  AOI222_X1 U258 ( .A1(D[61]), .A2(net70125), .B1(E[61]), .B2(net78774), .C1(
        B[61]), .C2(net88405), .ZN(n21) );
  NAND2_X1 U259 ( .A1(n18), .A2(n19), .ZN(Y[62]) );
  AOI22_X1 U260 ( .A1(C[62]), .A2(n181), .B1(A[62]), .B2(net70175), .ZN(n18)
         );
  AOI222_X1 U261 ( .A1(D[62]), .A2(net70129), .B1(E[62]), .B2(net78774), .C1(
        B[62]), .C2(net70149), .ZN(n19) );
  NAND2_X1 U262 ( .A1(n16), .A2(n17), .ZN(Y[63]) );
  AOI22_X1 U263 ( .A1(C[63]), .A2(net72882), .B1(A[63]), .B2(net70175), .ZN(
        n16) );
  AOI222_X1 U264 ( .A1(D[63]), .A2(net70123), .B1(E[63]), .B2(net78774), .C1(
        B[63]), .C2(net88405), .ZN(n17) );
  AOI22_X1 U265 ( .A1(C[28]), .A2(net72880), .B1(A[28]), .B2(net70175), .ZN(
        n94) );
  CLKBUF_X1 U266 ( .A(n8), .Z(net72878) );
  AOI22_X1 U267 ( .A1(C[27]), .A2(n181), .B1(A[27]), .B2(net70175), .ZN(n96)
         );
  AOI222_X1 U268 ( .A1(D[27]), .A2(net70119), .B1(E[27]), .B2(net70133), .C1(
        B[27]), .C2(net91117), .ZN(n97) );
  NAND2_X1 U269 ( .A1(n76), .A2(n77), .ZN(Y[36]) );
  AOI222_X1 U270 ( .A1(D[36]), .A2(net70121), .B1(E[36]), .B2(n191), .C1(B[36]), .C2(net70149), .ZN(n77) );
  AOI22_X1 U271 ( .A1(C[0]), .A2(net72879), .B1(A[0]), .B2(net70175), .ZN(n134) );
  AOI222_X1 U272 ( .A1(D[1]), .A2(net70125), .B1(E[1]), .B2(n185), .C1(B[1]), 
        .C2(net84586), .ZN(n113) );
  AOI222_X1 U273 ( .A1(D[0]), .A2(net70129), .B1(E[0]), .B2(n185), .C1(B[0]), 
        .C2(net70149), .ZN(n135) );
  AOI22_X1 U274 ( .A1(C[1]), .A2(net72880), .B1(A[1]), .B2(net70175), .ZN(n112) );
  AOI222_X1 U275 ( .A1(D[2]), .A2(net70119), .B1(net70137), .B2(E[2]), .C1(
        B[2]), .C2(net70151), .ZN(n91) );
  NAND2_X1 U276 ( .A1(n134), .A2(n135), .ZN(Y[0]) );
  NAND2_X1 U277 ( .A1(n112), .A2(n113), .ZN(Y[1]) );
  AOI22_X1 U278 ( .A1(C[23]), .A2(net72880), .B1(A[23]), .B2(net70175), .ZN(
        n104) );
  NAND2_X1 U279 ( .A1(n94), .A2(n95), .ZN(Y[28]) );
  NAND2_X1 U280 ( .A1(n86), .A2(n87), .ZN(Y[31]) );
  AOI22_X1 U281 ( .A1(C[34]), .A2(net72879), .B1(A[34]), .B2(net70175), .ZN(
        n80) );
  AOI22_X1 U282 ( .A1(C[35]), .A2(net72882), .B1(A[35]), .B2(net70175), .ZN(
        n78) );
  AOI22_X1 U283 ( .A1(C[33]), .A2(net72882), .B1(A[33]), .B2(net70175), .ZN(
        n82) );
  AOI22_X1 U284 ( .A1(C[32]), .A2(n181), .B1(A[32]), .B2(net70175), .ZN(n84)
         );
  NAND2_X1 U285 ( .A1(n110), .A2(n111), .ZN(Y[20]) );
  AOI22_X1 U286 ( .A1(C[20]), .A2(net72879), .B1(A[20]), .B2(net70175), .ZN(
        n110) );
  AOI222_X1 U287 ( .A1(D[24]), .A2(net70119), .B1(E[24]), .B2(net70133), .C1(
        B[24]), .C2(net70151), .ZN(n103) );
  AOI22_X1 U288 ( .A1(C[31]), .A2(net72882), .B1(A[31]), .B2(net70175), .ZN(
        n86) );
  AOI222_X1 U289 ( .A1(D[3]), .A2(net70127), .B1(n184), .B2(E[3]), .C1(B[3]), 
        .C2(n182), .ZN(n69) );
endmodule


module Booth_Encoder_15 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   net83782, net87822, n4, n5, n6, n7, n8, n9, n10, n11;

  AND3_X2 U3 ( .A1(net83782), .A2(n6), .A3(i[2]), .ZN(o[2]) );
  OAI22_X1 U4 ( .A1(n4), .A2(n5), .B1(i[2]), .B2(n6), .ZN(o[1]) );
  INV_X1 U5 ( .A(i[2]), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n7), .A2(n8), .ZN(n4) );
  NAND2_X1 U7 ( .A1(i[0]), .A2(i[1]), .ZN(n8) );
  OR2_X1 U8 ( .A1(i[0]), .A2(i[1]), .ZN(n7) );
  AOI21_X1 U9 ( .B1(net87822), .B2(n6), .A(i[2]), .ZN(o[0]) );
  NAND2_X1 U10 ( .A1(i[0]), .A2(i[1]), .ZN(n6) );
  OR2_X1 U11 ( .A1(i[0]), .A2(i[1]), .ZN(n9) );
  OR2_X1 U12 ( .A1(i[0]), .A2(i[1]), .ZN(n10) );
  NAND2_X1 U13 ( .A1(n9), .A2(n11), .ZN(net87822) );
  NAND2_X1 U14 ( .A1(n10), .A2(n8), .ZN(net83782) );
  NAND2_X1 U15 ( .A1(i[0]), .A2(i[1]), .ZN(n11) );
endmodule


module MUX_booth_N64_15 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n14, n19, n69, n91, net71113, net71107, net71131, net71129, net71127,
         net71133, net71143, net71141, net71139, net71155, net71151, net71149,
         net71161, net84042, net84040, net85007, net85229, net86459, net89101,
         net89100, net89698, net89956, net90207, net90236, net90297, net90563,
         net90582, net90716, net90902, net90854, net91896, net99153, net99466,
         net99641, net99605, net90852, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307;

  AND2_X2 U1 ( .A1(n139), .A2(net90852), .ZN(net99153) );
  NAND2_X1 U2 ( .A1(n235), .A2(n234), .ZN(Y[32]) );
  INV_X1 U3 ( .A(D[2]), .ZN(n171) );
  INV_X1 U4 ( .A(D[3]), .ZN(n172) );
  BUF_X2 U5 ( .A(net71107), .Z(net89956) );
  NAND2_X1 U6 ( .A1(n222), .A2(n221), .ZN(Y[26]) );
  INV_X1 U7 ( .A(n158), .ZN(net71129) );
  AND2_X2 U8 ( .A1(n154), .A2(n153), .ZN(n139) );
  CLKBUF_X1 U9 ( .A(net99466), .Z(net71127) );
  BUF_X1 U10 ( .A(net99466), .Z(net90716) );
  AND2_X1 U11 ( .A1(net90852), .A2(n139), .ZN(n141) );
  AND2_X2 U12 ( .A1(n150), .A2(n161), .ZN(net71107) );
  BUF_X1 U13 ( .A(sel[1]), .Z(n161) );
  INV_X1 U14 ( .A(n157), .ZN(n140) );
  AND2_X1 U15 ( .A1(D[11]), .A2(net71113), .ZN(n142) );
  AND2_X1 U16 ( .A1(n141), .A2(E[11]), .ZN(n143) );
  AND2_X1 U17 ( .A1(B[11]), .A2(net71139), .ZN(n144) );
  NOR3_X1 U18 ( .A1(n142), .A2(n143), .A3(n144), .ZN(n189) );
  BUF_X1 U19 ( .A(net90236), .Z(net71113) );
  AND2_X1 U20 ( .A1(D[6]), .A2(net89956), .ZN(n145) );
  AND2_X1 U21 ( .A1(n141), .A2(E[6]), .ZN(n146) );
  AND2_X1 U22 ( .A1(B[6]), .A2(net99605), .ZN(n147) );
  NOR3_X1 U23 ( .A1(n145), .A2(n146), .A3(n147), .ZN(n165) );
  INV_X1 U24 ( .A(n158), .ZN(n148) );
  AND2_X1 U25 ( .A1(n160), .A2(n156), .ZN(n149) );
  CLKBUF_X1 U26 ( .A(net90207), .Z(net71155) );
  CLKBUF_X3 U27 ( .A(net85007), .Z(net71161) );
  NAND2_X1 U28 ( .A1(n155), .A2(sel[1]), .ZN(n154) );
  NOR2_X1 U29 ( .A1(sel[2]), .A2(sel[1]), .ZN(n156) );
  INV_X1 U30 ( .A(sel[1]), .ZN(n151) );
  NAND2_X1 U31 ( .A1(n150), .A2(n161), .ZN(net90852) );
  NOR3_X1 U32 ( .A1(n140), .A2(n161), .A3(n160), .ZN(net85007) );
  NAND2_X1 U33 ( .A1(net90852), .A2(n139), .ZN(n158) );
  NOR2_X1 U34 ( .A1(sel[0]), .A2(sel[2]), .ZN(n155) );
  INV_X1 U35 ( .A(sel[0]), .ZN(n152) );
  BUF_X2 U36 ( .A(net89101), .Z(n163) );
  INV_X1 U37 ( .A(n154), .ZN(net90207) );
  INV_X2 U38 ( .A(n159), .ZN(net89100) );
  INV_X1 U39 ( .A(net90207), .ZN(n159) );
  INV_X1 U40 ( .A(n152), .ZN(n160) );
  INV_X1 U41 ( .A(sel[2]), .ZN(n157) );
  NOR2_X1 U42 ( .A1(n152), .A2(sel[2]), .ZN(n150) );
  AND2_X1 U43 ( .A1(n154), .A2(n153), .ZN(n162) );
  CLKBUF_X1 U44 ( .A(net71139), .Z(n164) );
  NAND2_X1 U45 ( .A1(n157), .A2(n151), .ZN(n153) );
  NAND2_X1 U46 ( .A1(n14), .A2(n165), .ZN(Y[6]) );
  CLKBUF_X1 U47 ( .A(n149), .Z(net99605) );
  AOI222_X1 U48 ( .A1(D[62]), .A2(net91896), .B1(E[62]), .B2(net71127), .C1(
        B[62]), .C2(net99605), .ZN(n19) );
  AND2_X1 U49 ( .A1(net71107), .A2(D[5]), .ZN(net86459) );
  NOR2_X1 U50 ( .A1(net71107), .A2(net99641), .ZN(net85229) );
  AND2_X1 U51 ( .A1(n162), .A2(net90852), .ZN(net71133) );
  NAND2_X1 U52 ( .A1(n139), .A2(E[7]), .ZN(net99641) );
  BUF_X1 U53 ( .A(n149), .Z(net71141) );
  BUF_X2 U54 ( .A(net90297), .Z(net71143) );
  CLKBUF_X1 U55 ( .A(net71139), .Z(net90563) );
  INV_X1 U56 ( .A(net84040), .ZN(net84042) );
  INV_X1 U57 ( .A(net90854), .ZN(net99466) );
  INV_X1 U58 ( .A(net99153), .ZN(net90854) );
  AND2_X1 U59 ( .A1(D[12]), .A2(net90236), .ZN(n166) );
  AND2_X1 U60 ( .A1(E[12]), .A2(net99153), .ZN(n167) );
  AND2_X1 U61 ( .A1(B[12]), .A2(n149), .ZN(n168) );
  NOR3_X1 U62 ( .A1(n166), .A2(n167), .A3(n168), .ZN(n191) );
  BUF_X1 U63 ( .A(net71107), .Z(net90236) );
  BUF_X2 U64 ( .A(n149), .Z(net71139) );
  BUF_X2 U65 ( .A(net90236), .Z(net91896) );
  CLKBUF_X1 U66 ( .A(net99466), .Z(net89698) );
  NAND2_X1 U67 ( .A1(n149), .A2(B[3]), .ZN(n174) );
  NAND2_X1 U68 ( .A1(n149), .A2(B[2]), .ZN(n173) );
  OAI21_X1 U69 ( .B1(n172), .B2(net90902), .A(n174), .ZN(n170) );
  AOI21_X1 U70 ( .B1(net99153), .B2(E[3]), .A(n170), .ZN(n69) );
  OAI21_X1 U71 ( .B1(n171), .B2(net90902), .A(n173), .ZN(n169) );
  AOI21_X1 U72 ( .B1(net71127), .B2(E[2]), .A(n169), .ZN(n91) );
  BUF_X2 U73 ( .A(net71143), .Z(net90582) );
  INV_X1 U74 ( .A(net71107), .ZN(net90902) );
  CLKBUF_X1 U75 ( .A(net90716), .Z(net71131) );
  NAND2_X1 U76 ( .A1(n224), .A2(n223), .ZN(Y[27]) );
  CLKBUF_X1 U77 ( .A(n149), .Z(net90297) );
  NAND2_X1 U78 ( .A1(n307), .A2(n306), .ZN(Y[9]) );
  BUF_X1 U79 ( .A(net90207), .Z(net89101) );
  NAND2_X1 U80 ( .A1(n188), .A2(n187), .ZN(Y[10]) );
  BUF_X1 U81 ( .A(net90207), .Z(net71149) );
  BUF_X1 U82 ( .A(net90207), .Z(net71151) );
  AND2_X1 U83 ( .A1(net71107), .A2(D[4]), .ZN(n175) );
  AND2_X1 U84 ( .A1(net71133), .A2(E[4]), .ZN(n176) );
  AND2_X1 U85 ( .A1(B[4]), .A2(n149), .ZN(n177) );
  NOR3_X1 U86 ( .A1(n176), .A2(n175), .A3(n177), .ZN(n271) );
  AND2_X1 U87 ( .A1(net71133), .A2(E[5]), .ZN(n178) );
  AND2_X1 U88 ( .A1(B[5]), .A2(n149), .ZN(n179) );
  NOR3_X1 U89 ( .A1(n178), .A2(net86459), .A3(n179), .ZN(n293) );
  AND2_X1 U90 ( .A1(D[20]), .A2(net89956), .ZN(n180) );
  AND2_X1 U91 ( .A1(E[20]), .A2(net99466), .ZN(n181) );
  AND2_X1 U92 ( .A1(B[20]), .A2(net90563), .ZN(n182) );
  NOR3_X1 U93 ( .A1(n180), .A2(n181), .A3(n182), .ZN(n209) );
  AND2_X1 U94 ( .A1(net71107), .A2(D[7]), .ZN(n183) );
  AND2_X1 U95 ( .A1(B[7]), .A2(n149), .ZN(n184) );
  NOR3_X1 U96 ( .A1(net85229), .A2(n183), .A3(n184), .ZN(n302) );
  INV_X1 U97 ( .A(net71139), .ZN(net84040) );
  NAND2_X1 U98 ( .A1(n302), .A2(n303), .ZN(Y[7]) );
  NAND2_X1 U99 ( .A1(n293), .A2(n294), .ZN(Y[5]) );
  NAND2_X1 U100 ( .A1(n271), .A2(n272), .ZN(Y[4]) );
  NAND2_X1 U101 ( .A1(n243), .A2(n242), .ZN(Y[36]) );
  AOI22_X1 U102 ( .A1(C[36]), .A2(net71151), .B1(A[36]), .B2(net71161), .ZN(
        n243) );
  AOI222_X1 U103 ( .A1(D[36]), .A2(net91896), .B1(E[36]), .B2(net71129), .C1(
        B[36]), .C2(net90582), .ZN(n242) );
  AOI22_X1 U104 ( .A1(C[37]), .A2(net89100), .B1(A[37]), .B2(net71161), .ZN(
        n245) );
  AOI22_X1 U105 ( .A1(C[7]), .A2(net71149), .B1(A[7]), .B2(net71161), .ZN(n303) );
  NAND2_X1 U106 ( .A1(n305), .A2(n304), .ZN(Y[8]) );
  AOI22_X1 U107 ( .A1(C[8]), .A2(net71155), .B1(A[8]), .B2(net71161), .ZN(n305) );
  AOI222_X1 U108 ( .A1(D[8]), .A2(net90236), .B1(net99153), .B2(E[8]), .C1(
        B[8]), .C2(n149), .ZN(n304) );
  NAND2_X1 U109 ( .A1(n249), .A2(n248), .ZN(Y[39]) );
  AOI22_X1 U110 ( .A1(C[39]), .A2(net71151), .B1(A[39]), .B2(net71161), .ZN(
        n249) );
  AOI222_X1 U111 ( .A1(D[39]), .A2(net91896), .B1(E[39]), .B2(net90716), .C1(
        B[39]), .C2(net84042), .ZN(n248) );
  NAND2_X1 U112 ( .A1(n241), .A2(n240), .ZN(Y[35]) );
  AOI22_X1 U113 ( .A1(C[35]), .A2(n163), .B1(A[35]), .B2(net71161), .ZN(n241)
         );
  AOI222_X1 U114 ( .A1(D[35]), .A2(net91896), .B1(E[35]), .B2(net71131), .C1(
        B[35]), .C2(net71143), .ZN(n240) );
  AOI22_X1 U115 ( .A1(C[4]), .A2(net90207), .B1(A[4]), .B2(net71161), .ZN(n272) );
  NAND2_X1 U116 ( .A1(n256), .A2(n255), .ZN(Y[42]) );
  AOI22_X1 U117 ( .A1(C[42]), .A2(net89101), .B1(A[42]), .B2(net71161), .ZN(
        n256) );
  AOI222_X1 U118 ( .A1(D[42]), .A2(net91896), .B1(E[42]), .B2(net71129), .C1(
        B[42]), .C2(net84042), .ZN(n255) );
  NAND2_X1 U119 ( .A1(n262), .A2(n261), .ZN(Y[45]) );
  AOI22_X1 U120 ( .A1(C[45]), .A2(n163), .B1(A[45]), .B2(net71161), .ZN(n262)
         );
  AOI222_X1 U121 ( .A1(D[45]), .A2(net91896), .B1(E[45]), .B2(net71127), .C1(
        B[45]), .C2(net84042), .ZN(n261) );
  NAND2_X1 U122 ( .A1(n264), .A2(n263), .ZN(Y[46]) );
  AOI22_X1 U123 ( .A1(C[46]), .A2(net71151), .B1(A[46]), .B2(net71161), .ZN(
        n264) );
  AOI222_X1 U124 ( .A1(D[46]), .A2(net91896), .B1(E[46]), .B2(net71127), .C1(
        B[46]), .C2(net90563), .ZN(n263) );
  AOI222_X1 U125 ( .A1(D[32]), .A2(net91896), .B1(E[32]), .B2(net71127), .C1(
        B[32]), .C2(net84042), .ZN(n234) );
  AOI22_X1 U126 ( .A1(C[32]), .A2(net89100), .B1(A[32]), .B2(net71161), .ZN(
        n235) );
  NAND2_X1 U127 ( .A1(n239), .A2(n238), .ZN(Y[34]) );
  AOI222_X1 U128 ( .A1(D[34]), .A2(net91896), .B1(E[34]), .B2(net71127), .C1(
        B[34]), .C2(net90563), .ZN(n238) );
  AOI22_X1 U129 ( .A1(C[34]), .A2(n163), .B1(A[34]), .B2(net71161), .ZN(n239)
         );
  NAND2_X1 U130 ( .A1(n237), .A2(n236), .ZN(Y[33]) );
  AOI22_X1 U131 ( .A1(C[33]), .A2(n163), .B1(A[33]), .B2(net71161), .ZN(n237)
         );
  NAND2_X1 U132 ( .A1(n220), .A2(n219), .ZN(Y[25]) );
  AOI22_X1 U133 ( .A1(C[25]), .A2(n163), .B1(A[25]), .B2(net71161), .ZN(n220)
         );
  AOI22_X1 U134 ( .A1(C[26]), .A2(net71151), .B1(A[26]), .B2(net71161), .ZN(
        n222) );
  NAND2_X1 U135 ( .A1(n191), .A2(n192), .ZN(Y[12]) );
  AOI22_X1 U136 ( .A1(C[12]), .A2(net90207), .B1(A[12]), .B2(net71161), .ZN(
        n192) );
  NAND2_X1 U137 ( .A1(n200), .A2(n199), .ZN(Y[16]) );
  AOI222_X1 U138 ( .A1(D[16]), .A2(net71113), .B1(E[16]), .B2(net71129), .C1(
        B[16]), .C2(net71143), .ZN(n199) );
  AOI22_X1 U139 ( .A1(C[16]), .A2(n163), .B1(A[16]), .B2(net71161), .ZN(n200)
         );
  NAND2_X1 U140 ( .A1(n252), .A2(n251), .ZN(Y[40]) );
  AOI22_X1 U141 ( .A1(C[40]), .A2(net89100), .B1(A[40]), .B2(net71161), .ZN(
        n252) );
  AOI222_X1 U142 ( .A1(D[40]), .A2(net91896), .B1(E[40]), .B2(net71129), .C1(
        B[40]), .C2(net84042), .ZN(n251) );
  NAND2_X1 U143 ( .A1(n247), .A2(n246), .ZN(Y[38]) );
  AOI22_X1 U144 ( .A1(C[38]), .A2(n163), .B1(A[38]), .B2(net71161), .ZN(n247)
         );
  AOI222_X1 U145 ( .A1(D[38]), .A2(net91896), .B1(E[38]), .B2(net90716), .C1(
        B[38]), .C2(net71143), .ZN(n246) );
  NAND2_X1 U146 ( .A1(n260), .A2(n259), .ZN(Y[44]) );
  AOI22_X1 U147 ( .A1(C[44]), .A2(net89100), .B1(A[44]), .B2(net71161), .ZN(
        n260) );
  AOI222_X1 U148 ( .A1(D[44]), .A2(net91896), .B1(E[44]), .B2(n148), .C1(B[44]), .C2(net84042), .ZN(n259) );
  NAND2_X1 U149 ( .A1(n254), .A2(n253), .ZN(Y[41]) );
  AOI22_X1 U150 ( .A1(C[41]), .A2(net71151), .B1(A[41]), .B2(net71161), .ZN(
        n254) );
  AOI222_X1 U151 ( .A1(D[41]), .A2(net91896), .B1(E[41]), .B2(net90716), .C1(
        B[41]), .C2(net71143), .ZN(n253) );
  NAND2_X1 U152 ( .A1(n258), .A2(n257), .ZN(Y[43]) );
  AOI22_X1 U153 ( .A1(C[43]), .A2(net89100), .B1(A[43]), .B2(net71161), .ZN(
        n258) );
  AOI222_X1 U154 ( .A1(D[43]), .A2(net91896), .B1(E[43]), .B2(net71127), .C1(
        B[43]), .C2(net84042), .ZN(n257) );
  NAND2_X1 U155 ( .A1(n266), .A2(n265), .ZN(Y[47]) );
  AOI22_X1 U156 ( .A1(C[47]), .A2(net89101), .B1(A[47]), .B2(net71161), .ZN(
        n266) );
  AOI222_X1 U157 ( .A1(D[47]), .A2(net91896), .B1(E[47]), .B2(net71127), .C1(
        B[47]), .C2(net84042), .ZN(n265) );
  AOI22_X1 U158 ( .A1(C[9]), .A2(net71155), .B1(A[9]), .B2(net71161), .ZN(n307) );
  AOI222_X1 U159 ( .A1(D[9]), .A2(net89956), .B1(E[9]), .B2(n141), .C1(B[9]), 
        .C2(net90297), .ZN(n306) );
  NAND2_X1 U160 ( .A1(n202), .A2(n201), .ZN(Y[17]) );
  AOI222_X1 U161 ( .A1(D[17]), .A2(net89956), .B1(E[17]), .B2(net99466), .C1(
        B[17]), .C2(net90563), .ZN(n201) );
  AOI22_X1 U162 ( .A1(C[17]), .A2(net71151), .B1(A[17]), .B2(net71161), .ZN(
        n202) );
  NAND2_X1 U163 ( .A1(n212), .A2(n211), .ZN(Y[21]) );
  AOI222_X1 U164 ( .A1(D[21]), .A2(net89956), .B1(E[21]), .B2(net89698), .C1(
        B[21]), .C2(net84042), .ZN(n211) );
  AOI22_X1 U165 ( .A1(C[21]), .A2(net89100), .B1(A[21]), .B2(net71161), .ZN(
        n212) );
  AOI22_X1 U166 ( .A1(C[10]), .A2(net89100), .B1(A[10]), .B2(net71161), .ZN(
        n188) );
  AOI222_X1 U167 ( .A1(D[10]), .A2(net89956), .B1(E[10]), .B2(net99466), .C1(
        B[10]), .C2(net71139), .ZN(n187) );
  NAND2_X1 U168 ( .A1(n190), .A2(n189), .ZN(Y[11]) );
  AOI22_X1 U169 ( .A1(C[11]), .A2(net89100), .B1(A[11]), .B2(net71161), .ZN(
        n190) );
  NAND2_X1 U170 ( .A1(n204), .A2(n203), .ZN(Y[18]) );
  AOI222_X1 U171 ( .A1(D[18]), .A2(net89956), .B1(E[18]), .B2(net89698), .C1(
        B[18]), .C2(net90582), .ZN(n203) );
  AOI22_X1 U172 ( .A1(C[18]), .A2(n163), .B1(A[18]), .B2(net71161), .ZN(n204)
         );
  NAND2_X1 U173 ( .A1(n198), .A2(n197), .ZN(Y[15]) );
  AOI222_X1 U174 ( .A1(D[15]), .A2(net89956), .B1(E[15]), .B2(net99466), .C1(
        B[15]), .C2(net71139), .ZN(n197) );
  AOI22_X1 U175 ( .A1(C[15]), .A2(net71151), .B1(A[15]), .B2(net71161), .ZN(
        n198) );
  NAND2_X1 U176 ( .A1(n206), .A2(n205), .ZN(Y[19]) );
  AOI222_X1 U177 ( .A1(D[19]), .A2(net89956), .B1(E[19]), .B2(net71129), .C1(
        B[19]), .C2(net71143), .ZN(n205) );
  AOI22_X1 U178 ( .A1(C[19]), .A2(net89100), .B1(A[19]), .B2(net71161), .ZN(
        n206) );
  AOI22_X1 U179 ( .A1(C[5]), .A2(net71149), .B1(A[5]), .B2(net71161), .ZN(n294) );
  NAND2_X1 U180 ( .A1(n231), .A2(n230), .ZN(Y[30]) );
  AOI22_X1 U181 ( .A1(C[30]), .A2(net89100), .B1(A[30]), .B2(net71161), .ZN(
        n231) );
  NAND2_X1 U182 ( .A1(n209), .A2(n210), .ZN(Y[20]) );
  AOI22_X1 U183 ( .A1(C[20]), .A2(n163), .B1(A[20]), .B2(net71161), .ZN(n210)
         );
  NAND2_X1 U184 ( .A1(n218), .A2(n217), .ZN(Y[24]) );
  AOI22_X1 U185 ( .A1(C[24]), .A2(net89100), .B1(A[24]), .B2(net71161), .ZN(
        n218) );
  AOI222_X1 U186 ( .A1(D[24]), .A2(net91896), .B1(E[24]), .B2(net89698), .C1(
        B[24]), .C2(net90582), .ZN(n217) );
  NAND2_X1 U187 ( .A1(n214), .A2(n213), .ZN(Y[22]) );
  AOI22_X1 U188 ( .A1(C[22]), .A2(net71151), .B1(A[22]), .B2(net71161), .ZN(
        n214) );
  AOI222_X1 U189 ( .A1(D[22]), .A2(net71113), .B1(E[22]), .B2(net90716), .C1(
        B[22]), .C2(net84042), .ZN(n213) );
  NAND2_X1 U190 ( .A1(n194), .A2(n193), .ZN(Y[13]) );
  AOI22_X1 U191 ( .A1(C[13]), .A2(net71151), .B1(A[13]), .B2(net71161), .ZN(
        n194) );
  AOI222_X1 U192 ( .A1(D[13]), .A2(net89956), .B1(n141), .B2(E[13]), .C1(B[13]), .C2(net71141), .ZN(n193) );
  NAND2_X1 U193 ( .A1(n196), .A2(n195), .ZN(Y[14]) );
  AOI22_X1 U194 ( .A1(C[14]), .A2(net89101), .B1(A[14]), .B2(net71161), .ZN(
        n196) );
  AOI222_X1 U195 ( .A1(D[14]), .A2(net71113), .B1(n148), .B2(E[14]), .C1(B[14]), .C2(net71139), .ZN(n195) );
  AOI22_X1 U196 ( .A1(C[6]), .A2(net89101), .B1(A[6]), .B2(net71161), .ZN(n14)
         );
  NAND2_X1 U197 ( .A1(n228), .A2(n227), .ZN(Y[29]) );
  AOI22_X1 U198 ( .A1(C[29]), .A2(n163), .B1(A[29]), .B2(net71161), .ZN(n228)
         );
  NAND2_X1 U199 ( .A1(n226), .A2(n225), .ZN(Y[28]) );
  AOI22_X1 U200 ( .A1(C[28]), .A2(net89100), .B1(A[28]), .B2(net71161), .ZN(
        n226) );
  AOI222_X1 U201 ( .A1(D[28]), .A2(net91896), .B1(E[28]), .B2(net71129), .C1(
        B[28]), .C2(n164), .ZN(n225) );
  NAND2_X1 U202 ( .A1(n216), .A2(n215), .ZN(Y[23]) );
  AOI222_X1 U203 ( .A1(D[23]), .A2(net89956), .B1(E[23]), .B2(net89698), .C1(
        B[23]), .C2(net90582), .ZN(n215) );
  AOI22_X1 U204 ( .A1(C[23]), .A2(n163), .B1(A[23]), .B2(net71161), .ZN(n216)
         );
  AOI222_X1 U205 ( .A1(D[27]), .A2(net91896), .B1(E[27]), .B2(net90716), .C1(
        B[27]), .C2(n164), .ZN(n223) );
  AOI22_X1 U206 ( .A1(C[27]), .A2(n163), .B1(A[27]), .B2(net71161), .ZN(n224)
         );
  NAND2_X1 U207 ( .A1(n233), .A2(n232), .ZN(Y[31]) );
  AOI22_X1 U208 ( .A1(C[31]), .A2(n163), .B1(A[31]), .B2(net71161), .ZN(n233)
         );
  AOI222_X1 U209 ( .A1(D[31]), .A2(net91896), .B1(E[31]), .B2(net71131), .C1(
        B[31]), .C2(net90582), .ZN(n232) );
  NAND2_X1 U210 ( .A1(n282), .A2(n281), .ZN(Y[54]) );
  AOI222_X1 U211 ( .A1(D[54]), .A2(net91896), .B1(E[54]), .B2(net71127), .C1(
        B[54]), .C2(net71143), .ZN(n281) );
  NAND2_X1 U212 ( .A1(n284), .A2(n283), .ZN(Y[55]) );
  AOI222_X1 U213 ( .A1(D[55]), .A2(net91896), .B1(E[55]), .B2(net90716), .C1(
        B[55]), .C2(net71141), .ZN(n283) );
  NAND2_X1 U214 ( .A1(n286), .A2(n285), .ZN(Y[56]) );
  AOI222_X1 U215 ( .A1(D[56]), .A2(net91896), .B1(E[56]), .B2(net71127), .C1(
        B[56]), .C2(n164), .ZN(n285) );
  NAND2_X1 U216 ( .A1(n288), .A2(n287), .ZN(Y[57]) );
  AOI222_X1 U217 ( .A1(D[57]), .A2(net91896), .B1(E[57]), .B2(n148), .C1(B[57]), .C2(net71143), .ZN(n287) );
  NAND2_X1 U218 ( .A1(n290), .A2(n289), .ZN(Y[58]) );
  AOI222_X1 U219 ( .A1(D[58]), .A2(net91896), .B1(E[58]), .B2(net71129), .C1(
        B[58]), .C2(net71143), .ZN(n289) );
  NAND2_X1 U220 ( .A1(n268), .A2(n267), .ZN(Y[48]) );
  AOI22_X1 U221 ( .A1(C[48]), .A2(net89100), .B1(A[48]), .B2(net71161), .ZN(
        n268) );
  AOI222_X1 U222 ( .A1(D[48]), .A2(net91896), .B1(E[48]), .B2(net71129), .C1(
        B[48]), .C2(net71139), .ZN(n267) );
  NAND2_X1 U223 ( .A1(n270), .A2(n269), .ZN(Y[49]) );
  AOI22_X1 U224 ( .A1(C[49]), .A2(n163), .B1(A[49]), .B2(net71161), .ZN(n270)
         );
  AOI222_X1 U225 ( .A1(D[49]), .A2(net91896), .B1(E[49]), .B2(net90716), .C1(
        B[49]), .C2(net71143), .ZN(n269) );
  NAND2_X1 U226 ( .A1(n274), .A2(n273), .ZN(Y[50]) );
  AOI22_X1 U227 ( .A1(C[50]), .A2(net89100), .B1(A[50]), .B2(net71161), .ZN(
        n274) );
  AOI222_X1 U228 ( .A1(D[50]), .A2(net91896), .B1(E[50]), .B2(net71127), .C1(
        B[50]), .C2(net71139), .ZN(n273) );
  NAND2_X1 U229 ( .A1(n276), .A2(n275), .ZN(Y[51]) );
  AOI22_X1 U230 ( .A1(C[51]), .A2(net71151), .B1(A[51]), .B2(net71161), .ZN(
        n276) );
  AOI222_X1 U231 ( .A1(D[51]), .A2(net91896), .B1(E[51]), .B2(net71129), .C1(
        B[51]), .C2(net71139), .ZN(n275) );
  NAND2_X1 U232 ( .A1(n278), .A2(n277), .ZN(Y[52]) );
  AOI22_X1 U233 ( .A1(C[52]), .A2(net71155), .B1(A[52]), .B2(net71161), .ZN(
        n278) );
  AOI222_X1 U234 ( .A1(D[52]), .A2(net91896), .B1(E[52]), .B2(net71127), .C1(
        B[52]), .C2(n164), .ZN(n277) );
  NAND2_X1 U235 ( .A1(n280), .A2(n279), .ZN(Y[53]) );
  AOI22_X1 U236 ( .A1(C[53]), .A2(n163), .B1(A[53]), .B2(net71161), .ZN(n280)
         );
  AOI222_X1 U237 ( .A1(D[53]), .A2(net91896), .B1(E[53]), .B2(net71129), .C1(
        B[53]), .C2(n164), .ZN(n279) );
  NAND2_X1 U238 ( .A1(n292), .A2(n291), .ZN(Y[59]) );
  AOI222_X1 U239 ( .A1(D[59]), .A2(net91896), .B1(E[59]), .B2(net90716), .C1(
        B[59]), .C2(net71141), .ZN(n291) );
  NAND2_X1 U240 ( .A1(n296), .A2(n295), .ZN(Y[60]) );
  AOI22_X1 U241 ( .A1(C[60]), .A2(net89100), .B1(A[60]), .B2(net71161), .ZN(
        n296) );
  AOI222_X1 U242 ( .A1(D[60]), .A2(net91896), .B1(E[60]), .B2(net71127), .C1(
        B[60]), .C2(net71143), .ZN(n295) );
  NAND2_X1 U243 ( .A1(n298), .A2(n297), .ZN(Y[61]) );
  AOI22_X1 U244 ( .A1(C[61]), .A2(n163), .B1(A[61]), .B2(net71161), .ZN(n298)
         );
  AOI222_X1 U245 ( .A1(D[61]), .A2(net91896), .B1(E[61]), .B2(n148), .C1(B[61]), .C2(n164), .ZN(n297) );
  NAND2_X1 U246 ( .A1(n299), .A2(n19), .ZN(Y[62]) );
  NAND2_X1 U247 ( .A1(n301), .A2(n300), .ZN(Y[63]) );
  AOI222_X1 U248 ( .A1(D[63]), .A2(net91896), .B1(E[63]), .B2(net71129), .C1(
        B[63]), .C2(net71141), .ZN(n300) );
  NAND2_X1 U249 ( .A1(n186), .A2(n185), .ZN(Y[0]) );
  AOI22_X1 U250 ( .A1(C[0]), .A2(net71155), .B1(A[0]), .B2(net71161), .ZN(n186) );
  AOI222_X1 U251 ( .A1(D[0]), .A2(net91896), .B1(E[0]), .B2(net71127), .C1(
        B[0]), .C2(n164), .ZN(n185) );
  NAND2_X1 U252 ( .A1(n208), .A2(n207), .ZN(Y[1]) );
  AOI22_X1 U253 ( .A1(C[1]), .A2(net89101), .B1(A[1]), .B2(net71161), .ZN(n208) );
  AOI222_X1 U254 ( .A1(D[1]), .A2(net91896), .B1(E[1]), .B2(net90716), .C1(
        B[1]), .C2(net90297), .ZN(n207) );
  NAND2_X1 U255 ( .A1(n245), .A2(n244), .ZN(Y[37]) );
  AOI222_X1 U256 ( .A1(D[37]), .A2(net91896), .B1(E[37]), .B2(net71127), .C1(
        B[37]), .C2(net90563), .ZN(n244) );
  AOI222_X1 U257 ( .A1(D[29]), .A2(net91896), .B1(E[29]), .B2(net71127), .C1(
        B[29]), .C2(net90582), .ZN(n227) );
  AOI22_X1 U258 ( .A1(C[2]), .A2(net90207), .B1(A[2]), .B2(net71161), .ZN(n229) );
  NAND2_X1 U259 ( .A1(n250), .A2(n69), .ZN(Y[3]) );
  NAND2_X1 U260 ( .A1(n229), .A2(n91), .ZN(Y[2]) );
  AOI22_X1 U261 ( .A1(C[3]), .A2(net71149), .B1(A[3]), .B2(net71161), .ZN(n250) );
  AOI222_X1 U262 ( .A1(D[30]), .A2(net91896), .B1(E[30]), .B2(net71131), .C1(
        B[30]), .C2(net84042), .ZN(n230) );
  AOI222_X1 U263 ( .A1(D[25]), .A2(net91896), .B1(E[25]), .B2(net71129), .C1(
        B[25]), .C2(n164), .ZN(n219) );
  AOI22_X1 U264 ( .A1(C[63]), .A2(net71151), .B1(A[63]), .B2(net71161), .ZN(
        n301) );
  AOI22_X1 U265 ( .A1(C[62]), .A2(net89100), .B1(A[62]), .B2(net71161), .ZN(
        n299) );
  AOI22_X1 U266 ( .A1(C[59]), .A2(net71151), .B1(A[59]), .B2(net71161), .ZN(
        n292) );
  AOI22_X1 U267 ( .A1(C[58]), .A2(n163), .B1(A[58]), .B2(net71161), .ZN(n290)
         );
  AOI22_X1 U268 ( .A1(C[57]), .A2(n163), .B1(A[57]), .B2(net71161), .ZN(n288)
         );
  AOI22_X1 U269 ( .A1(C[56]), .A2(net89100), .B1(A[56]), .B2(net71161), .ZN(
        n286) );
  AOI22_X1 U270 ( .A1(C[55]), .A2(net71151), .B1(A[55]), .B2(net71161), .ZN(
        n284) );
  AOI22_X1 U271 ( .A1(C[54]), .A2(net89100), .B1(A[54]), .B2(net71161), .ZN(
        n282) );
  AOI222_X1 U272 ( .A1(D[26]), .A2(net91896), .B1(E[26]), .B2(net71127), .C1(
        B[26]), .C2(net84042), .ZN(n221) );
  AOI222_X1 U273 ( .A1(D[33]), .A2(net91896), .B1(E[33]), .B2(n148), .C1(B[33]), .C2(net90563), .ZN(n236) );
endmodule


module G_0 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n2) );
endmodule


module PG_0 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n2;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n2) );
  INV_X1 U3 ( .A(n2), .ZN(Gx) );
endmodule


module PG_944 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_943 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_942 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_941 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_940 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_939 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_938 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_937 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_936 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_935 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_934 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_933 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_932 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_931 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_930 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_929 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_928 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_927 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_926 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_925 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_924 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_923 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_922 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_921 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_920 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_919 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_918 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_917 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_916 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_915 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_254 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_914 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_913 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_912 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_911 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_910 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_909 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_908 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_907 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_906 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_905 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_904 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_903 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_902 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_901 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_900 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_253 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_899 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_898 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_897 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_896 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_895 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_894 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_893 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_252 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
endmodule


module G_251 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_892 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_891 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_890 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_889 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_888 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_887 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_250 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n3, n5;

  AND2_X1 U1 ( .A1(P_IK), .A2(G_K_1), .ZN(n3) );
  NOR2_X1 U2 ( .A1(n3), .A2(G_IK), .ZN(n5) );
  INV_X1 U3 ( .A(n5), .ZN(Gx) );
endmodule


module G_249 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_248 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_247 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
endmodule


module PG_886 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_885 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_884 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_883 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_246 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_245 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_244 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_243 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_242 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_241 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_240 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_239 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module carry_generator_N64_NPB4_0 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   n16, n17, \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n3, n4, n6, n7, n8, n9,
         n10, n11, n12, n14, n15;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(A[6]), .B(B[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U77 ( .A(B[59]), .B(A[59]), .Z(\PG_Network[0][0][59] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U81 ( .A(B[55]), .B(A[55]), .Z(\PG_Network[0][0][55] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U85 ( .A(B[51]), .B(A[51]), .Z(\PG_Network[0][0][51] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U88 ( .A(B[49]), .B(A[49]), .Z(\PG_Network[0][0][49] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U90 ( .A(B[47]), .B(A[47]), .Z(\PG_Network[0][0][47] ) );
  XOR2_X1 U91 ( .A(B[46]), .B(A[46]), .Z(\PG_Network[0][0][46] ) );
  XOR2_X1 U92 ( .A(B[45]), .B(A[45]), .Z(\PG_Network[0][0][45] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U94 ( .A(B[43]), .B(A[43]), .Z(\PG_Network[0][0][43] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(A[3]), .B(B[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U99 ( .A(B[39]), .B(A[39]), .Z(\PG_Network[0][0][39] ) );
  XOR2_X1 U100 ( .A(B[38]), .B(A[38]), .Z(\PG_Network[0][0][38] ) );
  XOR2_X1 U101 ( .A(B[37]), .B(A[37]), .Z(\PG_Network[0][0][37] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U103 ( .A(B[35]), .B(A[35]), .Z(\PG_Network[0][0][35] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U107 ( .A(A[31]), .B(B[31]), .Z(\PG_Network[0][0][31] ) );
  XOR2_X1 U108 ( .A(B[30]), .B(A[30]), .Z(\PG_Network[0][0][30] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U110 ( .A(B[29]), .B(A[29]), .Z(\PG_Network[0][0][29] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U112 ( .A(B[27]), .B(A[27]), .Z(\PG_Network[0][0][27] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U114 ( .A(B[25]), .B(A[25]), .Z(\PG_Network[0][0][25] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U116 ( .A(B[23]), .B(A[23]), .Z(\PG_Network[0][0][23] ) );
  XOR2_X1 U117 ( .A(A[22]), .B(B[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U121 ( .A(B[19]), .B(A[19]), .Z(\PG_Network[0][0][19] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(A[10]), .B(B[10]), .Z(\PG_Network[0][0][10] ) );
  G_0 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n14), .Gx(\PG_Network[1][1][1] ) );
  PG_0 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), 
        .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_944 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_943 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_942 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_941 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_940 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_939 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_938 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_937 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_936 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_935 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_934 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_933 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_932 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_931 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_930 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_929 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_928 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_927 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_926 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_925 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_924 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_923 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_922 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_921 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_920 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_919 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_918 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_917 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_916 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_915 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_254 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(n17) );
  PG_914 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_913 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_912 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_911 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_910 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_909 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_908 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_907 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_906 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_905 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_904 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_903 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_902 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_901 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_900 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_253 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(n17), .Gx(Co[1]) );
  PG_899 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_898 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_897 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_896 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_895 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_894 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_893 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_252 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), .G_K_1(Co[1]), .Gx(n16) );
  G_251 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_892 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_891 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_890 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][47] ), .Px(
        \PG_Network[4][0][47] ) );
  PG_889 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][43] ), .Px(
        \PG_Network[4][0][43] ) );
  PG_888 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][63] ), .Px(
        \PG_Network[4][0][63] ) );
  PG_887 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][59] ), .Px(
        \PG_Network[4][0][59] ) );
  G_250 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), .G_K_1(n6), .Gx(Co[7]) );
  G_249 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), .G_K_1(n6), .Gx(Co[6]) );
  G_248 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), .G_K_1(Co[3]), .Gx(Co[5]) );
  G_247 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), .G_K_1(n16), .Gx(Co[4]) );
  PG_886 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][63] ), .Px(
        \PG_Network[5][0][63] ) );
  PG_885 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][59] ), .Px(
        \PG_Network[5][0][59] ) );
  PG_884 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][55] ), .Px(
        \PG_Network[5][0][55] ) );
  PG_883 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][51] ), .Px(
        \PG_Network[5][0][51] ) );
  G_246 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), .G_K_1(n12), .Gx(Co[15]) );
  G_245 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), .G_K_1(n12), .Gx(Co[14]) );
  G_244 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), .G_K_1(n12), .Gx(Co[13]) );
  G_243 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), .G_K_1(n12), .Gx(Co[12]) );
  G_242 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), .G_K_1(n11), .Gx(Co[11]) );
  G_241 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), .G_K_1(n11), .Gx(Co[10]) );
  G_240 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), .G_K_1(Co[7]), .Gx(Co[9]) );
  G_239 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), .G_K_1(Co[7]), .Gx(Co[8]) );
  BUF_X2 U1 ( .A(n17), .Z(Co[0]) );
  BUF_X2 U2 ( .A(n16), .Z(Co[3]) );
  CLKBUF_X1 U3 ( .A(Co[3]), .Z(n6) );
  NAND2_X1 U4 ( .A1(A[15]), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(B[15]), .A2(n7), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n9), .A2(n10), .ZN(\PG_Network[0][0][15] ) );
  INV_X1 U7 ( .A(A[15]), .ZN(n7) );
  INV_X1 U8 ( .A(B[15]), .ZN(n8) );
  CLKBUF_X1 U9 ( .A(Co[7]), .Z(n11) );
  CLKBUF_X1 U10 ( .A(n11), .Z(n12) );
  AND2_X1 U11 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U12 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U13 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U14 ( .A1(B[7]), .A2(A[7]), .ZN(\PG_Network[0][1][7] ) );
  AND2_X1 U15 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U16 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U17 ( .A1(A[37]), .A2(B[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U18 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U19 ( .A1(A[35]), .A2(B[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U20 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U21 ( .A1(A[39]), .A2(B[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U22 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AND2_X1 U23 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U24 ( .A1(A[19]), .A2(B[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U25 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U26 ( .A1(B[11]), .A2(A[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U27 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U28 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U29 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AND2_X1 U30 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U31 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U32 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U33 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U34 ( .A1(A[25]), .A2(B[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U35 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U36 ( .A1(A[43]), .A2(B[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U37 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U38 ( .A1(A[41]), .A2(B[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U39 ( .A1(A[46]), .A2(B[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U40 ( .A1(A[47]), .A2(B[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U41 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U42 ( .A1(A[45]), .A2(B[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U43 ( .A1(B[5]), .A2(A[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U44 ( .A1(A[29]), .A2(B[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U45 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U46 ( .A1(A[15]), .A2(B[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U47 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U48 ( .A1(B[21]), .A2(A[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U49 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U50 ( .A1(A[51]), .A2(B[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U51 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U52 ( .A1(A[49]), .A2(B[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U53 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U54 ( .A1(A[59]), .A2(B[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U55 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
  AND2_X1 U56 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U57 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U58 ( .A1(A[53]), .A2(B[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U59 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U60 ( .A1(A[55]), .A2(B[55]), .ZN(\PG_Network[0][1][55] ) );
  INV_X1 U61 ( .A(n3), .ZN(n14) );
  AND2_X1 U62 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U63 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U64 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U65 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U66 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AOI21_X1 U67 ( .B1(A[0]), .B2(B[0]), .A(n15), .ZN(n3) );
  INV_X1 U125 ( .A(n4), .ZN(n15) );
  OAI21_X1 U131 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n4) );
  AND2_X1 U132 ( .A1(B[27]), .A2(A[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U133 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U134 ( .A1(B[23]), .A2(A[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U135 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U136 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  AND2_X1 U137 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U138 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U139 ( .A1(A[31]), .A2(B[31]), .ZN(\PG_Network[0][1][31] ) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n2) );
endmodule


module FA_1919 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1918 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1917 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1919 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1918 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1917 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1916 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1915 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1914 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1913 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_479 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1916 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1915 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1914 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1913 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_0 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n6, n7, n8, n9, n13;

  INV_X1 U1 ( .A(n7), .ZN(Y[2]) );
  AOI22_X1 U2 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n7) );
  INV_X1 U3 ( .A(n9), .ZN(Y[0]) );
  AOI22_X1 U4 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n9) );
  INV_X1 U5 ( .A(n8), .ZN(Y[1]) );
  AOI22_X1 U6 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n8) );
  INV_X1 U7 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n6) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_0 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_479 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_0 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1912 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n8, n9, n11, n12;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n11), .Z(n4) );
  NAND2_X1 U2 ( .A1(A), .A2(n6), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n5), .A2(B), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n7), .A2(n8), .ZN(n11) );
  INV_X1 U6 ( .A(A), .ZN(n5) );
  INV_X1 U7 ( .A(B), .ZN(n6) );
  CLKBUF_X1 U8 ( .A(A), .Z(n9) );
  AOI22_X1 U9 ( .A1(B), .A2(n9), .B1(n11), .B2(Ci), .ZN(n12) );
  INV_X1 U10 ( .A(n12), .ZN(Co) );
endmodule


module FA_1911 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6, n7, n8;

  XOR2_X1 U3 ( .A(n5), .B(n8), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  NAND2_X1 U1 ( .A1(n7), .A2(n6), .ZN(Co) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n5) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n8), .ZN(n7) );
endmodule


module FA_1910 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_1909 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(n4), .ZN(n7) );
endmodule


module RCA_N4_478 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1912 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1911 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1910 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1909 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1908 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1907 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1906 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1905 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_477 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1908 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1907 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1906 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1905 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_239 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U6 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U7 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U8 ( .A(sel), .ZN(n13) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n13), .ZN(n17) );
endmodule


module carry_select_block_NPB4_239 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_478 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_477 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_239 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1904 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  CLKBUF_X1 U1 ( .A(n8), .Z(n4) );
  CLKBUF_X1 U2 ( .A(A), .Z(n5) );
  CLKBUF_X1 U5 ( .A(B), .Z(n6) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n6), .A2(n5), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_1903 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_1902 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_1901 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_476 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1904 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1903 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1902 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1901 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1900 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1899 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1898 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1897 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_475 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1900 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1899 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1898 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1897 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_238 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U2 ( .A(n16), .ZN(Y[1]) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n5) );
  INV_X1 U4 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U5 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U6 ( .A(sel), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n14), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n14), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(n5), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
endmodule


module carry_select_block_NPB4_238 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_476 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_475 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_238 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1896 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  CLKBUF_X1 U1 ( .A(n8), .Z(n4) );
  CLKBUF_X1 U2 ( .A(A), .Z(n5) );
  CLKBUF_X1 U5 ( .A(B), .Z(n6) );
  AOI22_X1 U6 ( .A1(n6), .A2(n5), .B1(n8), .B2(Ci), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_1895 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1894 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1893 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n7), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_474 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1896 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1895 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1894 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1893 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1892 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1891 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n7), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  CLKBUF_X1 U1 ( .A(A), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n5), .A2(n4), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1890 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1889 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_473 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1892 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1891 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1890 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1889 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_237 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19;

  CLKBUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U4 ( .A(sel), .ZN(n10) );
  INV_X1 U5 ( .A(sel), .ZN(n11) );
  INV_X1 U6 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U7 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(n5), .A2(A[2]), .B1(n10), .B2(B[2]), .ZN(n18) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[1]), .B1(n11), .B2(B[1]), .ZN(n17) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[3]), .B1(n10), .B2(B[3]), .ZN(n19) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n11), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_237 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_474 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_473 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_237 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1888 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1887 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1886 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1885 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_472 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1888 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1887 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1886 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1885 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1884 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1883 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1882 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1881 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_471 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1884 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1883 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1882 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1881 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_236 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n11), .ZN(n5) );
  BUF_X1 U4 ( .A(sel), .Z(n11) );
  INV_X1 U5 ( .A(sel), .ZN(n10) );
  INV_X1 U6 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U7 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(n11), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(n11), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U10 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n10), .ZN(n17) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n10), .ZN(n16) );
endmodule


module carry_select_block_NPB4_236 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_472 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_471 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_236 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1880 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  CLKBUF_X1 U2 ( .A(A), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(n5), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1879 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1878 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1877 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_470 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1880 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1879 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1878 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1877 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1876 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1875 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1874 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1873 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_469 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1876 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1875 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1874 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1873 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_235 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U4 ( .A(sel), .ZN(n5) );
  INV_X1 U5 ( .A(n17), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[2]), .B1(B[2]), .B2(n5), .ZN(n17) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n5), .ZN(n16) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n14), .ZN(n15) );
  INV_X1 U9 ( .A(sel), .ZN(n14) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n5), .ZN(n18) );
endmodule


module carry_select_block_NPB4_235 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_470 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_469 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_235 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1872 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1871 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1870 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n7), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  NAND2_X1 U1 ( .A1(n5), .A2(n6), .ZN(Co) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U5 ( .A1(n7), .A2(Ci), .ZN(n6) );
endmodule


module FA_1869 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_468 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1872 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1871 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1870 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1869 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1868 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1867 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1866 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1865 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_467 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1868 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1867 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1866 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1865 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_234 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18;

  CLKBUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(sel), .ZN(n10) );
  INV_X1 U3 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U5 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U6 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n10), .ZN(n17) );
  AOI22_X1 U8 ( .A1(n5), .A2(A[3]), .B1(B[3]), .B2(n10), .ZN(n18) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n10), .ZN(n16) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n10), .ZN(n15) );
endmodule


module carry_select_block_NPB4_234 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_468 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_467 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_234 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1864 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(A), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n5) );
  AOI22_X1 U5 ( .A1(B), .A2(n4), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_1863 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1862 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1861 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_466 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1864 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1863 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1862 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1861 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1860 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1859 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1858 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1857 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_465 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1860 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1859 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1858 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1857 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_233 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(sel), .Z(n5) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(n10), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U9 ( .A1(n5), .A2(A[3]), .B1(B[3]), .B2(n15), .ZN(n19) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(A[0]), .A2(sel), .B1(n15), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_233 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_466 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_465 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_233 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1856 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  NAND2_X1 U1 ( .A1(A), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(n9) );
  INV_X1 U5 ( .A(A), .ZN(n4) );
  INV_X1 U6 ( .A(B), .ZN(n5) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
  INV_X1 U8 ( .A(n10), .ZN(Co) );
endmodule


module FA_1855 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1854 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1853 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_464 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1856 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1855 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1854 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1853 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1852 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1851 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1850 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1849 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_463 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1852 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1851 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1850 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1849 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_232 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n15), .ZN(Y[0]) );
  CLKBUF_X1 U2 ( .A(n14), .Z(n5) );
  INV_X1 U3 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n17) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(sel), .B1(n5), .B2(B[3]), .ZN(n18) );
  INV_X1 U10 ( .A(sel), .ZN(n14) );
endmodule


module carry_select_block_NPB4_232 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_464 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_463 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_232 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1848 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1847 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1846 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1845 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_462 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1848 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1847 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1846 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1845 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1844 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1843 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1842 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1841 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_461 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1844 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1843 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1842 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1841 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_231 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y[3]) );
  INV_X2 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U6 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n13), .ZN(n17) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(sel), .ZN(n13) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_231 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_462 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_461 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_231 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1840 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1839 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1838 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1837 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_460 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1840 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1839 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1838 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1837 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1836 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1835 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1834 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1833 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_459 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1836 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1835 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1834 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1833 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_230 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X2 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(sel), .ZN(n13) );
  INV_X1 U3 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U4 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U5 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U7 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_230 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_460 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_459 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_230 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1832 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1831 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1830 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1829 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_458 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1832 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1831 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1830 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1829 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1828 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1827 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1826 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1825 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_457 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1828 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1827 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1826 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1825 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_229 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_229 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_458 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_457 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_229 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1824 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1823 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1822 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1821 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_456 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1824 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1823 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1822 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1821 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1820 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1819 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1818 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1817 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_455 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1820 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1819 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1818 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1817 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_228 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_228 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_456 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_455 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_228 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1816 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1815 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1814 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1813 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_454 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1816 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1815 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1814 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1813 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1812 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1811 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1810 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1809 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_453 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1812 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1811 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1810 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1809 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_227 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_227 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_454 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_453 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_227 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1808 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1807 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1806 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1805 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_452 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1808 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1807 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1806 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1805 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1804 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1803 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1802 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1801 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_451 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1804 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1803 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1802 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1801 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_226 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_226 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_452 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_451 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_226 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1800 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1799 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1798 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1797 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_450 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1800 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1799 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1798 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1797 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1796 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1795 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1794 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1793 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_449 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1796 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1795 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1794 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1793 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_225 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_225 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_450 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_449 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_225 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_0 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_0 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_239 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_238 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_237 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_236 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_235 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_234 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_233 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_232 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_231 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_230 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), .S(S[43:40]) );
  carry_select_block_NPB4_229 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), .S(S[47:44]) );
  carry_select_block_NPB4_228 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), .S(S[51:48]) );
  carry_select_block_NPB4_227 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), .S(S[55:52]) );
  carry_select_block_NPB4_226 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), .S(S[59:56]) );
  carry_select_block_NPB4_225 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), .S(S[63:60]) );
endmodule


module P4_ADDER_N64_0 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_0 CGEN ( .A({A[63:25], n9, A[23:21], n2, A[19:17], 
        n17, A[15:13], n20, A[11:9], n22, A[7:5], n27, A[3:0]}), .B({B[63:33], 
        n21, B[31:21], n18, B[19:13], n5, B[11:9], n6, B[7:5], n13, B[3:0]}), 
        .Cin(Cin), .Co(CoutCgen) );
  sum_generator_N64_NPB4_0 SGEN ( .A({A[63:32], n12, A[30:16], n14, A[14:8], 
        n1, n3, A[5:4], n25, A[2:0]}), .B({B[63:32], n24, B[30:24], n11, 
        B[22:20], n15, B[18:16], n19, n4, B[13:11], n16, B[9:8], n8, n7, 
        B[5:4], n26, n10, B[1:0]}), .Ci({CoutCgen, Cin}), .S(S), .Co(Cout) );
  BUF_X1 U1 ( .A(B[14]), .Z(n4) );
  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(A[20]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(A[6]), .Z(n3) );
  CLKBUF_X1 U5 ( .A(B[12]), .Z(n5) );
  CLKBUF_X1 U6 ( .A(B[8]), .Z(n6) );
  BUF_X1 U7 ( .A(B[6]), .Z(n7) );
  CLKBUF_X1 U8 ( .A(B[7]), .Z(n8) );
  CLKBUF_X1 U9 ( .A(A[24]), .Z(n9) );
  CLKBUF_X1 U10 ( .A(B[2]), .Z(n10) );
  CLKBUF_X1 U11 ( .A(B[23]), .Z(n11) );
  CLKBUF_X1 U12 ( .A(A[31]), .Z(n12) );
  CLKBUF_X1 U13 ( .A(B[4]), .Z(n13) );
  CLKBUF_X1 U14 ( .A(A[15]), .Z(n14) );
  BUF_X1 U15 ( .A(B[19]), .Z(n15) );
  BUF_X1 U16 ( .A(B[10]), .Z(n16) );
  CLKBUF_X1 U17 ( .A(A[16]), .Z(n17) );
  CLKBUF_X1 U18 ( .A(B[20]), .Z(n18) );
  CLKBUF_X1 U19 ( .A(B[15]), .Z(n19) );
  CLKBUF_X1 U20 ( .A(A[12]), .Z(n20) );
  CLKBUF_X1 U21 ( .A(B[32]), .Z(n21) );
  CLKBUF_X1 U22 ( .A(A[8]), .Z(n22) );
  INV_X1 U23 ( .A(B[31]), .ZN(n23) );
  INV_X1 U24 ( .A(n23), .ZN(n24) );
  CLKBUF_X1 U25 ( .A(A[3]), .Z(n25) );
  CLKBUF_X1 U26 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U27 ( .A(A[4]), .Z(n27) );
endmodule


module Booth_Encoder_14 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_14 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305;

  NOR3_X1 U1 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U2 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  NOR4_X1 U3 ( .A1(n151), .A2(n145), .A3(n154), .A4(n167), .ZN(n139) );
  AOI222_X1 U4 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n158), .ZN(n298) );
  NAND2_X1 U5 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  NAND2_X1 U6 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI222_X1 U7 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n154), .ZN(n188) );
  AOI222_X1 U8 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n154), .ZN(n186) );
  BUF_X2 U9 ( .A(n165), .Z(n167) );
  BUF_X2 U10 ( .A(n152), .Z(n154) );
  CLKBUF_X1 U11 ( .A(n165), .Z(n169) );
  CLKBUF_X1 U12 ( .A(n165), .Z(n168) );
  CLKBUF_X1 U13 ( .A(n152), .Z(n156) );
  CLKBUF_X1 U14 ( .A(n152), .Z(n155) );
  CLKBUF_X1 U15 ( .A(n303), .Z(n166) );
  CLKBUF_X1 U16 ( .A(n302), .Z(n153) );
  BUF_X1 U17 ( .A(n139), .Z(n159) );
  BUF_X1 U18 ( .A(n139), .Z(n163) );
  BUF_X1 U19 ( .A(n139), .Z(n160) );
  BUF_X1 U20 ( .A(n139), .Z(n162) );
  BUF_X1 U21 ( .A(n139), .Z(n161) );
  BUF_X1 U22 ( .A(n153), .Z(n157) );
  BUF_X1 U23 ( .A(n153), .Z(n158) );
  BUF_X1 U24 ( .A(n166), .Z(n171) );
  BUF_X1 U25 ( .A(n166), .Z(n170) );
  CLKBUF_X1 U26 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U27 ( .A(n301), .Z(n148) );
  CLKBUF_X1 U28 ( .A(n301), .Z(n146) );
  CLKBUF_X1 U29 ( .A(n301), .Z(n147) );
  BUF_X1 U30 ( .A(n303), .Z(n165) );
  BUF_X1 U31 ( .A(n302), .Z(n152) );
  CLKBUF_X1 U32 ( .A(n301), .Z(n149) );
  CLKBUF_X1 U33 ( .A(n300), .Z(n142) );
  CLKBUF_X1 U34 ( .A(n300), .Z(n143) );
  CLKBUF_X1 U35 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U36 ( .A(n300), .Z(n141) );
  CLKBUF_X1 U37 ( .A(n300), .Z(n140) );
  INV_X1 U38 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U39 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n303) );
  AND3_X1 U40 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U41 ( .A(sel[2]), .ZN(n173) );
  NAND2_X1 U42 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  AOI22_X1 U43 ( .A1(C[32]), .A2(n149), .B1(A[32]), .B2(n143), .ZN(n225) );
  NAND2_X1 U44 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI22_X1 U45 ( .A1(C[39]), .A2(n148), .B1(A[39]), .B2(n142), .ZN(n239) );
  AOI222_X1 U46 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n156), .ZN(n238) );
  NAND2_X1 U47 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI22_X1 U48 ( .A1(C[45]), .A2(n148), .B1(A[45]), .B2(n142), .ZN(n253) );
  AOI222_X1 U49 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n157), .ZN(n252) );
  NAND2_X1 U50 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI22_X1 U51 ( .A1(C[46]), .A2(n147), .B1(A[46]), .B2(n141), .ZN(n255) );
  AOI222_X1 U52 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n157), .ZN(n254) );
  NAND2_X1 U53 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U54 ( .A1(C[6]), .A2(n146), .B1(A[6]), .B2(n140), .ZN(n295) );
  NAND2_X1 U55 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI22_X1 U56 ( .A1(C[35]), .A2(n149), .B1(A[35]), .B2(n143), .ZN(n231) );
  NAND2_X1 U57 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U58 ( .A1(C[7]), .A2(n146), .B1(A[7]), .B2(n140), .ZN(n297) );
  NAND2_X1 U59 ( .A1(n305), .A2(n304), .ZN(Y[9]) );
  AOI22_X1 U60 ( .A1(C[9]), .A2(n148), .B1(A[9]), .B2(n142), .ZN(n305) );
  NAND2_X1 U61 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  AOI22_X1 U62 ( .A1(C[40]), .A2(n148), .B1(A[40]), .B2(n142), .ZN(n243) );
  AOI222_X1 U63 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n156), .ZN(n242) );
  NAND2_X1 U64 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI22_X1 U65 ( .A1(C[37]), .A2(n148), .B1(A[37]), .B2(n142), .ZN(n235) );
  AOI222_X1 U66 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n156), .ZN(n234) );
  NAND2_X1 U67 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  AOI22_X1 U68 ( .A1(C[44]), .A2(n148), .B1(A[44]), .B2(n142), .ZN(n251) );
  AOI222_X1 U69 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n157), .ZN(n250) );
  NAND2_X1 U70 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI22_X1 U71 ( .A1(C[41]), .A2(n148), .B1(A[41]), .B2(n142), .ZN(n245) );
  AOI222_X1 U72 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n156), .ZN(n244) );
  NAND2_X1 U73 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI22_X1 U74 ( .A1(C[42]), .A2(n148), .B1(A[42]), .B2(n142), .ZN(n247) );
  AOI222_X1 U75 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n156), .ZN(n246) );
  NAND2_X1 U76 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI22_X1 U77 ( .A1(C[43]), .A2(n148), .B1(A[43]), .B2(n142), .ZN(n249) );
  AOI222_X1 U78 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n156), .ZN(n248) );
  NAND2_X1 U79 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U80 ( .A1(C[11]), .A2(n151), .B1(A[11]), .B2(n145), .ZN(n179) );
  AOI222_X1 U81 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n154), .ZN(n178) );
  NAND2_X1 U82 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U83 ( .A1(C[15]), .A2(n150), .B1(A[15]), .B2(n144), .ZN(n187) );
  NAND2_X1 U84 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI222_X1 U85 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n155), .ZN(n204) );
  AOI22_X1 U86 ( .A1(C[23]), .A2(n150), .B1(A[23]), .B2(n144), .ZN(n205) );
  NAND2_X1 U87 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  AOI22_X1 U88 ( .A1(C[16]), .A2(n150), .B1(A[16]), .B2(n144), .ZN(n189) );
  NAND2_X1 U89 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI22_X1 U90 ( .A1(C[38]), .A2(n148), .B1(A[38]), .B2(n142), .ZN(n237) );
  AOI222_X1 U91 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n156), .ZN(n236) );
  NAND2_X1 U92 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U93 ( .A1(C[10]), .A2(n151), .B1(A[10]), .B2(n145), .ZN(n177) );
  AOI222_X1 U94 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n154), .ZN(n176) );
  NAND2_X1 U95 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U96 ( .A1(C[14]), .A2(n150), .B1(A[14]), .B2(n144), .ZN(n185) );
  AOI222_X1 U97 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n154), .ZN(n184) );
  NAND2_X1 U98 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI222_X1 U99 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n154), .ZN(n192) );
  AOI22_X1 U100 ( .A1(C[18]), .A2(n150), .B1(A[18]), .B2(n144), .ZN(n193) );
  NAND2_X1 U101 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI222_X1 U102 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n155), .ZN(n202) );
  AOI22_X1 U103 ( .A1(C[22]), .A2(n150), .B1(A[22]), .B2(n144), .ZN(n203) );
  NAND2_X1 U104 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI222_X1 U105 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n156), .ZN(n228) );
  AOI22_X1 U106 ( .A1(C[34]), .A2(n149), .B1(A[34]), .B2(n143), .ZN(n229) );
  NAND2_X1 U107 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI22_X1 U108 ( .A1(C[26]), .A2(n149), .B1(A[26]), .B2(n143), .ZN(n211) );
  AOI222_X1 U109 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n155), .ZN(n210) );
  NAND2_X1 U110 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U111 ( .A1(C[30]), .A2(n149), .B1(A[30]), .B2(n143), .ZN(n221) );
  AOI222_X1 U112 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n155), .ZN(n220) );
  NAND2_X1 U113 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U114 ( .A1(C[13]), .A2(n151), .B1(A[13]), .B2(n145), .ZN(n183) );
  AOI222_X1 U115 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n154), .ZN(n182) );
  NAND2_X1 U116 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI222_X1 U117 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n154), .ZN(n190) );
  AOI22_X1 U118 ( .A1(C[17]), .A2(n150), .B1(A[17]), .B2(n144), .ZN(n191) );
  NAND2_X1 U119 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI222_X1 U120 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n155), .ZN(n200) );
  AOI22_X1 U121 ( .A1(C[21]), .A2(n150), .B1(A[21]), .B2(n144), .ZN(n201) );
  NAND2_X1 U122 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI222_X1 U123 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n155), .ZN(n208) );
  AOI22_X1 U124 ( .A1(C[25]), .A2(n149), .B1(A[25]), .B2(n143), .ZN(n209) );
  NAND2_X1 U125 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI222_X1 U126 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n155), .ZN(n216) );
  AOI22_X1 U127 ( .A1(C[29]), .A2(n149), .B1(A[29]), .B2(n143), .ZN(n217) );
  NAND2_X1 U128 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  AOI22_X1 U129 ( .A1(C[20]), .A2(n150), .B1(A[20]), .B2(n144), .ZN(n199) );
  AOI222_X1 U130 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n155), .ZN(n198) );
  NAND2_X1 U131 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI22_X1 U132 ( .A1(C[8]), .A2(n146), .B1(A[8]), .B2(n140), .ZN(n299) );
  AOI222_X1 U133 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n154), .ZN(n194) );
  AOI22_X1 U134 ( .A1(C[19]), .A2(n150), .B1(A[19]), .B2(n144), .ZN(n195) );
  NAND2_X1 U135 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  AOI22_X1 U136 ( .A1(C[28]), .A2(n149), .B1(A[28]), .B2(n143), .ZN(n215) );
  NAND2_X1 U137 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI22_X1 U138 ( .A1(C[27]), .A2(n149), .B1(A[27]), .B2(n143), .ZN(n213) );
  NAND2_X1 U139 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI22_X1 U140 ( .A1(C[31]), .A2(n149), .B1(A[31]), .B2(n143), .ZN(n223) );
  AOI222_X1 U141 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n156), .ZN(n232) );
  AOI22_X1 U142 ( .A1(C[36]), .A2(n148), .B1(A[36]), .B2(n142), .ZN(n233) );
  NAND2_X1 U143 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  AOI22_X1 U144 ( .A1(C[24]), .A2(n150), .B1(A[24]), .B2(n144), .ZN(n207) );
  AOI222_X1 U145 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n155), .ZN(n206) );
  NAND2_X1 U146 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  AOI22_X1 U147 ( .A1(C[12]), .A2(n151), .B1(A[12]), .B2(n145), .ZN(n181) );
  AOI222_X1 U148 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n154), .ZN(n180) );
  NAND2_X1 U149 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI22_X1 U150 ( .A1(C[33]), .A2(n149), .B1(A[33]), .B2(n143), .ZN(n227) );
  AOI222_X1 U151 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n156), .ZN(n226) );
  NAND2_X1 U152 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI22_X1 U153 ( .A1(C[47]), .A2(n147), .B1(A[47]), .B2(n141), .ZN(n257) );
  AOI222_X1 U154 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n157), .ZN(n256) );
  NAND2_X1 U155 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  AOI22_X1 U156 ( .A1(C[48]), .A2(n147), .B1(A[48]), .B2(n141), .ZN(n259) );
  AOI222_X1 U157 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n157), .ZN(n258) );
  NAND2_X1 U158 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  AOI22_X1 U159 ( .A1(C[52]), .A2(n147), .B1(A[52]), .B2(n141), .ZN(n269) );
  AOI222_X1 U160 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n157), .ZN(n268) );
  NAND2_X1 U161 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI22_X1 U162 ( .A1(C[49]), .A2(n147), .B1(A[49]), .B2(n141), .ZN(n261) );
  AOI222_X1 U163 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n157), .ZN(n260) );
  NAND2_X1 U164 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI22_X1 U165 ( .A1(C[50]), .A2(n147), .B1(A[50]), .B2(n141), .ZN(n265) );
  AOI222_X1 U166 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n157), .ZN(n264) );
  NAND2_X1 U167 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  AOI22_X1 U168 ( .A1(C[51]), .A2(n147), .B1(A[51]), .B2(n141), .ZN(n267) );
  AOI222_X1 U169 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n157), .ZN(n266) );
  NAND2_X1 U170 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  AOI22_X1 U171 ( .A1(C[56]), .A2(n147), .B1(A[56]), .B2(n141), .ZN(n277) );
  AOI222_X1 U172 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n158), .ZN(n276) );
  NAND2_X1 U173 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  AOI22_X1 U174 ( .A1(C[53]), .A2(n147), .B1(A[53]), .B2(n141), .ZN(n271) );
  AOI222_X1 U175 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n157), .ZN(n270) );
  NAND2_X1 U176 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI22_X1 U177 ( .A1(C[54]), .A2(n147), .B1(A[54]), .B2(n141), .ZN(n273) );
  AOI222_X1 U178 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n157), .ZN(n272) );
  NAND2_X1 U179 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI22_X1 U180 ( .A1(C[55]), .A2(n147), .B1(A[55]), .B2(n141), .ZN(n275) );
  AOI222_X1 U181 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n157), .ZN(n274) );
  NAND2_X1 U182 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  AOI22_X1 U183 ( .A1(C[57]), .A2(n146), .B1(A[57]), .B2(n140), .ZN(n279) );
  AOI222_X1 U184 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n158), .ZN(n278) );
  NAND2_X1 U185 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U186 ( .A1(C[60]), .A2(n146), .B1(A[60]), .B2(n140), .ZN(n287) );
  AOI222_X1 U187 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n158), .ZN(n286) );
  NAND2_X1 U188 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U189 ( .A1(C[61]), .A2(n146), .B1(A[61]), .B2(n140), .ZN(n289) );
  AOI222_X1 U190 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n158), .ZN(n288) );
  NAND2_X1 U191 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI22_X1 U192 ( .A1(C[58]), .A2(n146), .B1(A[58]), .B2(n140), .ZN(n281) );
  AOI222_X1 U193 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n158), .ZN(n280) );
  NAND2_X1 U194 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U195 ( .A1(C[62]), .A2(n146), .B1(A[62]), .B2(n140), .ZN(n291) );
  AOI222_X1 U196 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n158), .ZN(n290) );
  NAND2_X1 U197 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U198 ( .A1(C[59]), .A2(n146), .B1(A[59]), .B2(n140), .ZN(n283) );
  AOI222_X1 U199 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n158), .ZN(n282) );
  NAND2_X1 U200 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U201 ( .A1(C[63]), .A2(n146), .B1(A[63]), .B2(n140), .ZN(n293) );
  AOI222_X1 U202 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n158), .ZN(n292) );
  NAND2_X1 U203 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U204 ( .A1(C[0]), .A2(n146), .B1(A[0]), .B2(n140), .ZN(n175) );
  AOI222_X1 U205 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n154), .ZN(n174) );
  NAND2_X1 U206 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U207 ( .A1(C[1]), .A2(n150), .B1(A[1]), .B2(n144), .ZN(n197) );
  AOI222_X1 U208 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n154), .ZN(n196) );
  NAND2_X1 U209 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U210 ( .A1(C[2]), .A2(n149), .B1(A[2]), .B2(n143), .ZN(n219) );
  AOI222_X1 U211 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n155), .ZN(n218) );
  NAND2_X1 U212 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U213 ( .A1(C[3]), .A2(n148), .B1(A[3]), .B2(n142), .ZN(n241) );
  AOI222_X1 U214 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n156), .ZN(n240) );
  AOI222_X1 U215 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n155), .ZN(n222) );
  AOI22_X1 U216 ( .A1(C[4]), .A2(n147), .B1(A[4]), .B2(n141), .ZN(n263) );
  NAND2_X1 U217 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  NAND2_X1 U218 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U219 ( .A1(C[5]), .A2(n146), .B1(A[5]), .B2(n140), .ZN(n285) );
  AOI222_X1 U220 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n158), .ZN(n294) );
  AOI222_X1 U221 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n157), .ZN(n262) );
  AOI222_X1 U222 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n158), .ZN(n304) );
  AOI222_X1 U223 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n156), .ZN(n224) );
  AOI222_X1 U224 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n158), .ZN(n284) );
  AOI222_X1 U225 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n155), .ZN(n212) );
  AOI222_X1 U226 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n155), .ZN(n214) );
  AOI222_X1 U227 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n156), .ZN(n230) );
  AOI222_X1 U228 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n158), .ZN(n296) );
  CLKBUF_X1 U229 ( .A(n300), .Z(n145) );
  CLKBUF_X1 U230 ( .A(n301), .Z(n151) );
  CLKBUF_X1 U231 ( .A(n139), .Z(n164) );
endmodule


module G_238 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_882 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_881 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_880 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_879 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_878 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_877 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_876 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_875 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_874 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_873 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_872 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_871 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_870 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_869 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_868 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_867 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_866 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_865 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_864 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_863 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_862 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_861 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_860 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_859 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_858 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_857 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_856 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_855 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_854 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_853 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_852 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_237 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_851 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_850 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_849 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_848 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_847 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_846 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  OR2_X1 U2 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_845 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_844 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_843 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_842 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_841 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_840 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_839 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_838 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_837 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_236 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_836 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_835 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_834 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_833 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_832 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_831 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_830 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_235 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_234 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module PG_829 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_828 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_827 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_826 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_825 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_824 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_233 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_232 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_231 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module G_230 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_823 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_822 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_821 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_820 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_229 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_228 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_227 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_226 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_225 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_224 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module G_223 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_222 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module carry_generator_N64_NPB4_14 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   n17, \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n12, n13, n14, n15, n16;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U77 ( .A(B[59]), .B(A[59]), .Z(\PG_Network[0][0][59] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U81 ( .A(B[55]), .B(A[55]), .Z(\PG_Network[0][0][55] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U85 ( .A(B[51]), .B(A[51]), .Z(\PG_Network[0][0][51] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U88 ( .A(B[49]), .B(A[49]), .Z(\PG_Network[0][0][49] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U90 ( .A(B[47]), .B(A[47]), .Z(\PG_Network[0][0][47] ) );
  XOR2_X1 U91 ( .A(B[46]), .B(A[46]), .Z(\PG_Network[0][0][46] ) );
  XOR2_X1 U92 ( .A(B[45]), .B(A[45]), .Z(\PG_Network[0][0][45] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U94 ( .A(B[43]), .B(A[43]), .Z(\PG_Network[0][0][43] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U99 ( .A(B[39]), .B(A[39]), .Z(\PG_Network[0][0][39] ) );
  XOR2_X1 U100 ( .A(B[38]), .B(A[38]), .Z(\PG_Network[0][0][38] ) );
  XOR2_X1 U101 ( .A(B[37]), .B(A[37]), .Z(\PG_Network[0][0][37] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U103 ( .A(B[35]), .B(A[35]), .Z(\PG_Network[0][0][35] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U107 ( .A(B[31]), .B(A[31]), .Z(\PG_Network[0][0][31] ) );
  XOR2_X1 U108 ( .A(B[30]), .B(A[30]), .Z(\PG_Network[0][0][30] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U110 ( .A(B[29]), .B(A[29]), .Z(\PG_Network[0][0][29] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U112 ( .A(B[27]), .B(A[27]), .Z(\PG_Network[0][0][27] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U114 ( .A(B[25]), .B(A[25]), .Z(\PG_Network[0][0][25] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U116 ( .A(B[23]), .B(A[23]), .Z(\PG_Network[0][0][23] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U125 ( .A(B[15]), .B(A[15]), .Z(\PG_Network[0][0][15] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_238 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n13), .Gx(\PG_Network[1][1][1] ) );
  PG_882 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_881 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_880 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_879 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_878 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_877 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_876 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_875 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_874 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_873 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_872 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_871 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_870 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_869 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_868 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_867 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_866 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_865 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_864 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_863 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_862 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_861 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_860 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_859 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_858 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_857 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_856 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_855 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_854 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_853 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_852 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_237 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_851 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_850 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_849 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_848 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_847 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_846 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_845 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_844 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_843 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_842 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_841 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_840 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_839 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_838 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_837 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_236 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_836 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_835 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_834 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_833 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_832 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_831 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_830 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_235 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), .G_K_1(Co[1]), .Gx(n17) );
  G_234 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_829 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_828 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_827 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][47] ), .Px(
        \PG_Network[4][0][47] ) );
  PG_826 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][43] ), .Px(
        \PG_Network[4][0][43] ) );
  PG_825 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][63] ), .Px(
        \PG_Network[4][0][63] ) );
  PG_824 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][59] ), .Px(
        \PG_Network[4][0][59] ) );
  G_233 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), .G_K_1(n9), .Gx(Co[7]) );
  G_232 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), .G_K_1(n9), .Gx(Co[6]) );
  G_231 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), .G_K_1(Co[3]), .Gx(Co[5]) );
  G_230 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), .G_K_1(n17), .Gx(Co[4]) );
  PG_823 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][63] ), .Px(
        \PG_Network[5][0][63] ) );
  PG_822 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][59] ), .Px(
        \PG_Network[5][0][59] ) );
  PG_821 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][55] ), .Px(
        \PG_Network[5][0][55] ) );
  PG_820 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][51] ), .Px(
        \PG_Network[5][0][51] ) );
  G_229 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), .G_K_1(n12), .Gx(Co[15]) );
  G_228 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), .G_K_1(n12), .Gx(Co[14]) );
  G_227 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), .G_K_1(n12), .Gx(Co[13]) );
  G_226 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), .G_K_1(n12), .Gx(Co[12]) );
  G_225 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), .G_K_1(n12), .Gx(Co[11]) );
  G_224 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), .G_K_1(n12), .Gx(Co[10]) );
  G_223 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), .G_K_1(n12), .Gx(Co[9]) );
  G_222 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), .G_K_1(Co[7]), .Gx(Co[8]) );
  BUF_X2 U1 ( .A(Co[7]), .Z(n12) );
  NAND2_X1 U2 ( .A1(B[19]), .A2(n6), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n5), .A2(A[19]), .ZN(n8) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(\PG_Network[0][0][19] ) );
  INV_X1 U5 ( .A(B[19]), .ZN(n5) );
  INV_X1 U6 ( .A(A[19]), .ZN(n6) );
  INV_X1 U7 ( .A(A[34]), .ZN(n10) );
  CLKBUF_X1 U8 ( .A(Co[3]), .Z(n9) );
  BUF_X2 U9 ( .A(n17), .Z(Co[3]) );
  XNOR2_X1 U10 ( .A(B[34]), .B(n10), .ZN(\PG_Network[0][0][34] ) );
  AND2_X1 U11 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U12 ( .A1(A[35]), .A2(B[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U13 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U14 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U15 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U16 ( .A1(B[11]), .A2(A[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U17 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U18 ( .A1(A[41]), .A2(B[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U19 ( .A1(A[43]), .A2(B[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U20 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U21 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U22 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U23 ( .A1(B[7]), .A2(A[7]), .ZN(\PG_Network[0][1][7] ) );
  AND2_X1 U24 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AND2_X1 U25 ( .A1(B[23]), .A2(A[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U26 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U27 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U28 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U29 ( .A1(B[9]), .A2(A[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U30 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U31 ( .A1(A[19]), .A2(B[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U32 ( .A1(A[47]), .A2(B[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U33 ( .A1(A[46]), .A2(B[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U34 ( .A1(A[45]), .A2(B[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U35 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U36 ( .A1(B[13]), .A2(A[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U37 ( .A1(B[14]), .A2(A[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U38 ( .A1(B[15]), .A2(A[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U39 ( .A1(A[25]), .A2(B[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U40 ( .A1(A[37]), .A2(B[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U41 ( .A1(A[29]), .A2(B[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U42 ( .A1(B[20]), .A2(A[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U43 ( .A1(A[21]), .A2(B[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U44 ( .A1(A[49]), .A2(B[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U45 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U46 ( .A1(A[51]), .A2(B[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U47 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U48 ( .A1(A[59]), .A2(B[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U49 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U50 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
  AND2_X1 U51 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U52 ( .A1(A[53]), .A2(B[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U53 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U54 ( .A1(A[55]), .A2(B[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U55 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U56 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U57 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U58 ( .A(n16), .ZN(n13) );
  AND2_X1 U59 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U60 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U61 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U62 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U63 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AOI21_X1 U64 ( .B1(A[0]), .B2(B[0]), .A(n14), .ZN(n16) );
  INV_X1 U65 ( .A(n15), .ZN(n14) );
  OAI21_X1 U66 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n15) );
  AND2_X1 U67 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U104 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U121 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U131 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U132 ( .A1(B[31]), .A2(A[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U133 ( .A1(B[27]), .A2(A[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U134 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U135 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U136 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U137 ( .A1(B[12]), .A2(A[12]), .ZN(\PG_Network[0][1][12] ) );
  AND2_X1 U138 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
endmodule


module FA_1792 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1791 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1790 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1789 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_448 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1792 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1791 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1790 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1789 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1788 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1787 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1786 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1785 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_447 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1788 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1787 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1786 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1785 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_224 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U2 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U4 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U5 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U7 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_224 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_448 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_447 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_224 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1784 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1783 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1782 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1781 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_446 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1784 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1783 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1782 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1781 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1780 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1779 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n5), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1778 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1777 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_445 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1780 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1779 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1778 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1777 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_223 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U2 ( .A(sel), .ZN(n13) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_223 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2;
  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_446 UADDER1 ( .A(A), .B({B[3:2], n1, n2}), .Ci(1'b1), .S(S1) );
  RCA_N4_445 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_223 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
  CLKBUF_X1 U3 ( .A(B[1]), .Z(n1) );
  CLKBUF_X1 U4 ( .A(B[0]), .Z(n2) );
endmodule


module FA_1776 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1775 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1774 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1773 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_444 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1776 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1775 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1774 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1773 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1772 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1771 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1770 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1769 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_443 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1772 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1771 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1770 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1769 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_222 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n18), .ZN(Y[2]) );
  BUF_X1 U3 ( .A(sel), .Z(n10) );
  BUF_X1 U4 ( .A(n15), .Z(n5) );
  INV_X1 U5 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U7 ( .A(sel), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(n10), .B1(B[1]), .B2(n5), .ZN(n17) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
endmodule


module carry_select_block_NPB4_222 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_444 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_443 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_222 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1768 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n5), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1767 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1766 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1765 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n4), .B2(n6), .ZN(n7) );
endmodule


module RCA_N4_442 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1768 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1767 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1766 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1765 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1764 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1763 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1762 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1761 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_441 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1764 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1763 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1762 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1761 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_221 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  CLKBUF_X1 U1 ( .A(n10), .Z(n5) );
  BUF_X1 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U5 ( .A(sel), .ZN(n15) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U8 ( .A1(n10), .A2(A[1]), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n15), .ZN(n19) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X2 U11 ( .A(n16), .ZN(Y[0]) );
endmodule


module carry_select_block_NPB4_221 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_442 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_441 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_221 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1760 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n5) );
  AOI22_X1 U5 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_1759 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1758 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1757 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_440 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1760 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1759 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1758 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1757 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1756 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1755 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1754 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1753 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_439 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1756 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1755 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1754 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1753 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_220 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n18), .ZN(Y[2]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n5) );
  INV_X1 U3 ( .A(sel), .ZN(n10) );
  INV_X1 U4 ( .A(sel), .ZN(n11) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n10), .ZN(n17) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[0]), .B1(n11), .B2(B[0]), .ZN(n16) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n10), .ZN(n19) );
  INV_X2 U11 ( .A(n17), .ZN(Y[1]) );
endmodule


module carry_select_block_NPB4_220 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_440 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_439 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_220 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1752 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XNOR2_X1 U1 ( .A(B), .B(n5), .ZN(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1751 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1750 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1749 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_438 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1752 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1751 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1750 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1749 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1748 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1747 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1746 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1745 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_437 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1748 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1747 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1746 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1745 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_219 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U4 ( .A(sel), .ZN(n10) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U6 ( .A(sel), .ZN(n15) );
  INV_X1 U7 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U9 ( .A1(n5), .A2(A[1]), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n10), .B2(B[0]), .ZN(n16) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n15), .ZN(n19) );
endmodule


module carry_select_block_NPB4_219 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_438 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_437 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_219 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1744 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1743 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1742 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1741 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_436 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1744 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1743 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1742 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1741 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1740 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1739 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1738 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1737 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_435 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1740 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1739 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1738 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1737 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_218 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  CLKBUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U3 ( .A(sel), .ZN(n10) );
  INV_X1 U4 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n15), .ZN(n17) );
  INV_X1 U8 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(n5), .A2(A[3]), .B1(B[3]), .B2(n15), .ZN(n19) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n10), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_218 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_436 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_435 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_218 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1736 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1735 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1734 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1733 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_434 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1736 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1735 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1734 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1733 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1732 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1731 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1730 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1729 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_433 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1732 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1731 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1730 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1729 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_217 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  CLKBUF_X1 U1 ( .A(n15), .Z(n5) );
  INV_X1 U2 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[0]) );
  CLKBUF_X1 U4 ( .A(sel), .Z(n10) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[1]), .B1(n15), .B2(B[1]), .ZN(n17) );
  INV_X1 U9 ( .A(sel), .ZN(n15) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
  INV_X1 U11 ( .A(n19), .ZN(Y[3]) );
endmodule


module carry_select_block_NPB4_217 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_434 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_433 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_217 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1728 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1727 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1726 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1725 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_432 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1728 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1727 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1726 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1725 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1724 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1723 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1722 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1721 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_431 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1724 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1723 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1722 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1721 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_216 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U6 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U7 ( .A(sel), .ZN(n13) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n13), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_216 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_432 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_431 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_216 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1720 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(n4) );
  NAND2_X1 U2 ( .A1(n8), .A2(Ci), .ZN(n5) );
  AND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(n9) );
  XOR2_X1 U6 ( .A(A), .B(B), .Z(n6) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_1719 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1718 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1717 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_430 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1720 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1719 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1718 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1717 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1716 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1715 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1714 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1713 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_429 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1716 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1715 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1714 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1713 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_215 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n10), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n10) );
  INV_X1 U4 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_215 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_430 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_429 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_215 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1712 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1711 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1710 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1709 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_428 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1712 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1711 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1710 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1709 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1708 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1707 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1706 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1705 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_427 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1708 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1707 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1706 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1705 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_214 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(sel), .ZN(n5) );
  INV_X1 U3 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n16) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n17) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n5), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(n5), .B2(B[0]), .ZN(n14) );
endmodule


module carry_select_block_NPB4_214 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_428 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_427 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_214 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1704 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1703 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1702 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1701 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_426 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1704 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1703 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1702 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1701 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1700 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1699 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1698 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1697 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_425 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1700 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1699 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1698 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1697 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_213 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18;

  BUF_X1 U1 ( .A(n10), .Z(n5) );
  INV_X1 U2 ( .A(sel), .ZN(n10) );
  INV_X1 U3 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U4 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n18) );
  INV_X1 U5 ( .A(n17), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n17) );
  INV_X1 U7 ( .A(n16), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n5), .ZN(n16) );
  INV_X1 U9 ( .A(n15), .ZN(Y[0]) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n10), .ZN(n15) );
endmodule


module carry_select_block_NPB4_213 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_426 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_425 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_213 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1696 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1695 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1694 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1693 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_424 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1696 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1695 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1694 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1693 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1692 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1691 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1690 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1689 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_423 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1692 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1691 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1690 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1689 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_212 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_212 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_424 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_423 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_212 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1688 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1687 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1686 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1685 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_422 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1688 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1687 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1686 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1685 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1684 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1683 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1682 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1681 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_421 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1684 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1683 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1682 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1681 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_211 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_211 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_422 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_421 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_211 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1680 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1679 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1678 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1677 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_420 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1680 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1679 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1678 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1677 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1676 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1675 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1674 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1673 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_419 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1676 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1675 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1674 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1673 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_210 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_210 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_420 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_419 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_210 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1672 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1671 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1670 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1669 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_418 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1672 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1671 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1670 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1669 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1668 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1667 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1666 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1665 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_417 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1668 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1667 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1666 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1665 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_209 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_209 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_418 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_417 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_209 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_14 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_224 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_223 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_222 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_221 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_220 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_219 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_218 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_217 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_216 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_215 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_214 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), .S(S[43:40]) );
  carry_select_block_NPB4_213 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), .S(S[47:44]) );
  carry_select_block_NPB4_212 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), .S(S[51:48]) );
  carry_select_block_NPB4_211 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), .S(S[55:52]) );
  carry_select_block_NPB4_210 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), .S(S[59:56]) );
  carry_select_block_NPB4_209 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), .S(S[63:60]) );
endmodule


module P4_ADDER_N64_14 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_14 CGEN ( .A(A), .B({B[63:29], n13, B[27:21], n8, 
        B[19:17], n5, B[15:13], n11, B[11:0]}), .Cin(Cin), .Co(CoutCgen) );
  sum_generator_N64_NPB4_14 SGEN ( .A(A), .B({B[63:30], n10, B[28], n2, n4, 
        B[25:24], n7, B[22], n6, B[20], n1, B[18:16], n12, B[14:12], n9, 
        B[10:8], n14, B[6:0]}), .Ci({CoutCgen, Cin}), .S(S), .Co(Cout) );
  BUF_X1 U1 ( .A(B[29]), .Z(n10) );
  BUF_X1 U2 ( .A(B[12]), .Z(n11) );
  CLKBUF_X1 U3 ( .A(B[19]), .Z(n1) );
  CLKBUF_X1 U4 ( .A(B[27]), .Z(n2) );
  INV_X1 U5 ( .A(B[26]), .ZN(n3) );
  INV_X1 U6 ( .A(n3), .ZN(n4) );
  CLKBUF_X1 U7 ( .A(B[16]), .Z(n5) );
  BUF_X2 U8 ( .A(B[21]), .Z(n6) );
  BUF_X1 U9 ( .A(B[20]), .Z(n8) );
  CLKBUF_X1 U10 ( .A(B[23]), .Z(n7) );
  CLKBUF_X1 U11 ( .A(B[11]), .Z(n9) );
  CLKBUF_X1 U12 ( .A(B[7]), .Z(n14) );
  CLKBUF_X1 U13 ( .A(B[15]), .Z(n12) );
  CLKBUF_X1 U14 ( .A(B[28]), .Z(n13) );
endmodule


module Booth_Encoder_13 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_13 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305;

  NAND2_X1 U1 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  NAND2_X1 U2 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  NAND2_X1 U3 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  NAND2_X1 U4 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  NAND2_X1 U5 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  NOR3_X1 U6 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U7 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  NOR4_X1 U8 ( .A1(n151), .A2(n145), .A3(n154), .A4(n167), .ZN(n139) );
  BUF_X1 U9 ( .A(n152), .Z(n154) );
  BUF_X1 U10 ( .A(n165), .Z(n167) );
  AOI222_X4 U11 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n154), .ZN(n176) );
  AOI222_X1 U12 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n154), .ZN(n192) );
  CLKBUF_X1 U13 ( .A(n165), .Z(n169) );
  CLKBUF_X1 U14 ( .A(n152), .Z(n156) );
  CLKBUF_X1 U15 ( .A(n303), .Z(n166) );
  CLKBUF_X1 U16 ( .A(n302), .Z(n153) );
  BUF_X1 U17 ( .A(n139), .Z(n159) );
  BUF_X1 U18 ( .A(n139), .Z(n162) );
  BUF_X1 U19 ( .A(n139), .Z(n160) );
  BUF_X1 U20 ( .A(n139), .Z(n161) );
  BUF_X1 U21 ( .A(n139), .Z(n163) );
  BUF_X1 U22 ( .A(n153), .Z(n157) );
  BUF_X1 U23 ( .A(n166), .Z(n170) );
  BUF_X1 U24 ( .A(n152), .Z(n155) );
  BUF_X1 U25 ( .A(n165), .Z(n168) );
  BUF_X1 U26 ( .A(n153), .Z(n158) );
  BUF_X1 U27 ( .A(n166), .Z(n171) );
  BUF_X1 U28 ( .A(n303), .Z(n165) );
  BUF_X1 U29 ( .A(n302), .Z(n152) );
  CLKBUF_X1 U30 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U31 ( .A(n301), .Z(n148) );
  CLKBUF_X1 U32 ( .A(n301), .Z(n149) );
  CLKBUF_X1 U33 ( .A(n301), .Z(n147) );
  CLKBUF_X1 U34 ( .A(n301), .Z(n146) );
  CLKBUF_X1 U35 ( .A(n300), .Z(n143) );
  CLKBUF_X1 U36 ( .A(n300), .Z(n142) );
  CLKBUF_X1 U37 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U38 ( .A(n300), .Z(n141) );
  CLKBUF_X1 U39 ( .A(n300), .Z(n140) );
  INV_X1 U40 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U41 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n303) );
  AND3_X1 U42 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U43 ( .A(sel[2]), .ZN(n173) );
  AOI22_X1 U44 ( .A1(C[8]), .A2(n146), .B1(A[8]), .B2(n140), .ZN(n299) );
  NAND2_X1 U45 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U46 ( .A1(C[11]), .A2(n151), .B1(A[11]), .B2(n145), .ZN(n179) );
  NAND2_X1 U47 ( .A1(n305), .A2(n304), .ZN(Y[9]) );
  AOI22_X1 U48 ( .A1(C[9]), .A2(n148), .B1(A[9]), .B2(n142), .ZN(n305) );
  NAND2_X1 U49 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U50 ( .A1(C[10]), .A2(n151), .B1(A[10]), .B2(n145), .ZN(n177) );
  NAND2_X1 U51 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  AOI22_X1 U52 ( .A1(C[12]), .A2(n151), .B1(A[12]), .B2(n145), .ZN(n181) );
  AOI222_X1 U53 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n154), .ZN(n180) );
  NAND2_X1 U54 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  AOI22_X1 U55 ( .A1(C[40]), .A2(n148), .B1(A[40]), .B2(n142), .ZN(n243) );
  AOI222_X1 U56 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n156), .ZN(n242) );
  AOI22_X1 U57 ( .A1(C[32]), .A2(n149), .B1(A[32]), .B2(n143), .ZN(n225) );
  AOI222_X1 U58 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n156), .ZN(n224) );
  NAND2_X1 U59 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI22_X1 U60 ( .A1(C[35]), .A2(n149), .B1(A[35]), .B2(n143), .ZN(n231) );
  AOI222_X1 U61 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n156), .ZN(n230) );
  NAND2_X1 U62 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI22_X1 U63 ( .A1(C[39]), .A2(n148), .B1(A[39]), .B2(n142), .ZN(n239) );
  AOI222_X1 U64 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n156), .ZN(n238) );
  NAND2_X1 U65 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI22_X1 U66 ( .A1(C[41]), .A2(n148), .B1(A[41]), .B2(n142), .ZN(n245) );
  AOI222_X1 U67 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n156), .ZN(n244) );
  NAND2_X1 U68 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI22_X1 U69 ( .A1(C[42]), .A2(n148), .B1(A[42]), .B2(n142), .ZN(n247) );
  AOI222_X1 U70 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n156), .ZN(n246) );
  NAND2_X1 U71 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI22_X1 U72 ( .A1(C[43]), .A2(n148), .B1(A[43]), .B2(n142), .ZN(n249) );
  AOI222_X1 U73 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n156), .ZN(n248) );
  NAND2_X1 U74 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI22_X1 U75 ( .A1(C[29]), .A2(n149), .B1(A[29]), .B2(n143), .ZN(n217) );
  NAND2_X1 U76 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI22_X1 U77 ( .A1(C[45]), .A2(n148), .B1(A[45]), .B2(n142), .ZN(n253) );
  AOI222_X1 U78 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n157), .ZN(n252) );
  NAND2_X1 U79 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  AOI22_X1 U80 ( .A1(C[48]), .A2(n147), .B1(A[48]), .B2(n141), .ZN(n259) );
  AOI222_X1 U81 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n157), .ZN(n258) );
  NAND2_X1 U82 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI22_X1 U83 ( .A1(C[46]), .A2(n147), .B1(A[46]), .B2(n141), .ZN(n255) );
  AOI222_X1 U84 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n157), .ZN(n254) );
  NAND2_X1 U85 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI22_X1 U86 ( .A1(C[47]), .A2(n147), .B1(A[47]), .B2(n141), .ZN(n257) );
  AOI222_X1 U87 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n157), .ZN(n256) );
  NAND2_X1 U88 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  AOI22_X1 U89 ( .A1(C[51]), .A2(n147), .B1(A[51]), .B2(n141), .ZN(n267) );
  AOI222_X1 U90 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n157), .ZN(n266) );
  NAND2_X1 U91 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI22_X1 U92 ( .A1(C[49]), .A2(n147), .B1(A[49]), .B2(n141), .ZN(n261) );
  AOI222_X1 U93 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n157), .ZN(n260) );
  NAND2_X1 U94 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  AOI22_X1 U95 ( .A1(C[53]), .A2(n147), .B1(A[53]), .B2(n141), .ZN(n271) );
  AOI222_X1 U96 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n157), .ZN(n270) );
  NAND2_X1 U97 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI22_X1 U98 ( .A1(C[55]), .A2(n147), .B1(A[55]), .B2(n141), .ZN(n275) );
  AOI222_X1 U99 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n157), .ZN(n274) );
  AOI22_X1 U100 ( .A1(C[16]), .A2(n150), .B1(A[16]), .B2(n144), .ZN(n189) );
  AOI222_X1 U101 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n154), .ZN(n188) );
  AOI222_X1 U102 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n155), .ZN(n206) );
  AOI22_X1 U103 ( .A1(C[24]), .A2(n150), .B1(A[24]), .B2(n144), .ZN(n207) );
  NAND2_X1 U104 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI22_X1 U105 ( .A1(C[50]), .A2(n147), .B1(A[50]), .B2(n141), .ZN(n265) );
  AOI222_X1 U106 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n157), .ZN(n264) );
  NAND2_X1 U107 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  AOI22_X1 U108 ( .A1(C[52]), .A2(n147), .B1(A[52]), .B2(n141), .ZN(n269) );
  AOI222_X1 U109 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n157), .ZN(n268) );
  NAND2_X1 U110 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI22_X1 U111 ( .A1(C[54]), .A2(n147), .B1(A[54]), .B2(n141), .ZN(n273) );
  AOI222_X1 U112 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n157), .ZN(n272) );
  NAND2_X1 U113 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI22_X1 U114 ( .A1(C[17]), .A2(n150), .B1(A[17]), .B2(n144), .ZN(n191) );
  AOI222_X1 U115 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n154), .ZN(n190) );
  NAND2_X1 U116 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U117 ( .A1(C[15]), .A2(n150), .B1(A[15]), .B2(n144), .ZN(n187) );
  AOI222_X1 U118 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n154), .ZN(n186) );
  NAND2_X1 U119 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI22_X1 U120 ( .A1(C[18]), .A2(n150), .B1(A[18]), .B2(n144), .ZN(n193) );
  NAND2_X1 U121 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI222_X1 U122 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n154), .ZN(n194) );
  AOI22_X1 U123 ( .A1(C[19]), .A2(n150), .B1(A[19]), .B2(n144), .ZN(n195) );
  NAND2_X1 U124 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI222_X1 U125 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n155), .ZN(n204) );
  AOI22_X1 U126 ( .A1(C[23]), .A2(n150), .B1(A[23]), .B2(n144), .ZN(n205) );
  NAND2_X1 U127 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI22_X1 U128 ( .A1(C[37]), .A2(n148), .B1(A[37]), .B2(n142), .ZN(n235) );
  NAND2_X1 U129 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U130 ( .A1(C[30]), .A2(n149), .B1(A[30]), .B2(n143), .ZN(n221) );
  NAND2_X1 U131 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI22_X1 U132 ( .A1(C[33]), .A2(n149), .B1(A[33]), .B2(n143), .ZN(n227) );
  NAND2_X1 U133 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI22_X1 U134 ( .A1(C[34]), .A2(n149), .B1(A[34]), .B2(n143), .ZN(n229) );
  NAND2_X1 U135 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI222_X1 U136 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n156), .ZN(n236) );
  AOI22_X1 U137 ( .A1(C[38]), .A2(n148), .B1(A[38]), .B2(n142), .ZN(n237) );
  NAND2_X1 U138 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  AOI22_X1 U139 ( .A1(C[44]), .A2(n148), .B1(A[44]), .B2(n142), .ZN(n251) );
  AOI222_X1 U140 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n157), .ZN(n250) );
  NAND2_X1 U141 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  AOI222_X1 U142 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n155), .ZN(n198) );
  AOI22_X1 U143 ( .A1(C[20]), .A2(n150), .B1(A[20]), .B2(n144), .ZN(n199) );
  NAND2_X1 U144 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI222_X1 U145 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n155), .ZN(n210) );
  AOI22_X1 U146 ( .A1(C[26]), .A2(n149), .B1(A[26]), .B2(n143), .ZN(n211) );
  NAND2_X1 U147 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U148 ( .A1(C[13]), .A2(n151), .B1(A[13]), .B2(n145), .ZN(n183) );
  AOI222_X1 U149 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n154), .ZN(n182) );
  NAND2_X1 U150 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI222_X1 U151 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n155), .ZN(n200) );
  AOI22_X1 U152 ( .A1(C[21]), .A2(n150), .B1(A[21]), .B2(n144), .ZN(n201) );
  NAND2_X1 U153 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI222_X1 U154 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n155), .ZN(n208) );
  AOI22_X1 U155 ( .A1(C[25]), .A2(n149), .B1(A[25]), .B2(n143), .ZN(n209) );
  NAND2_X1 U156 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U157 ( .A1(C[14]), .A2(n150), .B1(A[14]), .B2(n144), .ZN(n185) );
  AOI222_X1 U158 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n154), .ZN(n184) );
  NAND2_X1 U159 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI22_X1 U160 ( .A1(C[22]), .A2(n150), .B1(A[22]), .B2(n144), .ZN(n203) );
  AOI222_X1 U161 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n155), .ZN(n202) );
  AOI222_X1 U162 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n156), .ZN(n232) );
  AOI22_X1 U163 ( .A1(C[36]), .A2(n148), .B1(A[36]), .B2(n142), .ZN(n233) );
  NAND2_X1 U164 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  AOI22_X1 U165 ( .A1(C[28]), .A2(n149), .B1(A[28]), .B2(n143), .ZN(n215) );
  AOI222_X1 U166 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n155), .ZN(n214) );
  NAND2_X1 U167 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI222_X1 U168 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n155), .ZN(n212) );
  AOI22_X1 U169 ( .A1(C[27]), .A2(n149), .B1(A[27]), .B2(n143), .ZN(n213) );
  NAND2_X1 U170 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI222_X1 U171 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n155), .ZN(n222) );
  AOI22_X1 U172 ( .A1(C[31]), .A2(n149), .B1(A[31]), .B2(n143), .ZN(n223) );
  NAND2_X1 U173 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI22_X1 U174 ( .A1(C[58]), .A2(n146), .B1(A[58]), .B2(n140), .ZN(n281) );
  AOI222_X1 U175 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n158), .ZN(n280) );
  NAND2_X1 U176 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  AOI22_X1 U177 ( .A1(C[57]), .A2(n146), .B1(A[57]), .B2(n140), .ZN(n279) );
  AOI222_X1 U178 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n158), .ZN(n278) );
  NAND2_X1 U179 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  AOI22_X1 U180 ( .A1(C[56]), .A2(n147), .B1(A[56]), .B2(n141), .ZN(n277) );
  AOI222_X1 U181 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n158), .ZN(n276) );
  NAND2_X1 U182 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U183 ( .A1(C[60]), .A2(n146), .B1(A[60]), .B2(n140), .ZN(n287) );
  AOI222_X1 U184 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n158), .ZN(n286) );
  NAND2_X1 U185 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U186 ( .A1(C[61]), .A2(n146), .B1(A[61]), .B2(n140), .ZN(n289) );
  AOI222_X1 U187 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n158), .ZN(n288) );
  NAND2_X1 U188 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U189 ( .A1(C[59]), .A2(n146), .B1(A[59]), .B2(n140), .ZN(n283) );
  AOI222_X1 U190 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n158), .ZN(n282) );
  NAND2_X1 U191 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U192 ( .A1(C[62]), .A2(n146), .B1(A[62]), .B2(n140), .ZN(n291) );
  AOI222_X1 U193 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n158), .ZN(n290) );
  NAND2_X1 U194 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U195 ( .A1(C[63]), .A2(n146), .B1(A[63]), .B2(n140), .ZN(n293) );
  AOI222_X1 U196 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n158), .ZN(n292) );
  NAND2_X1 U197 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U198 ( .A1(C[0]), .A2(n146), .B1(A[0]), .B2(n140), .ZN(n175) );
  AOI222_X1 U199 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n154), .ZN(n174) );
  NAND2_X1 U200 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U201 ( .A1(C[4]), .A2(n147), .B1(A[4]), .B2(n141), .ZN(n263) );
  AOI222_X1 U202 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n157), .ZN(n262) );
  NAND2_X1 U203 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U204 ( .A1(C[1]), .A2(n150), .B1(A[1]), .B2(n144), .ZN(n197) );
  AOI222_X1 U205 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n154), .ZN(n196) );
  NAND2_X1 U206 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U207 ( .A1(C[5]), .A2(n146), .B1(A[5]), .B2(n140), .ZN(n285) );
  AOI222_X1 U208 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n158), .ZN(n284) );
  NAND2_X1 U209 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U210 ( .A1(C[2]), .A2(n149), .B1(A[2]), .B2(n143), .ZN(n219) );
  AOI222_X1 U211 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n155), .ZN(n218) );
  NAND2_X1 U212 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U213 ( .A1(C[3]), .A2(n148), .B1(A[3]), .B2(n142), .ZN(n241) );
  AOI222_X1 U214 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n156), .ZN(n240) );
  AOI222_X1 U215 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n156), .ZN(n226) );
  AOI222_X1 U216 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n158), .ZN(n294) );
  AOI22_X1 U217 ( .A1(C[6]), .A2(n146), .B1(A[6]), .B2(n140), .ZN(n295) );
  NAND2_X1 U218 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  NAND2_X1 U219 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U220 ( .A1(C[7]), .A2(n146), .B1(A[7]), .B2(n140), .ZN(n297) );
  AOI222_X1 U221 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n158), .ZN(n298) );
  AOI222_X1 U222 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n154), .ZN(n178) );
  AOI222_X1 U223 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n156), .ZN(n228) );
  AOI222_X1 U224 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n158), .ZN(n296) );
  AOI222_X1 U225 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n155), .ZN(n216) );
  AOI222_X1 U226 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n155), .ZN(n220) );
  AOI222_X1 U227 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n156), .ZN(n234) );
  AOI222_X1 U228 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n158), .ZN(n304) );
  CLKBUF_X1 U229 ( .A(n300), .Z(n145) );
  CLKBUF_X1 U230 ( .A(n301), .Z(n151) );
  CLKBUF_X1 U231 ( .A(n139), .Z(n164) );
endmodule


module G_221 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_819 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_818 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_817 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3, n5;

  CLKBUF_X1 U1 ( .A(P_IK), .Z(n3) );
  INV_X1 U2 ( .A(n5), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n5) );
  AND2_X1 U4 ( .A1(P_K_1), .A2(n3), .ZN(Px) );
endmodule


module PG_816 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_815 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_814 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_813 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_812 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_811 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_810 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_809 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_808 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_807 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_806 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_805 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_804 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_803 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_802 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_801 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_800 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_799 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_798 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_797 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_796 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_795 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_794 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_793 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_792 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_791 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_790 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_789 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_220 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_788 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_787 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_786 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_785 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_784 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_783 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_782 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_781 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_780 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_779 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_778 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_777 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_776 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_775 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_774 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_219 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_773 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_772 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_771 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_770 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_769 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_768 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_767 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_218 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_217 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
endmodule


module PG_766 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_765 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_764 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_763 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_762 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_761 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_216 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_215 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_214 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
endmodule


module G_213 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_760 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_759 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_758 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_757 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_212 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_211 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_210 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_209 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_208 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_207 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_206 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_205 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module carry_generator_N64_NPB4_13 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   n22, \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n11, n12, n14, n15, n16, n17, n18, n19, n20, n21;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U77 ( .A(B[59]), .B(A[59]), .Z(\PG_Network[0][0][59] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U81 ( .A(B[55]), .B(A[55]), .Z(\PG_Network[0][0][55] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U85 ( .A(B[51]), .B(A[51]), .Z(\PG_Network[0][0][51] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U88 ( .A(B[49]), .B(A[49]), .Z(\PG_Network[0][0][49] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U90 ( .A(B[47]), .B(A[47]), .Z(\PG_Network[0][0][47] ) );
  XOR2_X1 U91 ( .A(B[46]), .B(A[46]), .Z(\PG_Network[0][0][46] ) );
  XOR2_X1 U92 ( .A(B[45]), .B(A[45]), .Z(\PG_Network[0][0][45] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U94 ( .A(B[43]), .B(A[43]), .Z(\PG_Network[0][0][43] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U100 ( .A(B[38]), .B(A[38]), .Z(\PG_Network[0][0][38] ) );
  XOR2_X1 U101 ( .A(B[37]), .B(A[37]), .Z(\PG_Network[0][0][37] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U108 ( .A(B[30]), .B(A[30]), .Z(\PG_Network[0][0][30] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U110 ( .A(B[29]), .B(A[29]), .Z(\PG_Network[0][0][29] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U114 ( .A(B[25]), .B(A[25]), .Z(\PG_Network[0][0][25] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_221 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n18), .Gx(\PG_Network[1][1][1] ) );
  PG_819 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_818 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_817 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_816 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_815 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_814 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_813 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_812 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_811 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_810 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_809 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_808 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_807 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_806 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_805 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_804 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_803 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_802 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_801 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_800 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_799 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_798 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_797 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_796 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_795 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_794 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_793 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_792 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_791 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_790 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_789 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_220 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_788 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_787 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_786 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_785 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_784 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_783 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_782 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_781 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_780 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_779 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_778 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_777 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_776 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_775 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_774 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_219 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_773 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_772 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_771 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_770 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_769 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_768 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_767 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_218 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), .G_K_1(Co[1]), .Gx(n22) );
  G_217 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_766 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_765 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_764 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][47] ), .Px(
        \PG_Network[4][0][47] ) );
  PG_763 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][43] ), .Px(
        \PG_Network[4][0][43] ) );
  PG_762 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][63] ), .Px(
        \PG_Network[4][0][63] ) );
  PG_761 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][59] ), .Px(
        \PG_Network[4][0][59] ) );
  G_216 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), .G_K_1(n15), .Gx(Co[7]) );
  G_215 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), .G_K_1(n15), .Gx(Co[6]) );
  G_214 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), .G_K_1(Co[3]), .Gx(Co[5]) );
  G_213 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), .G_K_1(n22), .Gx(Co[4]) );
  PG_760 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][63] ), .Px(
        \PG_Network[5][0][63] ) );
  PG_759 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][59] ), .Px(
        \PG_Network[5][0][59] ) );
  PG_758 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][55] ), .Px(
        \PG_Network[5][0][55] ) );
  PG_757 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][51] ), .Px(
        \PG_Network[5][0][51] ) );
  G_212 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), .G_K_1(n5), .Gx(Co[15]) );
  G_211 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), .G_K_1(n5), .Gx(Co[14]) );
  G_210 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), .G_K_1(n5), .Gx(Co[13]) );
  G_209 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), .G_K_1(n5), .Gx(Co[12]) );
  G_208 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), .G_K_1(n5), .Gx(Co[11]) );
  G_207 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), .G_K_1(n16), .Gx(Co[10]) );
  G_206 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), .G_K_1(n16), .Gx(Co[9]) );
  G_205 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), .G_K_1(Co[7]), .Gx(Co[8]) );
  BUF_X1 U1 ( .A(n22), .Z(Co[3]) );
  INV_X1 U2 ( .A(A[11]), .ZN(n11) );
  INV_X1 U3 ( .A(A[35]), .ZN(n17) );
  INV_X1 U4 ( .A(A[27]), .ZN(n14) );
  INV_X1 U5 ( .A(A[31]), .ZN(n7) );
  INV_X1 U6 ( .A(A[39]), .ZN(n6) );
  INV_X1 U7 ( .A(A[15]), .ZN(n12) );
  INV_X1 U8 ( .A(A[19]), .ZN(n9) );
  INV_X1 U9 ( .A(A[23]), .ZN(n10) );
  INV_X1 U10 ( .A(A[7]), .ZN(n8) );
  CLKBUF_X1 U11 ( .A(n16), .Z(n5) );
  CLKBUF_X1 U12 ( .A(Co[7]), .Z(n16) );
  XNOR2_X1 U13 ( .A(B[39]), .B(n6), .ZN(\PG_Network[0][0][39] ) );
  CLKBUF_X1 U14 ( .A(Co[3]), .Z(n15) );
  XNOR2_X1 U15 ( .A(B[31]), .B(n7), .ZN(\PG_Network[0][0][31] ) );
  XNOR2_X1 U16 ( .A(B[7]), .B(n8), .ZN(\PG_Network[0][0][7] ) );
  XNOR2_X1 U17 ( .A(B[19]), .B(n9), .ZN(\PG_Network[0][0][19] ) );
  XNOR2_X1 U18 ( .A(B[23]), .B(n10), .ZN(\PG_Network[0][0][23] ) );
  XNOR2_X1 U19 ( .A(B[11]), .B(n11), .ZN(\PG_Network[0][0][11] ) );
  XNOR2_X1 U20 ( .A(B[15]), .B(n12), .ZN(\PG_Network[0][0][15] ) );
  XNOR2_X1 U21 ( .A(B[27]), .B(n14), .ZN(\PG_Network[0][0][27] ) );
  XNOR2_X1 U22 ( .A(B[35]), .B(n17), .ZN(\PG_Network[0][0][35] ) );
  AND2_X1 U23 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U24 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U25 ( .A1(A[11]), .A2(B[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U26 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U27 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U28 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U29 ( .A1(A[43]), .A2(B[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U30 ( .A1(A[41]), .A2(B[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U31 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U32 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U33 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U34 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U35 ( .A1(B[19]), .A2(A[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U36 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AND2_X1 U37 ( .A1(B[13]), .A2(A[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U38 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U39 ( .A1(B[15]), .A2(A[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U40 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U41 ( .A1(B[7]), .A2(A[7]), .ZN(\PG_Network[0][1][7] ) );
  AND2_X1 U42 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U43 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U44 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U45 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U46 ( .A1(A[25]), .A2(B[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U47 ( .A1(A[46]), .A2(B[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U48 ( .A1(A[47]), .A2(B[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U49 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U50 ( .A1(A[45]), .A2(B[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U51 ( .A1(A[49]), .A2(B[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U52 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U53 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U54 ( .A1(A[51]), .A2(B[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U55 ( .A1(A[29]), .A2(B[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U56 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AND2_X1 U57 ( .A1(B[23]), .A2(A[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U58 ( .A1(A[37]), .A2(B[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U59 ( .A1(B[21]), .A2(A[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U60 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U61 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U62 ( .A1(A[59]), .A2(B[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U63 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
  AND2_X1 U64 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U65 ( .A1(A[53]), .A2(B[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U66 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U67 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U70 ( .A1(A[55]), .A2(B[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U99 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U103 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U107 ( .A(n21), .ZN(n18) );
  AND2_X1 U112 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U116 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U121 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U125 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U129 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U131 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U132 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AOI21_X1 U133 ( .B1(A[0]), .B2(B[0]), .A(n19), .ZN(n21) );
  INV_X1 U134 ( .A(n20), .ZN(n19) );
  OAI21_X1 U135 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n20) );
  AND2_X1 U136 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U137 ( .A1(A[27]), .A2(B[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U138 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U139 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U140 ( .A1(A[31]), .A2(B[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U141 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U142 ( .A1(A[35]), .A2(B[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U143 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
endmodule


module FA_1664 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1663 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1662 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1661 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_416 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1664 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1663 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1662 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1661 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1660 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1659 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1658 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1657 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_415 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1660 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1659 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1658 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1657 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_208 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U2 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_208 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_416 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_415 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_208 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1656 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1655 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1654 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1653 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_414 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1656 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1655 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1654 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1653 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1652 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1651 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1650 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1649 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_413 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1652 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1651 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1650 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1649 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_207 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_207 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_414 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_413 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_207 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1648 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_1647 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1646 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1645 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  OR2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n6) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n8) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_412 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1648 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1647 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1646 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1645 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1644 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1643 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(n4), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1642 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1641 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_411 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1644 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1643 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1642 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1641 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_206 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U5 ( .A(sel), .ZN(n13) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n13), .ZN(n17) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_206 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_412 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_411 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_206 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1640 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  XOR2_X1 U2 ( .A(A), .B(n4), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1639 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1638 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1637 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(n4), .ZN(n7) );
endmodule


module RCA_N4_410 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1640 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1639 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1638 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1637 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1636 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1635 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1634 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1633 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_409 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1636 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1635 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1634 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1633 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_205 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19, n20;

  INV_X1 U1 ( .A(n19), .ZN(Y[2]) );
  INV_X1 U2 ( .A(n18), .ZN(Y[1]) );
  BUF_X1 U3 ( .A(n11), .Z(n5) );
  INV_X1 U4 ( .A(n5), .ZN(n10) );
  INV_X1 U5 ( .A(n17), .ZN(Y[0]) );
  INV_X1 U6 ( .A(sel), .ZN(n11) );
  INV_X1 U7 ( .A(n20), .ZN(Y[3]) );
  INV_X1 U8 ( .A(sel), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n20) );
  AOI22_X1 U10 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n19) );
  AOI22_X1 U11 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n11), .ZN(n18) );
  AOI22_X1 U12 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n16), .ZN(n17) );
endmodule


module carry_select_block_NPB4_205 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_410 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_409 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_205 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1632 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1631 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1630 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1629 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_408 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1632 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1631 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1630 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1629 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1628 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1627 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1626 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1625 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_407 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1628 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1627 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1626 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1625 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_204 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n17), .ZN(Y[1]) );
  BUF_X1 U2 ( .A(n15), .Z(n10) );
  INV_X1 U3 ( .A(n18), .ZN(Y[2]) );
  CLKBUF_X1 U4 ( .A(sel), .Z(n5) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U7 ( .A(sel), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n10), .ZN(n19) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[1]), .B1(n15), .B2(B[1]), .ZN(n17) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_204 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_408 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_407 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_204 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1624 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n4), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_1623 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net69247, n4, n5;
  assign Co = net69247;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(net69247) );
endmodule


module FA_1622 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1621 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  OR2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_406 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1624 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1623 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1622 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1621 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1620 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1619 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(n4), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1618 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1617 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_405 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1620 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1619 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1618 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1617 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_203 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U5 ( .A(sel), .ZN(n10) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n10), .ZN(n17) );
  INV_X1 U8 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n10), .ZN(n19) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_203 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_406 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_405 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_203 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1616 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_1615 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1614 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1613 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_404 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1616 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1615 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1614 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1613 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1612 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1611 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1610 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1609 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_403 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1612 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1611 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1610 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1609 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_202 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n12, n17, n18, n19, n20, n21;

  BUF_X1 U1 ( .A(sel), .Z(n12) );
  BUF_X1 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(n20), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n21), .ZN(Y[3]) );
  INV_X1 U5 ( .A(n10), .ZN(n5) );
  INV_X1 U6 ( .A(n19), .ZN(Y[1]) );
  INV_X1 U7 ( .A(n18), .ZN(Y[0]) );
  INV_X1 U8 ( .A(sel), .ZN(n11) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(n12), .B1(n17), .B2(B[2]), .ZN(n20) );
  AOI22_X1 U10 ( .A1(n12), .A2(A[1]), .B1(B[1]), .B2(n5), .ZN(n19) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n11), .B2(B[0]), .ZN(n18) );
  INV_X1 U12 ( .A(n10), .ZN(n17) );
  AOI22_X1 U13 ( .A1(A[3]), .A2(n12), .B1(B[3]), .B2(n17), .ZN(n21) );
endmodule


module carry_select_block_NPB4_202 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_404 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_403 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_202 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1608 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n5) );
  AOI22_X1 U5 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_1607 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1606 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1605 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_402 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1608 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1607 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1606 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1605 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1604 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1603 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1602 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1601 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_401 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1604 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1603 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1602 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1601 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_201 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U2 ( .A(sel), .ZN(n5) );
  INV_X1 U3 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n17) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n18) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n14), .ZN(n15) );
  INV_X1 U10 ( .A(sel), .ZN(n14) );
endmodule


module carry_select_block_NPB4_201 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_402 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_401 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_201 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1600 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(n4), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_1599 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1598 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1597 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_400 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1600 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1599 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1598 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1597 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1596 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1595 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1594 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1593 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_399 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1596 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1595 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1594 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1593 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_200 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n16), .ZN(Y[1]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n5) );
  INV_X2 U3 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U5 ( .A(sel), .ZN(n14) );
  INV_X1 U6 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n14), .ZN(n17) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(n5), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n14), .ZN(n18) );
endmodule


module carry_select_block_NPB4_200 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_400 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_399 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_200 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1592 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_1591 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1590 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1589 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_398 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1592 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1591 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1590 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1589 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1588 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1587 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1586 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1585 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_397 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1588 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1587 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1586 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1585 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_199 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(sel), .Z(n10) );
  INV_X1 U2 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U5 ( .A(sel), .ZN(n5) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n5), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n15), .ZN(n17) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(n10), .A2(A[3]), .B1(B[3]), .B2(n15), .ZN(n19) );
endmodule


module carry_select_block_NPB4_199 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_398 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_397 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_199 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1584 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1583 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1582 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1581 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_396 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1584 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1583 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1582 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1581 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1580 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1579 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1578 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1577 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_395 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1580 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1579 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1578 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1577 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_198 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U2 ( .A(sel), .ZN(n5) );
  INV_X1 U3 ( .A(n16), .ZN(Y[0]) );
  BUF_X1 U4 ( .A(n5), .Z(n10) );
  CLKBUF_X1 U5 ( .A(sel), .Z(n11) );
  INV_X1 U6 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U7 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n11), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n10), .ZN(n17) );
  AOI22_X1 U10 ( .A1(n11), .A2(A[3]), .B1(B[3]), .B2(n10), .ZN(n19) );
  AOI22_X1 U11 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n5), .ZN(n16) );
endmodule


module carry_select_block_NPB4_198 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_396 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_395 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_198 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1576 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1575 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1574 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1573 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_394 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1576 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1575 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1574 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1573 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1572 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1571 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1570 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1569 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_393 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1572 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1571 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1570 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1569 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_197 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  CLKBUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(n5), .ZN(n10) );
  INV_X1 U3 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U4 ( .A1(n5), .A2(A[3]), .B1(B[3]), .B2(n10), .ZN(n19) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n10), .ZN(n18) );
  INV_X1 U7 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(n5), .B1(B[1]), .B2(n15), .ZN(n17) );
  INV_X1 U9 ( .A(n16), .ZN(Y[0]) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_197 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_394 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_393 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_197 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1568 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1567 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1566 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1565 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_392 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1568 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1567 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1566 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1565 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1564 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1563 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1562 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1561 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_391 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1564 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1563 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1562 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1561 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_196 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(sel), .ZN(n13) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_196 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_392 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_391 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_196 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1560 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1559 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1558 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1557 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_390 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1560 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1559 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1558 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1557 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1556 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1555 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1554 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1553 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_389 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1556 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1555 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1554 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1553 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_195 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_195 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_390 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_389 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_195 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1552 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1551 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1550 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1549 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_388 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1552 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1551 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1550 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1549 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1548 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1547 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1546 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1545 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_387 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1548 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1547 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1546 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1545 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_194 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_194 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_388 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_387 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_194 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1544 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1543 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1542 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1541 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_386 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1544 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1543 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1542 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1541 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1540 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1539 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1538 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1537 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_385 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1540 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1539 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1538 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1537 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_193 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_193 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_386 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_385 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_193 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_13 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_208 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_207 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_206 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_205 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_204 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_203 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_202 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_201 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_200 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_199 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_198 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), .S(S[43:40]) );
  carry_select_block_NPB4_197 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), .S(S[47:44]) );
  carry_select_block_NPB4_196 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), .S(S[51:48]) );
  carry_select_block_NPB4_195 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), .S(S[55:52]) );
  carry_select_block_NPB4_194 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), .S(S[59:56]) );
  carry_select_block_NPB4_193 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), .S(S[63:60]) );
endmodule


module P4_ADDER_N64_13 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_13 CGEN ( .A(A), .B({B[63:37], n12, B[35:21], n15, 
        B[19:17], n11, B[15:0]}), .Cin(Cin), .Co(CoutCgen) );
  sum_generator_N64_NPB4_13 SGEN ( .A(A), .B({B[63:40], n14, B[38:32], n6, n8, 
        B[29:28], n4, B[26:24], n3, B[22:20], n5, B[18:16], n1, B[14:12], n10, 
        B[10:8], n2, B[6:0]}), .Ci({CoutCgen, Cin}), .S(S), .Co(Cout) );
  CLKBUF_X1 U1 ( .A(B[15]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(B[7]), .Z(n2) );
  CLKBUF_X1 U3 ( .A(B[23]), .Z(n3) );
  CLKBUF_X1 U4 ( .A(B[27]), .Z(n4) );
  CLKBUF_X1 U5 ( .A(B[19]), .Z(n5) );
  CLKBUF_X1 U6 ( .A(B[31]), .Z(n6) );
  INV_X1 U7 ( .A(B[30]), .ZN(n7) );
  INV_X1 U8 ( .A(n7), .ZN(n8) );
  INV_X1 U9 ( .A(B[11]), .ZN(n9) );
  INV_X1 U10 ( .A(n9), .ZN(n10) );
  CLKBUF_X1 U11 ( .A(B[16]), .Z(n11) );
  CLKBUF_X1 U12 ( .A(B[36]), .Z(n12) );
  INV_X1 U13 ( .A(B[39]), .ZN(n13) );
  INV_X1 U14 ( .A(n13), .ZN(n14) );
  CLKBUF_X1 U15 ( .A(B[20]), .Z(n15) );
endmodule


module Booth_Encoder_12 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_12 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305;

  NAND2_X1 U1 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  NAND2_X1 U2 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  NAND2_X1 U3 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  NAND2_X1 U4 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  NOR4_X1 U5 ( .A1(n151), .A2(n145), .A3(n154), .A4(n167), .ZN(n139) );
  NOR3_X1 U6 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U7 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  NAND2_X2 U8 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  NAND2_X2 U9 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  CLKBUF_X1 U10 ( .A(n165), .Z(n169) );
  CLKBUF_X1 U11 ( .A(n152), .Z(n156) );
  CLKBUF_X1 U12 ( .A(n165), .Z(n168) );
  CLKBUF_X1 U13 ( .A(n152), .Z(n155) );
  CLKBUF_X1 U14 ( .A(n303), .Z(n166) );
  CLKBUF_X1 U15 ( .A(n302), .Z(n153) );
  BUF_X1 U16 ( .A(n139), .Z(n161) );
  BUF_X1 U17 ( .A(n139), .Z(n160) );
  BUF_X1 U18 ( .A(n139), .Z(n162) );
  BUF_X1 U19 ( .A(n139), .Z(n159) );
  BUF_X1 U20 ( .A(n139), .Z(n163) );
  BUF_X1 U21 ( .A(n153), .Z(n157) );
  BUF_X1 U22 ( .A(n166), .Z(n170) );
  BUF_X1 U23 ( .A(n153), .Z(n158) );
  BUF_X1 U24 ( .A(n166), .Z(n171) );
  BUF_X1 U25 ( .A(n152), .Z(n154) );
  BUF_X1 U26 ( .A(n165), .Z(n167) );
  CLKBUF_X1 U27 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U28 ( .A(n301), .Z(n149) );
  CLKBUF_X1 U29 ( .A(n301), .Z(n148) );
  CLKBUF_X1 U30 ( .A(n301), .Z(n146) );
  BUF_X1 U31 ( .A(n303), .Z(n165) );
  BUF_X1 U32 ( .A(n302), .Z(n152) );
  CLKBUF_X1 U33 ( .A(n301), .Z(n147) );
  CLKBUF_X1 U34 ( .A(n300), .Z(n143) );
  CLKBUF_X1 U35 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U36 ( .A(n300), .Z(n141) );
  CLKBUF_X1 U37 ( .A(n300), .Z(n140) );
  CLKBUF_X1 U38 ( .A(n300), .Z(n142) );
  INV_X1 U39 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U40 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n303) );
  AND3_X1 U41 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U42 ( .A(sel[2]), .ZN(n173) );
  NAND2_X1 U43 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U44 ( .A1(C[11]), .A2(n151), .B1(A[11]), .B2(n145), .ZN(n179) );
  NAND2_X1 U45 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U46 ( .A1(C[10]), .A2(n151), .B1(A[10]), .B2(n145), .ZN(n177) );
  AOI22_X1 U47 ( .A1(C[12]), .A2(n151), .B1(A[12]), .B2(n145), .ZN(n181) );
  AOI222_X1 U48 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n154), .ZN(n180) );
  NAND2_X1 U49 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U50 ( .A1(C[15]), .A2(n150), .B1(A[15]), .B2(n144), .ZN(n187) );
  AOI222_X1 U51 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n154), .ZN(n186) );
  NAND2_X1 U52 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U53 ( .A1(C[14]), .A2(n150), .B1(A[14]), .B2(n144), .ZN(n185) );
  AOI222_X1 U54 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n154), .ZN(n184) );
  NAND2_X1 U55 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  AOI22_X1 U56 ( .A1(C[16]), .A2(n150), .B1(A[16]), .B2(n144), .ZN(n189) );
  AOI222_X1 U57 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n154), .ZN(n188) );
  AOI22_X1 U58 ( .A1(C[24]), .A2(n150), .B1(A[24]), .B2(n144), .ZN(n207) );
  AOI222_X1 U59 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n155), .ZN(n206) );
  NAND2_X1 U60 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  AOI22_X1 U61 ( .A1(C[28]), .A2(n149), .B1(A[28]), .B2(n143), .ZN(n215) );
  AOI222_X1 U62 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n155), .ZN(n214) );
  NAND2_X1 U63 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI22_X1 U64 ( .A1(C[23]), .A2(n150), .B1(A[23]), .B2(n144), .ZN(n205) );
  AOI222_X1 U65 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n155), .ZN(n204) );
  NAND2_X1 U66 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI22_X1 U67 ( .A1(C[26]), .A2(n149), .B1(A[26]), .B2(n143), .ZN(n211) );
  AOI222_X1 U68 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n155), .ZN(n210) );
  NAND2_X1 U69 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI22_X1 U70 ( .A1(C[27]), .A2(n149), .B1(A[27]), .B2(n143), .ZN(n213) );
  AOI222_X1 U71 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n155), .ZN(n212) );
  NAND2_X1 U72 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI22_X1 U73 ( .A1(C[31]), .A2(n149), .B1(A[31]), .B2(n143), .ZN(n223) );
  AOI222_X1 U74 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n155), .ZN(n222) );
  AOI222_X1 U75 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n158), .ZN(n298) );
  NAND2_X1 U76 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  AOI22_X1 U77 ( .A1(C[48]), .A2(n147), .B1(A[48]), .B2(n141), .ZN(n259) );
  AOI222_X1 U78 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n157), .ZN(n258) );
  NAND2_X1 U79 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI22_X1 U80 ( .A1(C[45]), .A2(n148), .B1(A[45]), .B2(n142), .ZN(n253) );
  AOI222_X1 U81 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n157), .ZN(n252) );
  NAND2_X1 U82 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI22_X1 U83 ( .A1(C[49]), .A2(n147), .B1(A[49]), .B2(n141), .ZN(n261) );
  AOI222_X1 U84 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n157), .ZN(n260) );
  NAND2_X1 U85 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI22_X1 U86 ( .A1(C[46]), .A2(n147), .B1(A[46]), .B2(n141), .ZN(n255) );
  AOI222_X1 U87 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n157), .ZN(n254) );
  NAND2_X1 U88 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI22_X1 U89 ( .A1(C[47]), .A2(n147), .B1(A[47]), .B2(n141), .ZN(n257) );
  AOI222_X1 U90 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n157), .ZN(n256) );
  NAND2_X1 U91 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  AOI22_X1 U92 ( .A1(C[52]), .A2(n147), .B1(A[52]), .B2(n141), .ZN(n269) );
  AOI222_X1 U93 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n157), .ZN(n268) );
  NAND2_X1 U94 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  AOI22_X1 U95 ( .A1(C[53]), .A2(n147), .B1(A[53]), .B2(n141), .ZN(n271) );
  AOI222_X1 U96 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n157), .ZN(n270) );
  NAND2_X1 U97 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI22_X1 U98 ( .A1(C[50]), .A2(n147), .B1(A[50]), .B2(n141), .ZN(n265) );
  AOI222_X1 U99 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n157), .ZN(n264) );
  NAND2_X1 U100 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI22_X1 U101 ( .A1(C[54]), .A2(n147), .B1(A[54]), .B2(n141), .ZN(n273) );
  AOI222_X1 U102 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n157), .ZN(n272) );
  NAND2_X1 U103 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  AOI22_X1 U104 ( .A1(C[51]), .A2(n147), .B1(A[51]), .B2(n141), .ZN(n267) );
  AOI222_X1 U105 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n157), .ZN(n266) );
  NAND2_X1 U106 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI22_X1 U107 ( .A1(C[55]), .A2(n147), .B1(A[55]), .B2(n141), .ZN(n275) );
  AOI222_X1 U108 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n157), .ZN(n274) );
  NAND2_X1 U109 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI22_X1 U110 ( .A1(C[34]), .A2(n149), .B1(A[34]), .B2(n143), .ZN(n229) );
  AOI222_X1 U111 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n156), .ZN(n228) );
  NAND2_X1 U112 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U113 ( .A1(C[30]), .A2(n149), .B1(A[30]), .B2(n143), .ZN(n221) );
  AOI222_X1 U114 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n155), .ZN(n220) );
  NAND2_X1 U115 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  AOI22_X1 U116 ( .A1(C[44]), .A2(n148), .B1(A[44]), .B2(n142), .ZN(n251) );
  AOI222_X1 U117 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n157), .ZN(n250) );
  NAND2_X1 U118 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI22_X1 U119 ( .A1(C[43]), .A2(n148), .B1(A[43]), .B2(n142), .ZN(n249) );
  AOI222_X1 U120 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n156), .ZN(n248) );
  NAND2_X1 U121 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI22_X1 U122 ( .A1(C[19]), .A2(n150), .B1(A[19]), .B2(n144), .ZN(n195) );
  AOI222_X1 U123 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n154), .ZN(n194) );
  NAND2_X1 U124 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI222_X1 U125 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n156), .ZN(n230) );
  AOI22_X1 U126 ( .A1(C[35]), .A2(n149), .B1(A[35]), .B2(n143), .ZN(n231) );
  NAND2_X1 U127 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U128 ( .A1(C[13]), .A2(n151), .B1(A[13]), .B2(n145), .ZN(n183) );
  NAND2_X1 U129 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI22_X1 U130 ( .A1(C[18]), .A2(n150), .B1(A[18]), .B2(n144), .ZN(n193) );
  AOI222_X1 U131 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n154), .ZN(n192) );
  NAND2_X1 U132 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI22_X1 U133 ( .A1(C[22]), .A2(n150), .B1(A[22]), .B2(n144), .ZN(n203) );
  AOI222_X1 U134 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n155), .ZN(n202) );
  NAND2_X1 U135 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI22_X1 U136 ( .A1(C[38]), .A2(n148), .B1(A[38]), .B2(n142), .ZN(n237) );
  AOI222_X1 U137 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n156), .ZN(n236) );
  NAND2_X1 U138 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI22_X1 U139 ( .A1(C[41]), .A2(n148), .B1(A[41]), .B2(n142), .ZN(n245) );
  AOI222_X1 U140 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n156), .ZN(n244) );
  NAND2_X1 U141 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI22_X1 U142 ( .A1(C[42]), .A2(n148), .B1(A[42]), .B2(n142), .ZN(n247) );
  AOI222_X1 U143 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n156), .ZN(n246) );
  AOI22_X1 U144 ( .A1(C[20]), .A2(n150), .B1(A[20]), .B2(n144), .ZN(n199) );
  AOI222_X1 U145 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n155), .ZN(n198) );
  NAND2_X1 U146 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI222_X1 U147 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n155), .ZN(n200) );
  AOI22_X1 U148 ( .A1(C[21]), .A2(n150), .B1(A[21]), .B2(n144), .ZN(n201) );
  NAND2_X1 U149 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI222_X1 U150 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n155), .ZN(n208) );
  AOI22_X1 U151 ( .A1(C[25]), .A2(n149), .B1(A[25]), .B2(n143), .ZN(n209) );
  NAND2_X1 U152 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI222_X1 U153 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n155), .ZN(n216) );
  AOI22_X1 U154 ( .A1(C[29]), .A2(n149), .B1(A[29]), .B2(n143), .ZN(n217) );
  NAND2_X1 U155 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI222_X1 U156 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n156), .ZN(n226) );
  AOI22_X1 U157 ( .A1(C[33]), .A2(n149), .B1(A[33]), .B2(n143), .ZN(n227) );
  NAND2_X1 U158 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI222_X1 U159 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n156), .ZN(n234) );
  AOI22_X1 U160 ( .A1(C[37]), .A2(n148), .B1(A[37]), .B2(n142), .ZN(n235) );
  NAND2_X1 U161 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI22_X1 U162 ( .A1(C[17]), .A2(n150), .B1(A[17]), .B2(n144), .ZN(n191) );
  AOI222_X1 U163 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n154), .ZN(n190) );
  AOI22_X1 U164 ( .A1(C[32]), .A2(n149), .B1(A[32]), .B2(n143), .ZN(n225) );
  AOI222_X1 U165 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n156), .ZN(n224) );
  AOI222_X1 U166 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n156), .ZN(n242) );
  AOI22_X1 U167 ( .A1(C[40]), .A2(n148), .B1(A[40]), .B2(n142), .ZN(n243) );
  NAND2_X1 U168 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI22_X1 U169 ( .A1(C[39]), .A2(n148), .B1(A[39]), .B2(n142), .ZN(n239) );
  AOI222_X1 U170 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n156), .ZN(n238) );
  AOI22_X1 U171 ( .A1(C[36]), .A2(n148), .B1(A[36]), .B2(n142), .ZN(n233) );
  AOI222_X1 U172 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n156), .ZN(n232) );
  NAND2_X1 U173 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  AOI22_X1 U174 ( .A1(C[56]), .A2(n147), .B1(A[56]), .B2(n141), .ZN(n277) );
  AOI222_X1 U175 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n158), .ZN(n276) );
  NAND2_X1 U176 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  AOI22_X1 U177 ( .A1(C[57]), .A2(n146), .B1(A[57]), .B2(n140), .ZN(n279) );
  AOI222_X1 U178 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n158), .ZN(n278) );
  NAND2_X1 U179 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI22_X1 U180 ( .A1(C[58]), .A2(n146), .B1(A[58]), .B2(n140), .ZN(n281) );
  AOI222_X1 U181 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n158), .ZN(n280) );
  NAND2_X1 U182 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U183 ( .A1(C[59]), .A2(n146), .B1(A[59]), .B2(n140), .ZN(n283) );
  AOI222_X1 U184 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n158), .ZN(n282) );
  NAND2_X1 U185 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U186 ( .A1(C[60]), .A2(n146), .B1(A[60]), .B2(n140), .ZN(n287) );
  AOI222_X1 U187 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n158), .ZN(n286) );
  NAND2_X1 U188 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U189 ( .A1(C[61]), .A2(n146), .B1(A[61]), .B2(n140), .ZN(n289) );
  AOI222_X1 U190 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n158), .ZN(n288) );
  NAND2_X1 U191 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U192 ( .A1(C[62]), .A2(n146), .B1(A[62]), .B2(n140), .ZN(n291) );
  AOI222_X1 U193 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n158), .ZN(n290) );
  NAND2_X1 U194 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U195 ( .A1(C[63]), .A2(n146), .B1(A[63]), .B2(n140), .ZN(n293) );
  AOI222_X1 U196 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n158), .ZN(n292) );
  NAND2_X1 U197 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U198 ( .A1(C[0]), .A2(n146), .B1(A[0]), .B2(n140), .ZN(n175) );
  AOI222_X1 U199 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n154), .ZN(n174) );
  NAND2_X1 U200 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U201 ( .A1(C[4]), .A2(n147), .B1(A[4]), .B2(n141), .ZN(n263) );
  AOI222_X1 U202 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n157), .ZN(n262) );
  NAND2_X1 U203 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U204 ( .A1(C[1]), .A2(n150), .B1(A[1]), .B2(n144), .ZN(n197) );
  AOI222_X1 U205 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n154), .ZN(n196) );
  NAND2_X1 U206 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U207 ( .A1(C[5]), .A2(n146), .B1(A[5]), .B2(n140), .ZN(n285) );
  AOI222_X1 U208 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n158), .ZN(n284) );
  NAND2_X1 U209 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U210 ( .A1(C[2]), .A2(n149), .B1(A[2]), .B2(n143), .ZN(n219) );
  AOI222_X1 U211 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n155), .ZN(n218) );
  NAND2_X1 U212 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U213 ( .A1(C[6]), .A2(n146), .B1(A[6]), .B2(n140), .ZN(n295) );
  AOI222_X1 U214 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n158), .ZN(n294) );
  NAND2_X1 U215 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U216 ( .A1(C[3]), .A2(n148), .B1(A[3]), .B2(n142), .ZN(n241) );
  AOI222_X1 U217 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n156), .ZN(n240) );
  NAND2_X1 U218 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U219 ( .A1(C[7]), .A2(n146), .B1(A[7]), .B2(n140), .ZN(n297) );
  AOI222_X1 U220 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n158), .ZN(n296) );
  AOI22_X1 U221 ( .A1(C[8]), .A2(n146), .B1(A[8]), .B2(n140), .ZN(n299) );
  NAND2_X1 U222 ( .A1(n305), .A2(n304), .ZN(Y[9]) );
  AOI22_X1 U223 ( .A1(C[9]), .A2(n148), .B1(A[9]), .B2(n142), .ZN(n305) );
  AOI222_X1 U224 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n154), .ZN(n176) );
  NAND2_X1 U225 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI222_X1 U226 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n154), .ZN(n182) );
  AOI222_X1 U227 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n158), .ZN(n304) );
  AOI222_X1 U228 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n154), .ZN(n178) );
  CLKBUF_X1 U229 ( .A(n300), .Z(n145) );
  CLKBUF_X1 U230 ( .A(n301), .Z(n151) );
  CLKBUF_X1 U231 ( .A(n139), .Z(n164) );
endmodule


module G_204 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_756 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_755 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_754 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_753 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_752 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_751 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_750 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_749 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_748 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_747 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_746 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3, n5;

  CLKBUF_X1 U1 ( .A(P_IK), .Z(n3) );
  AND2_X1 U2 ( .A1(n3), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n5) );
  INV_X1 U4 ( .A(n5), .ZN(Gx) );
endmodule


module PG_745 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_744 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_743 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_742 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_741 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_740 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_739 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_738 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_737 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_736 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_735 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_734 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_733 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_732 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_731 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_730 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_729 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_728 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_727 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_726 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_203 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_725 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_724 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_723 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_722 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_721 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_720 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_719 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_718 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_717 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_716 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_715 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_714 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_713 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_712 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_711 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_202 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_710 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_709 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_708 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_707 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_706 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_705 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_704 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_201 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_200 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_703 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_702 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_701 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3;

  OR2_X1 U1 ( .A1(n3), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_700 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_699 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_698 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_199 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_198 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_197 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module G_196 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_697 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_696 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_695 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_694 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module G_195 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_194 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_193 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_192 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_191 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_190 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_189 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_188 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module carry_generator_N64_NPB4_12 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U77 ( .A(B[59]), .B(A[59]), .Z(\PG_Network[0][0][59] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U81 ( .A(B[55]), .B(A[55]), .Z(\PG_Network[0][0][55] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U85 ( .A(B[51]), .B(A[51]), .Z(\PG_Network[0][0][51] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U88 ( .A(B[49]), .B(A[49]), .Z(\PG_Network[0][0][49] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U90 ( .A(B[47]), .B(A[47]), .Z(\PG_Network[0][0][47] ) );
  XOR2_X1 U91 ( .A(B[46]), .B(A[46]), .Z(\PG_Network[0][0][46] ) );
  XOR2_X1 U92 ( .A(B[45]), .B(A[45]), .Z(\PG_Network[0][0][45] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U100 ( .A(B[38]), .B(A[38]), .Z(\PG_Network[0][0][38] ) );
  XOR2_X1 U101 ( .A(B[37]), .B(A[37]), .Z(\PG_Network[0][0][37] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U110 ( .A(B[29]), .B(A[29]), .Z(\PG_Network[0][0][29] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_204 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n23), .Gx(\PG_Network[1][1][1] ) );
  PG_756 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_755 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_754 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_753 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_752 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_751 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_750 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_749 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_748 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_747 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_746 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_745 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_744 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_743 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_742 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_741 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_740 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_739 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_738 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_737 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_736 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_735 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_734 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_733 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_732 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_731 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_730 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_729 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_728 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_727 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_726 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_203 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_725 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_724 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_723 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_722 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_721 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_720 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_719 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_718 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_717 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_716 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_715 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_714 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_713 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_712 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_711 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_202 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_710 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_709 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_708 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_707 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_706 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_705 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_704 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_201 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), .G_K_1(Co[1]), .Gx(Co[3]) );
  G_200 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_703 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(n5), .P_K_1(\PG_Network[3][0][23] ), 
        .Gx(\PG_Network[4][1][31] ), .Px(\PG_Network[4][0][31] ) );
  PG_702 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_701 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(n8), .P_K_1(n9), .Gx(
        \PG_Network[4][1][47] ), .Px(\PG_Network[4][0][47] ) );
  PG_700 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(n19), .P_K_1(n9), .Gx(
        \PG_Network[4][1][43] ), .Px(\PG_Network[4][0][43] ) );
  PG_699 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][63] ), .Px(
        \PG_Network[4][0][63] ) );
  PG_698 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][59] ), .Px(
        \PG_Network[4][0][59] ) );
  G_199 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), .G_K_1(n6), .Gx(Co[7]) );
  G_198 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), .G_K_1(n6), .Gx(Co[6]) );
  G_197 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), .G_K_1(n6), .Gx(Co[5]) );
  G_196 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), .G_K_1(Co[3]), .Gx(Co[4]) );
  PG_697 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][63] ), .Px(
        \PG_Network[5][0][63] ) );
  PG_696 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][59] ), .Px(
        \PG_Network[5][0][59] ) );
  PG_695 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][55] ), .Px(
        \PG_Network[5][0][55] ) );
  PG_694 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][51] ), .Px(
        \PG_Network[5][0][51] ) );
  G_195 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), .G_K_1(n21), .Gx(Co[15]) );
  G_194 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), .G_K_1(n21), .Gx(Co[14]) );
  G_193 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), .G_K_1(n21), .Gx(Co[13]) );
  G_192 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), .G_K_1(n21), .Gx(Co[12]) );
  G_191 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), .G_K_1(n21), .Gx(Co[11]) );
  G_190 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), .G_K_1(n21), .Gx(Co[10]) );
  G_189 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), .G_K_1(n7), .Gx(Co[9]) );
  G_188 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), .G_K_1(Co[7]), .Gx(Co[8]) );
  CLKBUF_X1 U1 ( .A(\PG_Network[3][1][23] ), .Z(n5) );
  INV_X1 U2 ( .A(A[43]), .ZN(n11) );
  INV_X1 U3 ( .A(A[35]), .ZN(n14) );
  INV_X1 U4 ( .A(A[11]), .ZN(n15) );
  INV_X1 U5 ( .A(A[15]), .ZN(n20) );
  INV_X1 U6 ( .A(A[23]), .ZN(n18) );
  INV_X1 U7 ( .A(A[27]), .ZN(n16) );
  INV_X1 U8 ( .A(A[31]), .ZN(n17) );
  INV_X1 U9 ( .A(A[30]), .ZN(n13) );
  INV_X1 U10 ( .A(A[19]), .ZN(n12) );
  INV_X1 U11 ( .A(A[39]), .ZN(n22) );
  INV_X1 U12 ( .A(A[25]), .ZN(n10) );
  CLKBUF_X1 U13 ( .A(Co[3]), .Z(n6) );
  CLKBUF_X1 U14 ( .A(Co[7]), .Z(n7) );
  CLKBUF_X1 U15 ( .A(n19), .Z(n8) );
  CLKBUF_X1 U16 ( .A(\PG_Network[3][0][39] ), .Z(n9) );
  CLKBUF_X1 U17 ( .A(n7), .Z(n21) );
  XNOR2_X1 U18 ( .A(B[25]), .B(n10), .ZN(\PG_Network[0][0][25] ) );
  XNOR2_X1 U19 ( .A(B[43]), .B(n11), .ZN(\PG_Network[0][0][43] ) );
  XNOR2_X1 U20 ( .A(B[19]), .B(n12), .ZN(\PG_Network[0][0][19] ) );
  XNOR2_X1 U21 ( .A(B[30]), .B(n13), .ZN(\PG_Network[0][0][30] ) );
  XNOR2_X1 U22 ( .A(B[35]), .B(n14), .ZN(\PG_Network[0][0][35] ) );
  XNOR2_X1 U23 ( .A(B[11]), .B(n15), .ZN(\PG_Network[0][0][11] ) );
  XNOR2_X1 U24 ( .A(B[27]), .B(n16), .ZN(\PG_Network[0][0][27] ) );
  XNOR2_X1 U25 ( .A(B[31]), .B(n17), .ZN(\PG_Network[0][0][31] ) );
  XNOR2_X1 U26 ( .A(B[23]), .B(n18), .ZN(\PG_Network[0][0][23] ) );
  BUF_X1 U27 ( .A(\PG_Network[3][1][39] ), .Z(n19) );
  XNOR2_X1 U28 ( .A(B[15]), .B(n20), .ZN(\PG_Network[0][0][15] ) );
  XNOR2_X1 U29 ( .A(B[39]), .B(n22), .ZN(\PG_Network[0][0][39] ) );
  AND2_X1 U30 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U31 ( .A1(B[30]), .A2(A[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U32 ( .A1(B[31]), .A2(A[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U33 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U34 ( .A1(A[35]), .A2(B[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U35 ( .A1(A[46]), .A2(B[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U36 ( .A1(A[47]), .A2(B[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U37 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U38 ( .A1(B[15]), .A2(A[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U39 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U40 ( .A1(A[37]), .A2(B[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U41 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U42 ( .A1(B[11]), .A2(A[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U43 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U44 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U45 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AND2_X1 U46 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U47 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U48 ( .A1(B[19]), .A2(A[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U49 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U50 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U51 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U52 ( .A1(B[25]), .A2(A[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U53 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U54 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U55 ( .A1(A[45]), .A2(B[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U56 ( .A1(A[49]), .A2(B[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U57 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U58 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U59 ( .A1(A[51]), .A2(B[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U60 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U61 ( .A1(A[55]), .A2(B[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U62 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U63 ( .A1(A[43]), .A2(B[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U64 ( .A1(A[41]), .A2(B[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U65 ( .A1(A[29]), .A2(B[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U66 ( .A1(A[53]), .A2(B[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U67 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U94 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U99 ( .A1(B[21]), .A2(A[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U103 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AND2_X1 U107 ( .A1(B[23]), .A2(A[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U108 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U112 ( .A1(A[59]), .A2(B[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U114 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
  AND2_X1 U116 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U121 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U125 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U129 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U131 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U132 ( .A(n26), .ZN(n23) );
  AND2_X1 U133 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U134 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U135 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U136 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U137 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U138 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U139 ( .A1(A[7]), .A2(B[7]), .ZN(\PG_Network[0][1][7] ) );
  AOI21_X1 U140 ( .B1(A[0]), .B2(B[0]), .A(n24), .ZN(n26) );
  INV_X1 U141 ( .A(n25), .ZN(n24) );
  OAI21_X1 U142 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n25) );
  AND2_X1 U143 ( .A1(B[27]), .A2(A[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U144 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U145 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U146 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U147 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U148 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
endmodule


module FA_1536 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1535 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1534 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1533 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_384 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1536 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1535 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1534 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1533 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1532 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1531 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1530 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1529 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_383 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1532 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1531 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1530 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1529 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_192 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U2 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_192 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_384 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_383 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_192 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1528 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1527 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1526 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1525 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_382 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1528 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1527 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1526 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1525 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1524 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1523 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1522 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1521 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_381 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1524 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1523 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1522 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1521 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_191 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_191 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_382 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_381 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_191 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1520 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1519 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1518 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1517 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_380 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1520 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1519 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1518 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1517 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1516 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1515 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1514 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1513 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_379 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1516 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1515 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1514 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1513 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_190 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U2 ( .A(sel), .ZN(n13) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_190 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_380 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_379 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_190 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1512 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8, n9;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n5) );
  CLKBUF_X1 U2 ( .A(n9), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n7), .A2(n8), .ZN(Co) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(n7) );
  NAND2_X1 U7 ( .A1(n9), .A2(Ci), .ZN(n8) );
endmodule


module FA_1511 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1510 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1509 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_378 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1512 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1511 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1510 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1509 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1508 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1507 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1506 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1505 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_377 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1508 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1507 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1506 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1505 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_189 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n18), .ZN(Y[2]) );
  BUF_X1 U2 ( .A(sel), .Z(n5) );
  INV_X1 U3 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U4 ( .A(sel), .ZN(n10) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U6 ( .A(sel), .ZN(n15) );
  INV_X1 U7 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n10), .ZN(n19) );
  AOI22_X1 U10 ( .A1(n5), .A2(A[1]), .B1(B[1]), .B2(n10), .ZN(n17) );
  AOI22_X1 U11 ( .A1(A[0]), .A2(sel), .B1(n15), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_189 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_378 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_377 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_189 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1504 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n5) );
  AOI22_X1 U5 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_1503 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1502 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1501 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_376 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1504 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1503 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1502 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1501 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1500 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1499 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1498 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1497 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_375 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1500 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1499 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1498 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1497 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_188 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U3 ( .A(sel), .ZN(n5) );
  INV_X1 U4 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U6 ( .A(sel), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n14), .ZN(n17) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n5), .ZN(n15) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n14), .ZN(n18) );
endmodule


module carry_select_block_NPB4_188 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_376 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_375 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_188 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1496 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_1495 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1494 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1493 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  OR2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_374 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1496 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1495 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1494 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1493 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1492 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1491 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1490 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1489 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_373 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1492 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1491 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1490 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1489 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_187 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  CLKBUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U5 ( .A(sel), .ZN(n10) );
  INV_X1 U6 ( .A(sel), .ZN(n15) );
  AOI22_X1 U7 ( .A1(n5), .A2(A[2]), .B1(n10), .B2(B[2]), .ZN(n18) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[1]), .B1(n10), .B2(B[1]), .ZN(n17) );
  INV_X1 U9 ( .A(n16), .ZN(Y[0]) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(sel), .B1(n10), .B2(B[3]), .ZN(n19) );
endmodule


module carry_select_block_NPB4_187 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_374 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_373 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_187 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1488 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_1487 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1486 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1485 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  OR2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n7) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(n4), .ZN(n10) );
endmodule


module RCA_N4_372 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1488 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1487 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1486 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1485 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1484 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1483 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(n4), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1482 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1481 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_371 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1484 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1483 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1482 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1481 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_186 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U5 ( .A(sel), .ZN(n10) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(n5), .A2(A[2]), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[1]), .B1(n10), .B2(B[1]), .ZN(n17) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n10), .ZN(n19) );
endmodule


module carry_select_block_NPB4_186 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_372 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_371 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_186 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1480 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1479 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1478 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1477 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_370 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1480 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1479 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1478 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1477 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1476 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1475 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1474 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1473 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_369 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1476 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1475 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1474 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1473 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_185 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(sel), .Z(n10) );
  INV_X1 U2 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n10), .ZN(n5) );
  INV_X1 U4 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U7 ( .A1(n10), .A2(A[1]), .B1(B[1]), .B2(n15), .ZN(n17) );
  INV_X1 U8 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_185 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_370 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_369 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_185 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1472 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_1471 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1470 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1469 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_368 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1472 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1471 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1470 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1469 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1468 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1467 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1466 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1465 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_367 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1468 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1467 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1466 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1465 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_184 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n15), .ZN(Y[0]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n5) );
  INV_X1 U3 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U5 ( .A(n16), .ZN(Y[1]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n14), .ZN(n17) );
  AOI22_X1 U7 ( .A1(n5), .A2(A[1]), .B1(B[1]), .B2(n14), .ZN(n16) );
  INV_X1 U8 ( .A(sel), .ZN(n14) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n14), .ZN(n18) );
endmodule


module carry_select_block_NPB4_184 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_368 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_367 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_184 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1464 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(n4), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1463 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1462 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1461 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_366 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1464 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1463 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1462 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1461 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1460 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1459 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1458 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1457 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_365 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1460 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1459 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1458 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1457 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_183 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n16), .ZN(Y[0]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(n10), .ZN(n5) );
  INV_X1 U4 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(n15), .B2(B[1]), .ZN(n17) );
  INV_X1 U8 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_183 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_366 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_365 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_183 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1456 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6, n7, n8;

  XOR2_X1 U3 ( .A(n8), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n8) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U6 ( .A1(n8), .A2(Ci), .ZN(n7) );
endmodule


module FA_1455 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1454 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1453 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_364 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1456 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1455 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1454 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1453 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1452 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1451 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1450 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1449 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_363 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1452 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1451 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1450 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1449 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_182 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X2 U1 ( .A(n17), .ZN(Y[1]) );
  BUF_X2 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(n10), .ZN(n5) );
  INV_X1 U4 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U8 ( .A1(n10), .A2(A[1]), .B1(B[1]), .B2(n5), .ZN(n17) );
  INV_X1 U9 ( .A(sel), .ZN(n15) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U11 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
endmodule


module carry_select_block_NPB4_182 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_364 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_363 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_182 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1448 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1447 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1446 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1445 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_362 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1448 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1447 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1446 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1445 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1444 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1443 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1442 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1441 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_361 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1444 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1443 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1442 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1441 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_181 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n10), .ZN(n5) );
  BUF_X2 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U4 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(n10), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(n10), .B1(n15), .B2(B[1]), .ZN(n17) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_181 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_362 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_361 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_181 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1440 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1439 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1438 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1437 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_360 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1440 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1439 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1438 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1437 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1436 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1435 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1434 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1433 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_359 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1436 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1435 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1434 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1433 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_180 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n15), .ZN(Y[0]) );
  CLKBUF_X1 U2 ( .A(n14), .Z(n5) );
  INV_X1 U3 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U4 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n18) );
  INV_X1 U5 ( .A(n17), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n17) );
  INV_X1 U7 ( .A(n16), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n5), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
  INV_X1 U10 ( .A(sel), .ZN(n14) );
endmodule


module carry_select_block_NPB4_180 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_360 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_359 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_180 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1432 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1431 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1430 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1429 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_358 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1432 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1431 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1430 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1429 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1428 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1427 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1426 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1425 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_357 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1428 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1427 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1426 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1425 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_179 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_179 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_358 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_357 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_179 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1424 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1423 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1422 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1421 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_356 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1424 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1423 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1422 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1421 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1420 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1419 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1418 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1417 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_355 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1420 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1419 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1418 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1417 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_178 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_178 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_356 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_355 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_178 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1416 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1415 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1414 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1413 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_354 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1416 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1415 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1414 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1413 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1412 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1411 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1410 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1409 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_353 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1412 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1411 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1410 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1409 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_177 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_177 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_354 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_353 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_177 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_12 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_192 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_191 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_190 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_189 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_188 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_187 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_186 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_185 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_184 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_183 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_182 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), .S(S[43:40]) );
  carry_select_block_NPB4_181 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), .S(S[47:44]) );
  carry_select_block_NPB4_180 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), .S(S[51:48]) );
  carry_select_block_NPB4_179 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), .S(S[55:52]) );
  carry_select_block_NPB4_178 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), .S(S[59:56]) );
  carry_select_block_NPB4_177 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), .S(S[63:60]) );
endmodule


module P4_ADDER_N64_12 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_12 CGEN ( .A(A), .B({B[63:29], n23, B[27:25], n7, 
        B[23:21], n22, B[19:17], n21, B[15:13], n15, B[11:0]}), .Cin(Cin), 
        .Co(CoutCgen) );
  sum_generator_N64_NPB4_12 SGEN ( .A(A), .B({B[63:44], n10, B[42:40], n17, 
        B[38:36], n12, B[34:32], n1, n14, B[29:28], n9, n3, B[25:24], n20, n5, 
        B[21:20], n6, n11, B[17:16], n19, B[14:12], n13, B[10:0]}), .Ci({
        CoutCgen, Cin}), .S(S), .Co(Cout) );
  BUF_X1 U1 ( .A(B[18]), .Z(n11) );
  BUF_X1 U2 ( .A(B[30]), .Z(n14) );
  CLKBUF_X1 U3 ( .A(B[31]), .Z(n1) );
  INV_X1 U4 ( .A(B[26]), .ZN(n2) );
  INV_X1 U5 ( .A(n2), .ZN(n3) );
  CLKBUF_X1 U6 ( .A(B[39]), .Z(n4) );
  CLKBUF_X1 U7 ( .A(B[22]), .Z(n5) );
  CLKBUF_X1 U8 ( .A(B[19]), .Z(n6) );
  CLKBUF_X1 U9 ( .A(B[24]), .Z(n7) );
  INV_X1 U10 ( .A(B[27]), .ZN(n8) );
  INV_X1 U11 ( .A(n8), .ZN(n9) );
  CLKBUF_X1 U12 ( .A(B[11]), .Z(n13) );
  BUF_X1 U13 ( .A(B[28]), .Z(n23) );
  CLKBUF_X1 U14 ( .A(B[43]), .Z(n10) );
  CLKBUF_X1 U15 ( .A(B[35]), .Z(n12) );
  CLKBUF_X1 U16 ( .A(B[12]), .Z(n15) );
  INV_X1 U17 ( .A(n4), .ZN(n16) );
  INV_X1 U18 ( .A(n16), .ZN(n17) );
  INV_X1 U19 ( .A(B[15]), .ZN(n18) );
  INV_X1 U20 ( .A(n18), .ZN(n19) );
  CLKBUF_X1 U21 ( .A(B[23]), .Z(n20) );
  CLKBUF_X1 U22 ( .A(B[16]), .Z(n21) );
  CLKBUF_X1 U23 ( .A(B[20]), .Z(n22) );
endmodule


module Booth_Encoder_11 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_11 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305;

  NAND2_X1 U1 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  NAND2_X1 U2 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  NAND2_X2 U3 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  NAND2_X1 U4 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  NAND2_X1 U5 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  NOR3_X1 U6 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U7 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  NAND2_X1 U8 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  NAND2_X2 U9 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  NOR4_X1 U10 ( .A1(n151), .A2(n145), .A3(n154), .A4(n167), .ZN(n139) );
  BUF_X1 U11 ( .A(n139), .Z(n161) );
  BUF_X1 U12 ( .A(n139), .Z(n160) );
  BUF_X1 U13 ( .A(n139), .Z(n159) );
  BUF_X1 U14 ( .A(n139), .Z(n162) );
  BUF_X1 U15 ( .A(n139), .Z(n163) );
  BUF_X1 U16 ( .A(n152), .Z(n155) );
  BUF_X1 U17 ( .A(n152), .Z(n156) );
  BUF_X1 U18 ( .A(n165), .Z(n168) );
  BUF_X1 U19 ( .A(n152), .Z(n154) );
  BUF_X1 U20 ( .A(n165), .Z(n167) );
  BUF_X1 U21 ( .A(n153), .Z(n157) );
  BUF_X1 U22 ( .A(n165), .Z(n169) );
  BUF_X1 U23 ( .A(n166), .Z(n170) );
  BUF_X1 U24 ( .A(n153), .Z(n158) );
  BUF_X1 U25 ( .A(n166), .Z(n171) );
  CLKBUF_X1 U26 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U27 ( .A(n301), .Z(n149) );
  BUF_X1 U28 ( .A(n303), .Z(n165) );
  BUF_X1 U29 ( .A(n302), .Z(n152) );
  CLKBUF_X1 U30 ( .A(n301), .Z(n147) );
  CLKBUF_X1 U31 ( .A(n301), .Z(n148) );
  BUF_X1 U32 ( .A(n303), .Z(n166) );
  BUF_X1 U33 ( .A(n302), .Z(n153) );
  CLKBUF_X1 U34 ( .A(n301), .Z(n146) );
  BUF_X1 U35 ( .A(n300), .Z(n140) );
  BUF_X1 U36 ( .A(n300), .Z(n144) );
  BUF_X1 U37 ( .A(n300), .Z(n141) );
  BUF_X1 U38 ( .A(n300), .Z(n143) );
  BUF_X1 U39 ( .A(n300), .Z(n142) );
  INV_X1 U40 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U41 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n303) );
  AND3_X1 U42 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U43 ( .A(sel[2]), .ZN(n173) );
  AOI22_X1 U44 ( .A1(C[24]), .A2(n150), .B1(A[24]), .B2(n144), .ZN(n207) );
  AOI222_X1 U45 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n155), .ZN(n206) );
  NAND2_X1 U46 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI22_X1 U47 ( .A1(C[25]), .A2(n149), .B1(A[25]), .B2(n143), .ZN(n209) );
  AOI222_X1 U48 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n155), .ZN(n208) );
  NAND2_X1 U49 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI222_X1 U50 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n156), .ZN(n228) );
  AOI22_X1 U51 ( .A1(C[34]), .A2(n149), .B1(A[34]), .B2(n143), .ZN(n229) );
  NAND2_X1 U52 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U53 ( .A1(C[13]), .A2(n151), .B1(A[13]), .B2(n145), .ZN(n183) );
  NAND2_X1 U54 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U55 ( .A1(C[15]), .A2(n150), .B1(A[15]), .B2(n144), .ZN(n187) );
  NAND2_X1 U56 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  AOI22_X1 U57 ( .A1(C[48]), .A2(n147), .B1(A[48]), .B2(n141), .ZN(n259) );
  AOI222_X1 U58 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n157), .ZN(n258) );
  NAND2_X1 U59 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  AOI22_X1 U60 ( .A1(C[52]), .A2(n147), .B1(A[52]), .B2(n141), .ZN(n269) );
  AOI222_X1 U61 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n157), .ZN(n268) );
  NAND2_X1 U62 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI22_X1 U63 ( .A1(C[45]), .A2(n148), .B1(A[45]), .B2(n142), .ZN(n253) );
  AOI222_X1 U64 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n157), .ZN(n252) );
  NAND2_X1 U65 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI22_X1 U66 ( .A1(C[49]), .A2(n147), .B1(A[49]), .B2(n141), .ZN(n261) );
  AOI222_X1 U67 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n157), .ZN(n260) );
  NAND2_X1 U68 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI22_X1 U69 ( .A1(C[50]), .A2(n147), .B1(A[50]), .B2(n141), .ZN(n265) );
  AOI222_X1 U70 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n157), .ZN(n264) );
  NAND2_X1 U71 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI22_X1 U72 ( .A1(C[47]), .A2(n147), .B1(A[47]), .B2(n141), .ZN(n257) );
  AOI222_X1 U73 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n157), .ZN(n256) );
  NAND2_X1 U74 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  AOI22_X1 U75 ( .A1(C[51]), .A2(n147), .B1(A[51]), .B2(n141), .ZN(n267) );
  AOI222_X1 U76 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n157), .ZN(n266) );
  AOI22_X1 U77 ( .A1(C[16]), .A2(n150), .B1(A[16]), .B2(n144), .ZN(n189) );
  AOI222_X1 U78 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n154), .ZN(n188) );
  NAND2_X1 U79 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI22_X1 U80 ( .A1(C[17]), .A2(n150), .B1(A[17]), .B2(n144), .ZN(n191) );
  AOI222_X1 U81 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n154), .ZN(n190) );
  AOI22_X1 U82 ( .A1(C[29]), .A2(n149), .B1(A[29]), .B2(n143), .ZN(n217) );
  AOI222_X1 U83 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n155), .ZN(n216) );
  NAND2_X1 U84 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI22_X1 U85 ( .A1(C[18]), .A2(n150), .B1(A[18]), .B2(n144), .ZN(n193) );
  AOI222_X1 U86 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n154), .ZN(n192) );
  NAND2_X1 U87 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI22_X1 U88 ( .A1(C[26]), .A2(n149), .B1(A[26]), .B2(n143), .ZN(n211) );
  AOI222_X1 U89 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n155), .ZN(n210) );
  NAND2_X1 U90 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI222_X1 U91 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n155), .ZN(n212) );
  AOI22_X1 U92 ( .A1(C[27]), .A2(n149), .B1(A[27]), .B2(n143), .ZN(n213) );
  NAND2_X1 U93 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI222_X1 U94 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n155), .ZN(n204) );
  AOI22_X1 U95 ( .A1(C[23]), .A2(n150), .B1(A[23]), .B2(n144), .ZN(n205) );
  NAND2_X1 U96 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI222_X1 U97 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n156), .ZN(n230) );
  AOI22_X1 U98 ( .A1(C[35]), .A2(n149), .B1(A[35]), .B2(n143), .ZN(n231) );
  NAND2_X1 U99 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI22_X1 U100 ( .A1(C[19]), .A2(n150), .B1(A[19]), .B2(n144), .ZN(n195) );
  AOI222_X1 U101 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n154), .ZN(n194) );
  NAND2_X1 U102 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U103 ( .A1(C[14]), .A2(n150), .B1(A[14]), .B2(n144), .ZN(n185) );
  AOI222_X1 U104 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n154), .ZN(n184) );
  NAND2_X1 U105 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI222_X1 U106 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n156), .ZN(n234) );
  NAND2_X1 U107 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI222_X1 U108 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n156), .ZN(n226) );
  NAND2_X1 U109 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI222_X1 U110 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n156), .ZN(n244) );
  NAND2_X1 U111 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI222_X1 U112 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n156), .ZN(n246) );
  AOI22_X1 U113 ( .A1(C[42]), .A2(n148), .B1(A[42]), .B2(n142), .ZN(n247) );
  NAND2_X1 U114 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI22_X1 U115 ( .A1(C[46]), .A2(n147), .B1(A[46]), .B2(n141), .ZN(n255) );
  AOI222_X1 U116 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n157), .ZN(n254) );
  NAND2_X1 U117 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  AOI22_X1 U118 ( .A1(C[28]), .A2(n149), .B1(A[28]), .B2(n143), .ZN(n215) );
  AOI222_X1 U119 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n155), .ZN(n214) );
  NAND2_X1 U120 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  AOI22_X1 U121 ( .A1(C[32]), .A2(n149), .B1(A[32]), .B2(n143), .ZN(n225) );
  AOI222_X1 U122 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n156), .ZN(n224) );
  AOI22_X1 U123 ( .A1(C[20]), .A2(n150), .B1(A[20]), .B2(n144), .ZN(n199) );
  AOI222_X1 U124 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n155), .ZN(n198) );
  AOI222_X1 U125 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n156), .ZN(n236) );
  NAND2_X1 U126 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI22_X1 U127 ( .A1(C[21]), .A2(n150), .B1(A[21]), .B2(n144), .ZN(n201) );
  AOI222_X1 U128 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n155), .ZN(n200) );
  NAND2_X1 U129 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI22_X1 U130 ( .A1(C[22]), .A2(n150), .B1(A[22]), .B2(n144), .ZN(n203) );
  AOI222_X1 U131 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n155), .ZN(n202) );
  NAND2_X1 U132 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U133 ( .A1(C[30]), .A2(n149), .B1(A[30]), .B2(n143), .ZN(n221) );
  AOI222_X1 U134 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n155), .ZN(n220) );
  AOI22_X1 U135 ( .A1(C[12]), .A2(n151), .B1(A[12]), .B2(n145), .ZN(n181) );
  NAND2_X1 U136 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  AOI22_X1 U137 ( .A1(C[44]), .A2(n148), .B1(A[44]), .B2(n142), .ZN(n251) );
  AOI222_X1 U138 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n157), .ZN(n250) );
  NAND2_X1 U139 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI22_X1 U140 ( .A1(C[43]), .A2(n148), .B1(A[43]), .B2(n142), .ZN(n249) );
  AOI222_X1 U141 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n156), .ZN(n248) );
  NAND2_X1 U142 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  AOI22_X1 U143 ( .A1(C[36]), .A2(n148), .B1(A[36]), .B2(n142), .ZN(n233) );
  AOI222_X1 U144 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n156), .ZN(n232) );
  AOI22_X1 U145 ( .A1(C[40]), .A2(n148), .B1(A[40]), .B2(n142), .ZN(n243) );
  AOI222_X1 U146 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n156), .ZN(n242) );
  NAND2_X1 U147 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI222_X1 U148 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n156), .ZN(n238) );
  AOI22_X1 U149 ( .A1(C[39]), .A2(n148), .B1(A[39]), .B2(n142), .ZN(n239) );
  NAND2_X1 U150 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI222_X1 U151 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n155), .ZN(n222) );
  AOI22_X1 U152 ( .A1(C[31]), .A2(n149), .B1(A[31]), .B2(n143), .ZN(n223) );
  NAND2_X1 U153 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  AOI22_X1 U154 ( .A1(C[56]), .A2(n147), .B1(A[56]), .B2(n141), .ZN(n277) );
  AOI222_X1 U155 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n158), .ZN(n276) );
  NAND2_X1 U156 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  AOI22_X1 U157 ( .A1(C[53]), .A2(n147), .B1(A[53]), .B2(n141), .ZN(n271) );
  AOI222_X1 U158 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n157), .ZN(n270) );
  NAND2_X1 U159 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  AOI22_X1 U160 ( .A1(C[57]), .A2(n146), .B1(A[57]), .B2(n140), .ZN(n279) );
  AOI222_X1 U161 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n158), .ZN(n278) );
  NAND2_X1 U162 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI22_X1 U163 ( .A1(C[54]), .A2(n147), .B1(A[54]), .B2(n141), .ZN(n273) );
  AOI222_X1 U164 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n157), .ZN(n272) );
  NAND2_X1 U165 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI22_X1 U166 ( .A1(C[58]), .A2(n146), .B1(A[58]), .B2(n140), .ZN(n281) );
  AOI222_X1 U167 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n158), .ZN(n280) );
  NAND2_X1 U168 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI22_X1 U169 ( .A1(C[55]), .A2(n147), .B1(A[55]), .B2(n141), .ZN(n275) );
  AOI222_X1 U170 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n157), .ZN(n274) );
  NAND2_X1 U171 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U172 ( .A1(C[59]), .A2(n146), .B1(A[59]), .B2(n140), .ZN(n283) );
  AOI222_X1 U173 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n158), .ZN(n282) );
  NAND2_X1 U174 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U175 ( .A1(C[60]), .A2(n146), .B1(A[60]), .B2(n140), .ZN(n287) );
  AOI222_X1 U176 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n158), .ZN(n286) );
  NAND2_X1 U177 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U178 ( .A1(C[61]), .A2(n146), .B1(A[61]), .B2(n140), .ZN(n289) );
  AOI222_X1 U179 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n158), .ZN(n288) );
  NAND2_X1 U180 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U181 ( .A1(C[62]), .A2(n146), .B1(A[62]), .B2(n140), .ZN(n291) );
  AOI222_X1 U182 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n158), .ZN(n290) );
  NAND2_X1 U183 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U184 ( .A1(C[63]), .A2(n146), .B1(A[63]), .B2(n140), .ZN(n293) );
  AOI222_X1 U185 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n158), .ZN(n292) );
  NAND2_X1 U186 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U187 ( .A1(C[0]), .A2(n146), .B1(A[0]), .B2(n140), .ZN(n175) );
  AOI222_X1 U188 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n154), .ZN(n174) );
  NAND2_X1 U189 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U190 ( .A1(C[4]), .A2(n147), .B1(A[4]), .B2(n141), .ZN(n263) );
  AOI222_X1 U191 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n157), .ZN(n262) );
  NAND2_X1 U192 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI22_X1 U193 ( .A1(C[8]), .A2(n146), .B1(A[8]), .B2(n140), .ZN(n299) );
  AOI222_X1 U194 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n158), .ZN(n298) );
  NAND2_X1 U195 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U196 ( .A1(C[1]), .A2(n150), .B1(A[1]), .B2(n144), .ZN(n197) );
  AOI222_X1 U197 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n154), .ZN(n196) );
  NAND2_X1 U198 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U199 ( .A1(C[5]), .A2(n146), .B1(A[5]), .B2(n140), .ZN(n285) );
  AOI222_X1 U200 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n158), .ZN(n284) );
  NAND2_X1 U201 ( .A1(n305), .A2(n304), .ZN(Y[9]) );
  AOI22_X1 U202 ( .A1(C[9]), .A2(n148), .B1(A[9]), .B2(n142), .ZN(n305) );
  AOI222_X1 U203 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n158), .ZN(n304) );
  NAND2_X1 U204 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U205 ( .A1(C[2]), .A2(n149), .B1(A[2]), .B2(n143), .ZN(n219) );
  AOI222_X1 U206 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n155), .ZN(n218) );
  NAND2_X1 U207 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U208 ( .A1(C[6]), .A2(n146), .B1(A[6]), .B2(n140), .ZN(n295) );
  AOI222_X1 U209 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n158), .ZN(n294) );
  NAND2_X1 U210 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U211 ( .A1(C[3]), .A2(n148), .B1(A[3]), .B2(n142), .ZN(n241) );
  AOI222_X1 U212 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n156), .ZN(n240) );
  NAND2_X1 U213 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U214 ( .A1(C[7]), .A2(n146), .B1(A[7]), .B2(n140), .ZN(n297) );
  AOI222_X1 U215 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n158), .ZN(n296) );
  AOI22_X1 U216 ( .A1(C[38]), .A2(n148), .B1(A[38]), .B2(n142), .ZN(n237) );
  AOI22_X1 U217 ( .A1(C[37]), .A2(n148), .B1(A[37]), .B2(n142), .ZN(n235) );
  AOI22_X1 U218 ( .A1(C[10]), .A2(n151), .B1(A[10]), .B2(n145), .ZN(n177) );
  AOI222_X1 U219 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n154), .ZN(n176) );
  AOI22_X1 U220 ( .A1(C[11]), .A2(n151), .B1(A[11]), .B2(n145), .ZN(n179) );
  NAND2_X1 U221 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  NAND2_X1 U222 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI222_X1 U223 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n154), .ZN(n186) );
  AOI22_X1 U224 ( .A1(C[33]), .A2(n149), .B1(A[33]), .B2(n143), .ZN(n227) );
  AOI222_X1 U225 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n154), .ZN(n180) );
  AOI222_X1 U226 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n154), .ZN(n178) );
  AOI22_X1 U227 ( .A1(C[41]), .A2(n148), .B1(A[41]), .B2(n142), .ZN(n245) );
  AOI222_X1 U228 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n154), .ZN(n182) );
  CLKBUF_X1 U229 ( .A(n300), .Z(n145) );
  CLKBUF_X1 U230 ( .A(n301), .Z(n151) );
  CLKBUF_X1 U231 ( .A(n139), .Z(n164) );
endmodule


module G_187 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_693 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_692 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_691 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_690 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_689 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_688 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_687 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_686 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_685 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_684 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_683 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_682 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_681 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_680 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_679 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_678 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_677 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_676 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_675 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_674 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_673 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_672 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_671 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_670 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_669 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_668 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_667 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_666 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_665 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_664 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_663 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_186 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_662 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_661 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_660 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_659 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_658 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_657 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_656 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_655 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_654 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_653 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_652 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_651 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_650 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_649 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_648 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_185 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_647 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_646 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_645 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_644 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_643 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_642 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_641 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_184 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_183 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_640 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_639 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_638 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  OR2_X1 U2 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_637 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_636 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_635 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_182 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_181 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_180 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_179 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_634 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_633 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_632 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_631 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_178 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_177 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_176 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_175 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_174 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_173 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_172 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
endmodule


module G_171 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module carry_generator_N64_NPB4_11 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U77 ( .A(B[59]), .B(A[59]), .Z(\PG_Network[0][0][59] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U81 ( .A(B[55]), .B(A[55]), .Z(\PG_Network[0][0][55] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U85 ( .A(B[51]), .B(A[51]), .Z(\PG_Network[0][0][51] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U88 ( .A(B[49]), .B(A[49]), .Z(\PG_Network[0][0][49] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U91 ( .A(B[46]), .B(A[46]), .Z(\PG_Network[0][0][46] ) );
  XOR2_X1 U92 ( .A(B[45]), .B(A[45]), .Z(\PG_Network[0][0][45] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U108 ( .A(B[30]), .B(A[30]), .Z(\PG_Network[0][0][30] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U114 ( .A(B[25]), .B(A[25]), .Z(\PG_Network[0][0][25] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_187 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n31), .Gx(\PG_Network[1][1][1] ) );
  PG_693 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_692 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_691 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_690 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_689 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_688 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_687 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_686 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_685 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_684 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_683 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_682 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_681 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_680 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_679 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_678 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_677 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_676 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_675 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_674 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_673 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_672 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_671 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_670 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_669 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_668 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_667 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_666 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_665 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_664 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_663 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_186 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_662 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_661 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_660 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_659 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_658 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_657 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_656 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_655 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_654 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_653 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_652 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_651 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_650 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_649 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_648 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_185 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_647 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_646 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_645 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_644 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_643 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_642 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_641 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_184 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), .G_K_1(Co[1]), .Gx(Co[3]) );
  G_183 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_640 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_639 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_638 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(n30), 
        .Gx(\PG_Network[4][1][47] ), .Px(\PG_Network[4][0][47] ) );
  PG_637 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(n30), 
        .Gx(\PG_Network[4][1][43] ), .Px(\PG_Network[4][0][43] ) );
  PG_636 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][63] ), .Px(
        \PG_Network[4][0][63] ) );
  PG_635 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][59] ), .Px(
        \PG_Network[4][0][59] ) );
  G_182 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), .G_K_1(n17), .Gx(Co[7]) );
  G_181 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), .G_K_1(n17), .Gx(Co[6]) );
  G_180 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), .G_K_1(n21), .Gx(Co[5]) );
  G_179 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), .G_K_1(Co[3]), .Gx(Co[4]) );
  PG_634 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(n18), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][63] ), .Px(\PG_Network[5][0][63] ) );
  PG_633 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(n18), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][59] ), .Px(\PG_Network[5][0][59] ) );
  PG_632 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(n18), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][55] ), .Px(\PG_Network[5][0][55] ) );
  PG_631 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(n18), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][51] ), .Px(\PG_Network[5][0][51] ) );
  G_178 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), .G_K_1(n16), .Gx(Co[15]) );
  G_177 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), .G_K_1(n16), .Gx(Co[14]) );
  G_176 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), .G_K_1(n16), .Gx(Co[13]) );
  G_175 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), .G_K_1(n16), .Gx(Co[12]) );
  G_174 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), .G_K_1(n16), .Gx(Co[11]) );
  G_173 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), .G_K_1(n16), .Gx(Co[10]) );
  G_172 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), .G_K_1(n26), .Gx(Co[9]) );
  G_171 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), .G_K_1(Co[7]), .Gx(Co[8]) );
  INV_X1 U1 ( .A(A[20]), .ZN(n9) );
  BUF_X1 U2 ( .A(n26), .Z(n16) );
  NAND2_X1 U3 ( .A1(B[29]), .A2(n6), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n5), .A2(A[29]), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n7), .A2(n8), .ZN(\PG_Network[0][0][29] ) );
  INV_X1 U6 ( .A(B[29]), .ZN(n5) );
  INV_X1 U7 ( .A(A[29]), .ZN(n6) );
  XNOR2_X1 U8 ( .A(B[20]), .B(n9), .ZN(\PG_Network[0][0][20] ) );
  BUF_X1 U9 ( .A(Co[7]), .Z(n26) );
  NAND2_X1 U10 ( .A1(B[38]), .A2(n11), .ZN(n12) );
  NAND2_X1 U11 ( .A1(n10), .A2(A[38]), .ZN(n13) );
  NAND2_X1 U12 ( .A1(n12), .A2(n13), .ZN(\PG_Network[0][0][38] ) );
  INV_X1 U13 ( .A(B[38]), .ZN(n10) );
  INV_X1 U14 ( .A(A[38]), .ZN(n11) );
  INV_X1 U15 ( .A(A[15]), .ZN(n22) );
  INV_X1 U16 ( .A(A[47]), .ZN(n14) );
  INV_X1 U17 ( .A(A[35]), .ZN(n19) );
  INV_X1 U18 ( .A(A[37]), .ZN(n15) );
  INV_X1 U19 ( .A(A[27]), .ZN(n20) );
  INV_X1 U20 ( .A(A[23]), .ZN(n27) );
  INV_X1 U21 ( .A(A[19]), .ZN(n24) );
  INV_X1 U22 ( .A(A[21]), .ZN(n23) );
  INV_X1 U23 ( .A(A[43]), .ZN(n29) );
  INV_X1 U24 ( .A(A[39]), .ZN(n28) );
  INV_X1 U25 ( .A(A[31]), .ZN(n25) );
  XNOR2_X1 U26 ( .A(B[47]), .B(n14), .ZN(\PG_Network[0][0][47] ) );
  XNOR2_X1 U27 ( .A(B[37]), .B(n15), .ZN(\PG_Network[0][0][37] ) );
  BUF_X1 U28 ( .A(n21), .Z(n17) );
  CLKBUF_X1 U29 ( .A(\PG_Network[4][1][47] ), .Z(n18) );
  XNOR2_X1 U30 ( .A(B[35]), .B(n19), .ZN(\PG_Network[0][0][35] ) );
  XNOR2_X1 U31 ( .A(B[27]), .B(n20), .ZN(\PG_Network[0][0][27] ) );
  CLKBUF_X1 U32 ( .A(Co[3]), .Z(n21) );
  XNOR2_X1 U33 ( .A(B[15]), .B(n22), .ZN(\PG_Network[0][0][15] ) );
  XNOR2_X1 U34 ( .A(B[21]), .B(n23), .ZN(\PG_Network[0][0][21] ) );
  XNOR2_X1 U35 ( .A(B[19]), .B(n24), .ZN(\PG_Network[0][0][19] ) );
  XNOR2_X1 U36 ( .A(B[31]), .B(n25), .ZN(\PG_Network[0][0][31] ) );
  XNOR2_X1 U37 ( .A(B[23]), .B(n27), .ZN(\PG_Network[0][0][23] ) );
  XNOR2_X1 U38 ( .A(B[39]), .B(n28), .ZN(\PG_Network[0][0][39] ) );
  XNOR2_X1 U39 ( .A(B[43]), .B(n29), .ZN(\PG_Network[0][0][43] ) );
  CLKBUF_X1 U40 ( .A(\PG_Network[3][0][39] ), .Z(n30) );
  AND2_X1 U41 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U42 ( .A1(A[15]), .A2(B[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U43 ( .A1(A[46]), .A2(B[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U44 ( .A1(A[47]), .A2(B[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U45 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U46 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U47 ( .A1(B[21]), .A2(A[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U48 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U49 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AND2_X1 U50 ( .A1(B[23]), .A2(A[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U51 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U52 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U53 ( .A1(A[35]), .A2(B[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U54 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U55 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U56 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U57 ( .A1(B[27]), .A2(A[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U58 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U59 ( .A1(A[11]), .A2(B[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U60 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U61 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U62 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U63 ( .A1(A[37]), .A2(B[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U64 ( .A1(B[41]), .A2(A[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U65 ( .A1(A[45]), .A2(B[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U66 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U67 ( .A1(A[51]), .A2(B[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U90 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U94 ( .A1(A[49]), .A2(B[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U99 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U100 ( .A1(A[55]), .A2(B[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U101 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U103 ( .A1(B[19]), .A2(A[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U107 ( .A1(B[25]), .A2(A[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U110 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U112 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U116 ( .A1(B[29]), .A2(A[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U118 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U119 ( .A1(A[53]), .A2(B[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U121 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U125 ( .A1(A[59]), .A2(B[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U131 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
  AND2_X1 U132 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U133 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U134 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U135 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U136 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U137 ( .A(n34), .ZN(n31) );
  AND2_X1 U138 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U139 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U140 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U141 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U142 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U143 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U144 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U145 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U146 ( .A1(A[7]), .A2(B[7]), .ZN(\PG_Network[0][1][7] ) );
  AOI21_X1 U147 ( .B1(A[0]), .B2(B[0]), .A(n32), .ZN(n34) );
  INV_X1 U148 ( .A(n33), .ZN(n32) );
  OAI21_X1 U149 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n33) );
  AND2_X1 U150 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U151 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U152 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U153 ( .A1(B[31]), .A2(A[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U154 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AND2_X1 U155 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U156 ( .A1(B[43]), .A2(A[43]), .ZN(\PG_Network[0][1][43] ) );
endmodule


module FA_1408 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1407 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1406 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1405 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_352 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1408 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1407 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1406 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1405 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1404 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1403 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1402 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1401 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_351 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1404 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1403 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1402 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1401 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_176 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U2 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_176 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_352 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_351 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_176 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1400 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1399 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1398 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1397 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_350 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1400 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1399 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1398 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1397 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1396 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1395 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1394 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1393 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_349 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1396 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1395 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1394 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1393 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_175 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_175 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_350 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_349 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_175 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1392 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1391 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1390 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1389 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_348 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1392 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1391 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1390 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1389 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1388 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1387 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1386 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1385 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_347 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1388 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1387 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1386 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1385 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_174 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_174 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_348 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_347 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_174 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1384 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(n5), .B(B), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1383 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1382 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1381 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  OR2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_346 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1384 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1383 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1382 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1381 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1380 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1379 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1378 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1377 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_345 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1380 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1379 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1378 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1377 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_173 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U2 ( .A(sel), .ZN(n13) );
  AOI22_X1 U3 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U6 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U7 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(n17), .ZN(Y[3]) );
endmodule


module carry_select_block_NPB4_173 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_346 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_345 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_173 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1376 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1375 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1374 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1373 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_344 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1376 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1375 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1374 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1373 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1372 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1371 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1370 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1369 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_343 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1372 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1371 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1370 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1369 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_172 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n17), .ZN(Y[2]) );
  BUF_X1 U3 ( .A(n14), .Z(n5) );
  INV_X1 U4 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U6 ( .A(sel), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n5), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
endmodule


module carry_select_block_NPB4_172 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_344 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_343 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_172 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1368 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1367 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1366 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_1365 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_342 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1368 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1367 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1366 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1365 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1364 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1363 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1362 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1361 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_341 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1364 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1363 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1362 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1361 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_171 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n17), .ZN(Y[1]) );
  BUF_X1 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U6 ( .A(n10), .ZN(n5) );
  INV_X1 U7 ( .A(sel), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n15), .ZN(n16) );
endmodule


module carry_select_block_NPB4_171 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_342 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_341 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_171 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1360 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n9), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Co) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n9) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(n7) );
  NAND2_X1 U7 ( .A1(n9), .A2(Ci), .ZN(n8) );
endmodule


module FA_1359 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_1358 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1357 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_340 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1360 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1359 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1358 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1357 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1356 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1355 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1354 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1353 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_339 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1356 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1355 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1354 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1353 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_170 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19, n20;

  INV_X1 U1 ( .A(n19), .ZN(Y[2]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n5) );
  BUF_X1 U4 ( .A(sel), .Z(n11) );
  INV_X1 U5 ( .A(n17), .ZN(Y[0]) );
  INV_X1 U6 ( .A(n20), .ZN(Y[3]) );
  INV_X1 U7 ( .A(n18), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n11), .B1(n5), .B2(B[2]), .ZN(n19) );
  AOI22_X1 U9 ( .A1(n10), .A2(A[1]), .B1(B[1]), .B2(n16), .ZN(n18) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n11), .B1(B[3]), .B2(n5), .ZN(n20) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n16), .ZN(n17) );
  INV_X1 U12 ( .A(sel), .ZN(n16) );
endmodule


module carry_select_block_NPB4_170 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_340 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_339 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_170 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1352 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1351 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1350 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1349 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_338 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1352 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1351 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1350 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1349 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1348 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1347 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1346 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1345 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_337 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1348 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1347 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1346 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1345 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_169 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19, n20;

  INV_X1 U1 ( .A(n18), .ZN(Y[1]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n11) );
  INV_X1 U3 ( .A(sel), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(n10) );
  INV_X1 U5 ( .A(n17), .ZN(Y[0]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n11), .B1(B[2]), .B2(n10), .ZN(n19) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[1]), .B1(n16), .B2(B[1]), .ZN(n18) );
  INV_X1 U9 ( .A(n20), .ZN(Y[3]) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n5), .B2(B[0]), .ZN(n17) );
  INV_X1 U11 ( .A(sel), .ZN(n16) );
  AOI22_X1 U12 ( .A1(A[3]), .A2(n11), .B1(n10), .B2(B[3]), .ZN(n20) );
endmodule


module carry_select_block_NPB4_169 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_338 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_337 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_169 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1344 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n4) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_1343 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1342 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1341 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_336 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1344 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1343 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1342 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1341 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1340 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1339 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1338 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1337 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_335 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1340 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1339 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1338 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1337 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_168 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n17), .ZN(Y[1]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n5) );
  BUF_X1 U3 ( .A(n15), .Z(n10) );
  INV_X1 U4 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n15), .ZN(n17) );
  INV_X1 U8 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n10), .ZN(n19) );
endmodule


module carry_select_block_NPB4_168 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_336 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_335 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_168 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1336 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n5), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1335 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1334 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1333 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(n4), .ZN(n7) );
endmodule


module RCA_N4_334 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1336 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1335 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1334 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1333 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1332 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1331 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1330 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1329 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_333 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1332 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1331 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1330 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1329 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_167 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n17), .ZN(Y[1]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n5) );
  INV_X1 U3 ( .A(sel), .ZN(n10) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U6 ( .A(sel), .ZN(n15) );
  INV_X1 U7 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[1]), .B1(n10), .B2(B[1]), .ZN(n17) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n10), .ZN(n19) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_167 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_334 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_333 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_167 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1328 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6, n7, n8;

  XOR2_X1 U3 ( .A(n8), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n7) );
  OR2_X1 U2 ( .A1(n5), .A2(n6), .ZN(Co) );
  AND2_X1 U4 ( .A1(B), .A2(A), .ZN(n5) );
  AND2_X1 U5 ( .A1(n8), .A2(Ci), .ZN(n6) );
  XNOR2_X1 U6 ( .A(n7), .B(B), .ZN(n8) );
endmodule


module FA_1327 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1326 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1325 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  OR2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_332 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1328 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1327 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1326 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1325 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1324 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1323 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1322 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1321 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_331 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1324 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1323 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1322 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1321 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_166 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  BUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U5 ( .A(sel), .ZN(n14) );
  AOI22_X1 U6 ( .A1(n5), .A2(A[1]), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U7 ( .A1(n5), .A2(A[2]), .B1(B[2]), .B2(n14), .ZN(n17) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
  INV_X1 U9 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n14), .ZN(n18) );
endmodule


module carry_select_block_NPB4_166 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_332 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_331 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_166 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1320 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_1319 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1318 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1317 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_330 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1320 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1319 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1318 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1317 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1316 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1315 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1314 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1313 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_329 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1316 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1315 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1314 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1313 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_165 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(sel), .ZN(n5) );
  BUF_X1 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U6 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(n10), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n15), .ZN(n19) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n5), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_165 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_330 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_329 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_165 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1312 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1311 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1310 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1309 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_328 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1312 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1311 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1310 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1309 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1308 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1307 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1306 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1305 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_327 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1308 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1307 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1306 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1305 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_164 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n10), .ZN(n5) );
  INV_X1 U2 ( .A(n16), .ZN(Y[0]) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n10) );
  INV_X1 U4 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(n10), .A2(A[3]), .B1(B[3]), .B2(n15), .ZN(n19) );
endmodule


module carry_select_block_NPB4_164 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_328 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_327 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_164 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1304 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1303 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1302 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1301 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_326 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1304 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1303 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1302 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1301 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1300 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1299 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1298 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1297 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_325 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1300 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1299 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1298 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1297 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_163 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(sel), .ZN(n13) );
  INV_X1 U3 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U4 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U5 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U7 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_163 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_326 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_325 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_163 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1296 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1295 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1294 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1293 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_324 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1296 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1295 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1294 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1293 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1292 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1291 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1290 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1289 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_323 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1292 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1291 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1290 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1289 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_162 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_162 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_324 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_323 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_162 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1288 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1287 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1286 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1285 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_322 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1288 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1287 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1286 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1285 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1284 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1283 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1282 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1281 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_321 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1284 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1283 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1282 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1281 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_161 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_161 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_322 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_321 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_161 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_11 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_176 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_175 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_174 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_173 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_172 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_171 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_170 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_169 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_168 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_167 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_166 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), .S(S[43:40]) );
  carry_select_block_NPB4_165 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), .S(S[47:44]) );
  carry_select_block_NPB4_164 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), .S(S[51:48]) );
  carry_select_block_NPB4_163 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), .S(S[55:52]) );
  carry_select_block_NPB4_162 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), .S(S[59:56]) );
  carry_select_block_NPB4_161 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), .S(S[63:60]) );
endmodule


module P4_ADDER_N64_11 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_11 CGEN ( .A(A), .B({B[63:45], n4, B[43:41], n14, 
        B[39:37], n16, B[35:33], n17, B[31:29], n19, B[27:25], n2, B[23:21], 
        n15, B[19:17], n18, B[15:13], n1, B[11:0]}), .Cin(Cin), .Co(CoutCgen)
         );
  sum_generator_N64_NPB4_11 SGEN ( .A(A), .B({B[63:44], n8, B[42:40], n9, n3, 
        B[37:36], n7, B[34:32], n5, n10, B[29:28], n6, B[26:24], n13, B[22:20], 
        n11, B[18:16], n12, B[14:0]}), .Ci({CoutCgen, Cin}), .S(S), .Co(Cout)
         );
  CLKBUF_X1 U1 ( .A(B[12]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(B[24]), .Z(n2) );
  CLKBUF_X1 U3 ( .A(B[38]), .Z(n3) );
  CLKBUF_X1 U4 ( .A(B[36]), .Z(n16) );
  CLKBUF_X1 U5 ( .A(B[20]), .Z(n15) );
  CLKBUF_X1 U6 ( .A(B[44]), .Z(n4) );
  CLKBUF_X1 U7 ( .A(B[31]), .Z(n5) );
  CLKBUF_X1 U8 ( .A(B[27]), .Z(n6) );
  CLKBUF_X1 U9 ( .A(B[35]), .Z(n7) );
  CLKBUF_X1 U10 ( .A(B[43]), .Z(n8) );
  CLKBUF_X1 U11 ( .A(B[39]), .Z(n9) );
  BUF_X1 U12 ( .A(B[30]), .Z(n10) );
  CLKBUF_X1 U13 ( .A(B[19]), .Z(n11) );
  CLKBUF_X1 U14 ( .A(B[15]), .Z(n12) );
  CLKBUF_X1 U15 ( .A(B[23]), .Z(n13) );
  CLKBUF_X1 U16 ( .A(B[40]), .Z(n14) );
  CLKBUF_X1 U17 ( .A(B[32]), .Z(n17) );
  CLKBUF_X1 U18 ( .A(B[16]), .Z(n18) );
  CLKBUF_X1 U19 ( .A(B[28]), .Z(n19) );
endmodule


module Booth_Encoder_10 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_10 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306;

  NAND2_X1 U1 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  NAND2_X1 U2 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  NAND2_X1 U3 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  NAND2_X1 U4 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  NAND2_X1 U5 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  NOR3_X1 U6 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U7 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  BUF_X1 U8 ( .A(n158), .Z(n160) );
  BUF_X1 U9 ( .A(n158), .Z(n159) );
  BUF_X1 U10 ( .A(n158), .Z(n162) );
  BUF_X1 U11 ( .A(n158), .Z(n161) );
  BUF_X1 U12 ( .A(n158), .Z(n163) );
  BUF_X1 U13 ( .A(n303), .Z(n158) );
  NOR4_X1 U14 ( .A1(n150), .A2(n144), .A3(n153), .A4(n167), .ZN(n303) );
  BUF_X1 U15 ( .A(n151), .Z(n154) );
  BUF_X1 U16 ( .A(n165), .Z(n168) );
  BUF_X1 U17 ( .A(n151), .Z(n153) );
  BUF_X1 U18 ( .A(n165), .Z(n167) );
  BUF_X1 U19 ( .A(n151), .Z(n155) );
  BUF_X1 U20 ( .A(n152), .Z(n156) );
  BUF_X1 U21 ( .A(n165), .Z(n169) );
  BUF_X1 U22 ( .A(n166), .Z(n170) );
  BUF_X1 U23 ( .A(n152), .Z(n157) );
  BUF_X1 U24 ( .A(n166), .Z(n171) );
  BUF_X1 U25 ( .A(n301), .Z(n149) );
  BUF_X1 U26 ( .A(n304), .Z(n165) );
  BUF_X1 U27 ( .A(n302), .Z(n151) );
  BUF_X1 U28 ( .A(n301), .Z(n148) );
  BUF_X1 U29 ( .A(n301), .Z(n147) );
  BUF_X1 U30 ( .A(n304), .Z(n166) );
  BUF_X1 U31 ( .A(n302), .Z(n152) );
  BUF_X1 U32 ( .A(n301), .Z(n146) );
  BUF_X1 U33 ( .A(n301), .Z(n145) );
  BUF_X1 U34 ( .A(n300), .Z(n139) );
  BUF_X1 U35 ( .A(n300), .Z(n143) );
  BUF_X1 U36 ( .A(n300), .Z(n140) );
  BUF_X1 U37 ( .A(n300), .Z(n142) );
  BUF_X1 U38 ( .A(n300), .Z(n141) );
  INV_X1 U39 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U40 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n304) );
  AND3_X1 U41 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U42 ( .A(sel[2]), .ZN(n173) );
  NAND2_X1 U43 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  AOI22_X1 U44 ( .A1(C[20]), .A2(n149), .B1(A[20]), .B2(n143), .ZN(n199) );
  AOI222_X1 U45 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n154), .ZN(n198) );
  NAND2_X1 U46 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI22_X1 U47 ( .A1(C[23]), .A2(n149), .B1(A[23]), .B2(n143), .ZN(n205) );
  AOI222_X1 U48 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n154), .ZN(n204) );
  NAND2_X1 U49 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI22_X1 U50 ( .A1(C[27]), .A2(n148), .B1(A[27]), .B2(n142), .ZN(n213) );
  AOI222_X1 U51 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n154), .ZN(n212) );
  AOI222_X1 U52 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n153), .ZN(n180) );
  NAND2_X1 U53 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U54 ( .A1(C[14]), .A2(n149), .B1(A[14]), .B2(n143), .ZN(n185) );
  NAND2_X1 U55 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U56 ( .A1(C[15]), .A2(n149), .B1(A[15]), .B2(n143), .ZN(n187) );
  NAND2_X1 U57 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI22_X1 U58 ( .A1(C[17]), .A2(n149), .B1(A[17]), .B2(n143), .ZN(n191) );
  NAND2_X1 U59 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  AOI22_X1 U60 ( .A1(C[48]), .A2(n146), .B1(A[48]), .B2(n140), .ZN(n259) );
  AOI222_X1 U61 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n156), .ZN(n258) );
  NAND2_X1 U62 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI22_X1 U63 ( .A1(C[49]), .A2(n146), .B1(A[49]), .B2(n140), .ZN(n261) );
  AOI222_X1 U64 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n156), .ZN(n260) );
  NAND2_X1 U65 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI22_X1 U66 ( .A1(C[46]), .A2(n146), .B1(A[46]), .B2(n140), .ZN(n255) );
  AOI222_X1 U67 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n156), .ZN(n254) );
  NAND2_X1 U68 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI22_X1 U69 ( .A1(C[18]), .A2(n149), .B1(A[18]), .B2(n143), .ZN(n193) );
  AOI222_X1 U70 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n153), .ZN(n192) );
  NAND2_X1 U71 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U72 ( .A1(C[30]), .A2(n148), .B1(A[30]), .B2(n142), .ZN(n221) );
  AOI222_X1 U73 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n154), .ZN(n220) );
  AOI22_X1 U74 ( .A1(C[32]), .A2(n148), .B1(A[32]), .B2(n142), .ZN(n225) );
  AOI222_X1 U75 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n155), .ZN(n224) );
  NAND2_X1 U76 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI22_X1 U77 ( .A1(C[19]), .A2(n149), .B1(A[19]), .B2(n143), .ZN(n195) );
  AOI222_X1 U78 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n153), .ZN(n194) );
  NAND2_X1 U79 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI22_X1 U80 ( .A1(C[45]), .A2(n147), .B1(A[45]), .B2(n141), .ZN(n253) );
  AOI222_X1 U81 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n156), .ZN(n252) );
  NAND2_X1 U82 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI22_X1 U83 ( .A1(C[47]), .A2(n146), .B1(A[47]), .B2(n140), .ZN(n257) );
  AOI222_X1 U84 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n156), .ZN(n256) );
  NAND2_X1 U85 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI22_X1 U86 ( .A1(C[22]), .A2(n149), .B1(A[22]), .B2(n143), .ZN(n203) );
  AOI222_X1 U87 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n154), .ZN(n202) );
  NAND2_X1 U88 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI22_X1 U89 ( .A1(C[26]), .A2(n148), .B1(A[26]), .B2(n142), .ZN(n211) );
  AOI222_X1 U90 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n154), .ZN(n210) );
  NAND2_X1 U91 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI22_X1 U92 ( .A1(C[34]), .A2(n148), .B1(A[34]), .B2(n142), .ZN(n229) );
  AOI222_X1 U93 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n155), .ZN(n228) );
  NAND2_X1 U94 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI22_X1 U95 ( .A1(C[38]), .A2(n147), .B1(A[38]), .B2(n141), .ZN(n237) );
  AOI222_X1 U96 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n155), .ZN(n236) );
  NAND2_X1 U97 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI22_X1 U98 ( .A1(C[42]), .A2(n147), .B1(A[42]), .B2(n141), .ZN(n247) );
  AOI222_X1 U99 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n155), .ZN(n246) );
  AOI22_X1 U100 ( .A1(C[28]), .A2(n148), .B1(A[28]), .B2(n142), .ZN(n215) );
  AOI222_X1 U101 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n154), .ZN(n214) );
  NAND2_X1 U102 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI22_X1 U103 ( .A1(C[21]), .A2(n149), .B1(A[21]), .B2(n143), .ZN(n201) );
  AOI222_X1 U104 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n154), .ZN(n200) );
  NAND2_X1 U105 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI222_X1 U106 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n154), .ZN(n208) );
  AOI22_X1 U107 ( .A1(C[25]), .A2(n148), .B1(A[25]), .B2(n142), .ZN(n209) );
  NAND2_X1 U108 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI222_X1 U109 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n154), .ZN(n216) );
  AOI22_X1 U110 ( .A1(C[29]), .A2(n148), .B1(A[29]), .B2(n142), .ZN(n217) );
  NAND2_X1 U111 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI222_X1 U112 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n155), .ZN(n226) );
  AOI22_X1 U113 ( .A1(C[33]), .A2(n148), .B1(A[33]), .B2(n142), .ZN(n227) );
  NAND2_X1 U114 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI222_X1 U115 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n155), .ZN(n234) );
  AOI22_X1 U116 ( .A1(C[37]), .A2(n147), .B1(A[37]), .B2(n141), .ZN(n235) );
  NAND2_X1 U117 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  AOI22_X1 U118 ( .A1(C[16]), .A2(n149), .B1(A[16]), .B2(n143), .ZN(n189) );
  AOI222_X1 U119 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n153), .ZN(n188) );
  AOI22_X1 U120 ( .A1(C[36]), .A2(n147), .B1(A[36]), .B2(n141), .ZN(n233) );
  AOI222_X1 U121 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n155), .ZN(n232) );
  NAND2_X1 U122 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI222_X1 U123 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n155), .ZN(n230) );
  NAND2_X1 U124 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI222_X1 U125 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n155), .ZN(n238) );
  AOI222_X1 U126 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n156), .ZN(n250) );
  AOI22_X1 U127 ( .A1(C[44]), .A2(n147), .B1(A[44]), .B2(n141), .ZN(n251) );
  NAND2_X1 U128 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI222_X1 U129 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n155), .ZN(n248) );
  NAND2_X1 U130 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  AOI222_X1 U131 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n155), .ZN(n242) );
  AOI22_X1 U132 ( .A1(C[24]), .A2(n149), .B1(A[24]), .B2(n143), .ZN(n207) );
  AOI222_X1 U133 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n154), .ZN(n206) );
  NAND2_X1 U134 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI22_X1 U135 ( .A1(C[31]), .A2(n148), .B1(A[31]), .B2(n142), .ZN(n223) );
  AOI222_X1 U136 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n154), .ZN(n222) );
  NAND2_X1 U137 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI222_X1 U138 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n155), .ZN(n244) );
  AOI22_X1 U139 ( .A1(C[41]), .A2(n147), .B1(A[41]), .B2(n141), .ZN(n245) );
  NAND2_X1 U140 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  AOI22_X1 U141 ( .A1(C[52]), .A2(n146), .B1(A[52]), .B2(n140), .ZN(n269) );
  AOI222_X1 U142 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n156), .ZN(n268) );
  NAND2_X1 U143 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  AOI22_X1 U144 ( .A1(C[56]), .A2(n146), .B1(A[56]), .B2(n140), .ZN(n277) );
  AOI222_X1 U145 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n157), .ZN(n276) );
  NAND2_X1 U146 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  AOI22_X1 U147 ( .A1(C[53]), .A2(n146), .B1(A[53]), .B2(n140), .ZN(n271) );
  AOI222_X1 U148 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n156), .ZN(n270) );
  NAND2_X1 U149 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI22_X1 U150 ( .A1(C[54]), .A2(n146), .B1(A[54]), .B2(n140), .ZN(n273) );
  AOI222_X1 U151 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n156), .ZN(n272) );
  NAND2_X1 U152 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  AOI22_X1 U153 ( .A1(C[51]), .A2(n146), .B1(A[51]), .B2(n140), .ZN(n267) );
  AOI222_X1 U154 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n156), .ZN(n266) );
  NAND2_X1 U155 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI22_X1 U156 ( .A1(C[55]), .A2(n146), .B1(A[55]), .B2(n140), .ZN(n275) );
  AOI222_X1 U157 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n156), .ZN(n274) );
  NAND2_X1 U158 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI22_X1 U159 ( .A1(C[50]), .A2(n146), .B1(A[50]), .B2(n140), .ZN(n265) );
  AOI222_X1 U160 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n156), .ZN(n264) );
  NAND2_X1 U161 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U162 ( .A1(C[60]), .A2(n145), .B1(A[60]), .B2(n139), .ZN(n287) );
  AOI222_X1 U163 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n157), .ZN(n286) );
  NAND2_X1 U164 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  AOI22_X1 U165 ( .A1(C[57]), .A2(n145), .B1(A[57]), .B2(n139), .ZN(n279) );
  AOI222_X1 U166 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n157), .ZN(n278) );
  NAND2_X1 U167 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U168 ( .A1(C[61]), .A2(n145), .B1(A[61]), .B2(n139), .ZN(n289) );
  AOI222_X1 U169 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n157), .ZN(n288) );
  NAND2_X1 U170 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI22_X1 U171 ( .A1(C[58]), .A2(n145), .B1(A[58]), .B2(n139), .ZN(n281) );
  AOI222_X1 U172 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n157), .ZN(n280) );
  NAND2_X1 U173 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U174 ( .A1(C[62]), .A2(n145), .B1(A[62]), .B2(n139), .ZN(n291) );
  AOI222_X1 U175 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n157), .ZN(n290) );
  NAND2_X1 U176 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U177 ( .A1(C[59]), .A2(n145), .B1(A[59]), .B2(n139), .ZN(n283) );
  AOI222_X1 U178 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n157), .ZN(n282) );
  NAND2_X1 U179 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U180 ( .A1(C[63]), .A2(n145), .B1(A[63]), .B2(n139), .ZN(n293) );
  AOI222_X1 U181 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n157), .ZN(n292) );
  NAND2_X1 U182 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U183 ( .A1(C[0]), .A2(n145), .B1(A[0]), .B2(n139), .ZN(n175) );
  AOI222_X1 U184 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n153), .ZN(n174) );
  NAND2_X1 U185 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U186 ( .A1(C[4]), .A2(n146), .B1(A[4]), .B2(n140), .ZN(n263) );
  AOI222_X1 U187 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n156), .ZN(n262) );
  NAND2_X1 U188 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI22_X1 U189 ( .A1(C[8]), .A2(n145), .B1(A[8]), .B2(n139), .ZN(n299) );
  AOI222_X1 U190 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n157), .ZN(n298) );
  NAND2_X1 U191 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U192 ( .A1(C[1]), .A2(n149), .B1(A[1]), .B2(n143), .ZN(n197) );
  AOI222_X1 U193 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n153), .ZN(n196) );
  NAND2_X1 U194 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U195 ( .A1(C[5]), .A2(n145), .B1(A[5]), .B2(n139), .ZN(n285) );
  AOI222_X1 U196 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n157), .ZN(n284) );
  NAND2_X1 U197 ( .A1(n306), .A2(n305), .ZN(Y[9]) );
  AOI22_X1 U198 ( .A1(C[9]), .A2(n147), .B1(A[9]), .B2(n141), .ZN(n306) );
  AOI222_X1 U199 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n157), .ZN(n305) );
  NAND2_X1 U200 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U201 ( .A1(C[2]), .A2(n148), .B1(A[2]), .B2(n142), .ZN(n219) );
  AOI222_X1 U202 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n154), .ZN(n218) );
  NAND2_X1 U203 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U204 ( .A1(C[6]), .A2(n145), .B1(A[6]), .B2(n139), .ZN(n295) );
  AOI222_X1 U205 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n157), .ZN(n294) );
  NAND2_X1 U206 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U207 ( .A1(C[10]), .A2(n150), .B1(A[10]), .B2(n144), .ZN(n177) );
  AOI222_X1 U208 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n153), .ZN(n176) );
  NAND2_X1 U209 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U210 ( .A1(C[3]), .A2(n147), .B1(A[3]), .B2(n141), .ZN(n241) );
  AOI222_X1 U211 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n155), .ZN(n240) );
  NAND2_X1 U212 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U213 ( .A1(C[7]), .A2(n145), .B1(A[7]), .B2(n139), .ZN(n297) );
  AOI222_X1 U214 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n157), .ZN(n296) );
  NAND2_X1 U215 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U216 ( .A1(C[11]), .A2(n150), .B1(A[11]), .B2(n144), .ZN(n179) );
  AOI222_X1 U217 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n153), .ZN(n178) );
  AOI22_X1 U218 ( .A1(C[40]), .A2(n147), .B1(A[40]), .B2(n141), .ZN(n243) );
  AOI22_X1 U219 ( .A1(C[39]), .A2(n147), .B1(A[39]), .B2(n141), .ZN(n239) );
  AOI22_X1 U220 ( .A1(C[12]), .A2(n150), .B1(A[12]), .B2(n144), .ZN(n181) );
  AOI22_X1 U221 ( .A1(C[13]), .A2(n150), .B1(A[13]), .B2(n144), .ZN(n183) );
  NAND2_X1 U222 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  NAND2_X1 U223 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI222_X1 U224 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n153), .ZN(n190) );
  AOI22_X1 U225 ( .A1(C[35]), .A2(n148), .B1(A[35]), .B2(n142), .ZN(n231) );
  AOI222_X1 U226 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n153), .ZN(n184) );
  AOI222_X1 U227 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n153), .ZN(n182) );
  AOI22_X1 U228 ( .A1(C[43]), .A2(n147), .B1(A[43]), .B2(n141), .ZN(n249) );
  AOI222_X1 U229 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n153), .ZN(n186) );
  CLKBUF_X1 U230 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U231 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U232 ( .A(n158), .Z(n164) );
endmodule


module G_170 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_630 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_629 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_628 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_627 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_626 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_625 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_624 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_623 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_622 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_621 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_620 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_619 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_618 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_617 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_616 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_615 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_614 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_613 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_612 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_611 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_610 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_609 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_608 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_607 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_606 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_605 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_604 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_603 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_602 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_601 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_600 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_169 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_599 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_598 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_597 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_596 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_595 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_594 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_593 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_592 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_591 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_590 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_589 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_588 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_587 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_586 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_585 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_168 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_584 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_583 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_582 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3, n5;

  CLKBUF_X1 U1 ( .A(P_IK), .Z(n3) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n5), .ZN(Gx) );
  AOI21_X1 U4 ( .B1(G_K_1), .B2(n3), .A(G_IK), .ZN(n5) );
endmodule


module PG_581 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_580 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_579 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_578 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_167 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n3;

  OR2_X2 U1 ( .A1(G_IK), .A2(n3), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n3) );
endmodule


module G_166 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_577 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_576 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_575 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  OR2_X1 U2 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_574 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_573 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_572 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_165 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  OR2_X2 U2 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
endmodule


module G_164 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_163 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_162 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module PG_571 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_570 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_569 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_568 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_161 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_160 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_159 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_158 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  OR2_X1 U2 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
endmodule


module G_157 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_156 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_155 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_154 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module carry_generator_N64_NPB4_10 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U77 ( .A(B[59]), .B(A[59]), .Z(\PG_Network[0][0][59] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U81 ( .A(B[55]), .B(A[55]), .Z(\PG_Network[0][0][55] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U85 ( .A(B[51]), .B(A[51]), .Z(\PG_Network[0][0][51] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U88 ( .A(B[49]), .B(A[49]), .Z(\PG_Network[0][0][49] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U91 ( .A(B[46]), .B(A[46]), .Z(\PG_Network[0][0][46] ) );
  XOR2_X1 U92 ( .A(B[45]), .B(A[45]), .Z(\PG_Network[0][0][45] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U100 ( .A(B[38]), .B(A[38]), .Z(\PG_Network[0][0][38] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_170 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n26), .Gx(\PG_Network[1][1][1] ) );
  PG_630 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_629 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_628 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_627 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_626 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_625 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_624 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_623 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_622 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_621 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_620 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_619 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_618 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_617 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_616 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_615 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_614 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_613 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_612 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_611 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_610 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_609 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_608 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_607 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_606 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_605 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_604 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_603 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_602 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_601 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_600 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_169 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_599 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_598 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_597 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_596 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_595 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_594 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_593 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_592 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_591 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_590 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_589 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_588 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_587 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_586 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_585 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_168 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_584 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_583 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_582 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_581 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_580 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_579 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_578 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_167 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), .G_K_1(Co[1]), .Gx(Co[3]) );
  G_166 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_577 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_576 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_575 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(n6), .P_K_1(\PG_Network[3][0][39] ), 
        .Gx(\PG_Network[4][1][47] ), .Px(\PG_Network[4][0][47] ) );
  PG_574 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][43] ), .Px(
        \PG_Network[4][0][43] ) );
  PG_573 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][63] ), .Px(
        \PG_Network[4][0][63] ) );
  PG_572 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][59] ), .Px(
        \PG_Network[4][0][59] ) );
  G_165 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), .G_K_1(Co[3]), .Gx(Co[7]) );
  G_164 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), .G_K_1(Co[3]), .Gx(Co[6]) );
  G_163 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), .G_K_1(Co[3]), .Gx(Co[5]) );
  G_162 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), .G_K_1(Co[3]), .Gx(Co[4]) );
  PG_571 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(n17), .P_K_1(n9), .Gx(
        \PG_Network[5][1][63] ), .Px(\PG_Network[5][0][63] ) );
  PG_570 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(n17), .P_K_1(n9), .Gx(
        \PG_Network[5][1][59] ), .Px(\PG_Network[5][0][59] ) );
  PG_569 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(n17), .P_K_1(n9), .Gx(
        \PG_Network[5][1][55] ), .Px(\PG_Network[5][0][55] ) );
  PG_568 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(n17), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][51] ), .Px(\PG_Network[5][0][51] ) );
  G_161 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), .G_K_1(n19), .Gx(Co[15]) );
  G_160 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), .G_K_1(n19), .Gx(Co[14]) );
  G_159 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), .G_K_1(n19), .Gx(Co[13]) );
  G_158 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), .G_K_1(n19), .Gx(Co[12]) );
  G_157 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), .G_K_1(Co[7]), .Gx(Co[11]) );
  G_156 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), .G_K_1(Co[7]), .Gx(Co[10]) );
  G_155 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), .G_K_1(Co[7]), .Gx(Co[9]) );
  G_154 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), .G_K_1(Co[7]), .Gx(Co[8]) );
  CLKBUF_X1 U1 ( .A(B[42]), .Z(n5) );
  CLKBUF_X1 U2 ( .A(\PG_Network[3][1][39] ), .Z(n6) );
  INV_X1 U3 ( .A(A[47]), .ZN(n13) );
  INV_X1 U4 ( .A(A[26]), .ZN(n8) );
  INV_X1 U5 ( .A(A[37]), .ZN(n10) );
  INV_X1 U6 ( .A(A[35]), .ZN(n11) );
  INV_X1 U7 ( .A(A[23]), .ZN(n23) );
  INV_X1 U8 ( .A(A[27]), .ZN(n18) );
  INV_X1 U9 ( .A(A[15]), .ZN(n15) );
  INV_X1 U10 ( .A(A[30]), .ZN(n14) );
  INV_X1 U11 ( .A(A[19]), .ZN(n12) );
  INV_X1 U12 ( .A(A[25]), .ZN(n7) );
  INV_X1 U13 ( .A(A[29]), .ZN(n22) );
  INV_X1 U14 ( .A(A[39]), .ZN(n20) );
  INV_X1 U15 ( .A(A[43]), .ZN(n25) );
  INV_X1 U16 ( .A(A[31]), .ZN(n21) );
  INV_X1 U17 ( .A(A[41]), .ZN(n24) );
  INV_X1 U18 ( .A(A[36]), .ZN(n16) );
  XNOR2_X1 U19 ( .A(B[25]), .B(n7), .ZN(\PG_Network[0][0][25] ) );
  XNOR2_X1 U20 ( .A(B[26]), .B(n8), .ZN(\PG_Network[0][0][26] ) );
  CLKBUF_X1 U21 ( .A(\PG_Network[4][0][47] ), .Z(n9) );
  XNOR2_X1 U22 ( .A(B[37]), .B(n10), .ZN(\PG_Network[0][0][37] ) );
  XNOR2_X1 U23 ( .A(B[35]), .B(n11), .ZN(\PG_Network[0][0][35] ) );
  XNOR2_X1 U24 ( .A(B[19]), .B(n12), .ZN(\PG_Network[0][0][19] ) );
  XNOR2_X1 U25 ( .A(B[47]), .B(n13), .ZN(\PG_Network[0][0][47] ) );
  XNOR2_X1 U26 ( .A(B[30]), .B(n14), .ZN(\PG_Network[0][0][30] ) );
  XNOR2_X1 U27 ( .A(B[15]), .B(n15), .ZN(\PG_Network[0][0][15] ) );
  XNOR2_X1 U28 ( .A(B[36]), .B(n16), .ZN(\PG_Network[0][0][36] ) );
  CLKBUF_X1 U29 ( .A(\PG_Network[4][1][47] ), .Z(n17) );
  XNOR2_X1 U30 ( .A(B[27]), .B(n18), .ZN(\PG_Network[0][0][27] ) );
  CLKBUF_X1 U31 ( .A(Co[7]), .Z(n19) );
  XNOR2_X1 U32 ( .A(B[39]), .B(n20), .ZN(\PG_Network[0][0][39] ) );
  XNOR2_X1 U33 ( .A(B[31]), .B(n21), .ZN(\PG_Network[0][0][31] ) );
  XNOR2_X1 U34 ( .A(B[29]), .B(n22), .ZN(\PG_Network[0][0][29] ) );
  XNOR2_X1 U35 ( .A(B[23]), .B(n23), .ZN(\PG_Network[0][0][23] ) );
  XNOR2_X1 U36 ( .A(B[41]), .B(n24), .ZN(\PG_Network[0][0][41] ) );
  XNOR2_X1 U37 ( .A(B[43]), .B(n25), .ZN(\PG_Network[0][0][43] ) );
  AND2_X1 U38 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U39 ( .A1(A[51]), .A2(B[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U40 ( .A1(A[42]), .A2(n5), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U41 ( .A1(B[30]), .A2(A[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U42 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U43 ( .A1(B[19]), .A2(A[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U44 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U45 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AND2_X1 U46 ( .A1(B[23]), .A2(A[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U47 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U48 ( .A1(A[46]), .A2(B[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U49 ( .A1(A[47]), .A2(B[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U50 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AND2_X1 U51 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U52 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U53 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U54 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U55 ( .A1(A[21]), .A2(B[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U56 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U57 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U58 ( .A1(B[25]), .A2(A[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U59 ( .A1(A[45]), .A2(B[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U60 ( .A1(A[49]), .A2(B[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U61 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U62 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U63 ( .A1(A[55]), .A2(B[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U64 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U65 ( .A1(A[59]), .A2(B[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U66 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
  AND2_X1 U67 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U90 ( .A1(B[26]), .A2(A[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U94 ( .A1(B[27]), .A2(A[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U96 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U99 ( .A1(B[29]), .A2(A[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U101 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U102 ( .A1(A[53]), .A2(B[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U103 ( .A1(A[37]), .A2(B[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U107 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U108 ( .A1(B[15]), .A2(A[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U110 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U112 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U113 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U114 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U116 ( .A1(A[11]), .A2(B[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U121 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U125 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U131 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U132 ( .A(n29), .ZN(n26) );
  AND2_X1 U133 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U134 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U135 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U136 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U137 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U138 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U139 ( .A1(A[7]), .A2(B[7]), .ZN(\PG_Network[0][1][7] ) );
  AOI21_X1 U140 ( .B1(A[0]), .B2(B[0]), .A(n27), .ZN(n29) );
  INV_X1 U141 ( .A(n28), .ZN(n27) );
  OAI21_X1 U142 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n28) );
  AND2_X1 U143 ( .A1(B[31]), .A2(A[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U144 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U145 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U146 ( .A1(A[35]), .A2(B[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U147 ( .A1(B[41]), .A2(A[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U148 ( .A1(B[43]), .A2(A[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U149 ( .A1(B[24]), .A2(A[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U150 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U151 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
endmodule


module FA_1280 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1279 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1278 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1277 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_320 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1280 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1279 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1278 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1277 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1276 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1275 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1274 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1273 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_319 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1276 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1275 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1274 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1273 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_160 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U2 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_160 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_320 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_319 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_160 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1272 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1271 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1270 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1269 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_318 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1272 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1271 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1270 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1269 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1268 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1267 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1266 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1265 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_317 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1268 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1267 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1266 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1265 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_159 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_159 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_318 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_317 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_159 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1264 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1263 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1262 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1261 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_316 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1264 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1263 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1262 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1261 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1260 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1259 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1258 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1257 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_315 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1260 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1259 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1258 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1257 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_158 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_158 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_316 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_315 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_158 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1256 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_314 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1256 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1255 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1254 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1253 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1252 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1251 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1250 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1249 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_313 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1252 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1251 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1250 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1249 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_157 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_157 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_314 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_313 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_157 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_312 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1248 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1247 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1246 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1245 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1244 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1243 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1242 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1241 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_311 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1244 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1243 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1242 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1241 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_156 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U3 ( .A(sel), .ZN(n5) );
  INV_X1 U4 ( .A(n16), .ZN(Y[0]) );
  CLKBUF_X1 U5 ( .A(sel), .Z(n10) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(n10), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n5), .ZN(n16) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n15), .ZN(n19) );
endmodule


module carry_select_block_NPB4_156 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_312 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_311 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_156 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n5) );
  AOI22_X1 U5 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_1239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_310 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1240 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1239 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1238 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1237 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1236 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1235 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1234 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1233 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_309 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1236 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1235 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1234 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1233 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_155 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n17), .ZN(Y[2]) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n5) );
  INV_X1 U4 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n14), .ZN(n17) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n14), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
  INV_X1 U10 ( .A(sel), .ZN(n14) );
endmodule


module carry_select_block_NPB4_155 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_310 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_309 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_155 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n8), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_1231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_308 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1232 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1231 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1230 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1229 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1228 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1227 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1226 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1225 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_307 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1228 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1227 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1226 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1225 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_154 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n16), .ZN(Y[0]) );
  INV_X2 U2 ( .A(n18), .ZN(Y[2]) );
  BUF_X1 U3 ( .A(n15), .Z(n5) );
  BUF_X1 U4 ( .A(sel), .Z(n10) );
  INV_X1 U5 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U6 ( .A(sel), .ZN(n15) );
  INV_X1 U7 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(n10), .A2(A[2]), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U9 ( .A1(n10), .A2(A[1]), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
endmodule


module carry_select_block_NPB4_154 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_308 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_307 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_154 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_1223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n8, n10, n11;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n10) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n5), .A2(n10), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n8), .A2(n7), .ZN(S) );
  INV_X1 U6 ( .A(Ci), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(n6) );
  INV_X1 U8 ( .A(n11), .ZN(Co) );
  AOI22_X1 U9 ( .A1(B), .A2(A), .B1(n10), .B2(n4), .ZN(n11) );
endmodule


module RCA_N4_306 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1224 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1223 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1222 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1221 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1220 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1219 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1218 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1217 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_305 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1220 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1219 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1218 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1217 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_153 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19, n20;

  INV_X2 U1 ( .A(n18), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n17), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n11), .ZN(n5) );
  BUF_X1 U4 ( .A(sel), .Z(n11) );
  CLKBUF_X1 U5 ( .A(n16), .Z(n10) );
  INV_X1 U6 ( .A(n19), .ZN(Y[2]) );
  INV_X1 U7 ( .A(n20), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n11), .B1(B[2]), .B2(n5), .ZN(n19) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n16), .ZN(n18) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n11), .B1(B[3]), .B2(n10), .ZN(n20) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n16), .B2(B[0]), .ZN(n17) );
  INV_X1 U12 ( .A(sel), .ZN(n16) );
endmodule


module carry_select_block_NPB4_153 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_306 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_305 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_153 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1216 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(n4), .ZN(n8) );
  CLKBUF_X1 U4 ( .A(B), .Z(n5) );
  XOR2_X1 U5 ( .A(A), .B(n5), .Z(n6) );
  AOI22_X1 U6 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_1215 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1214 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1213 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_304 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1216 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1215 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1214 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1213 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1212 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1211 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1210 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1209 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_303 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1212 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1211 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1210 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1209 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_152 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U2 ( .A(sel), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n10) );
  INV_X1 U4 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n5), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
endmodule


module carry_select_block_NPB4_152 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_304 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_303 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_152 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1208 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_1207 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1206 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1205 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_302 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1208 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1207 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1206 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1205 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1204 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1203 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1202 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1201 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_301 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1204 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1203 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1202 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1201 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_151 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n16), .ZN(Y[0]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(sel), .ZN(n5) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n15), .ZN(n18) );
  INV_X1 U7 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[1]), .B1(n15), .B2(B[1]), .ZN(n17) );
  INV_X1 U9 ( .A(sel), .ZN(n15) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n15), .ZN(n19) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n5), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_151 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_302 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_301 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_151 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1200 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  XOR2_X1 U2 ( .A(A), .B(n4), .Z(n5) );
  AOI22_X1 U5 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_1199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_300 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1200 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1199 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1198 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1197 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1196 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1195 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  XOR2_X1 U2 ( .A(A), .B(n4), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1194 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1193 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_299 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1196 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1195 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1194 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1193 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_150 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(sel), .ZN(n5) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n5), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(n15), .B2(B[0]), .ZN(n16) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
endmodule


module carry_select_block_NPB4_150 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_300 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_299 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_150 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1192 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n7), .Z(S) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1191 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1190 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1189 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_298 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1192 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1191 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1190 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1189 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1188 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1187 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1186 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1185 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_297 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1188 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1187 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1186 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1185 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_149 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19, n20;

  CLKBUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(n17), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n5), .ZN(n10) );
  CLKBUF_X1 U4 ( .A(n5), .Z(n11) );
  INV_X1 U5 ( .A(n19), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n18), .ZN(Y[1]) );
  INV_X1 U7 ( .A(n20), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n11), .B1(B[2]), .B2(n10), .ZN(n19) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(n16), .B2(B[1]), .ZN(n18) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n11), .B1(B[3]), .B2(n10), .ZN(n20) );
  AOI22_X1 U11 ( .A1(A[0]), .A2(sel), .B1(n16), .B2(B[0]), .ZN(n17) );
  INV_X1 U12 ( .A(sel), .ZN(n16) );
endmodule


module carry_select_block_NPB4_149 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_298 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_297 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_149 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1184 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1183 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1182 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1181 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_296 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1184 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1183 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1182 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1181 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1180 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1179 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1178 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1177 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_295 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1180 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1179 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1178 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1177 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_148 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  CLKBUF_X1 U1 ( .A(n14), .Z(n5) );
  INV_X1 U2 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n16), .ZN(Y[1]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n17) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
  INV_X1 U10 ( .A(sel), .ZN(n14) );
endmodule


module carry_select_block_NPB4_148 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_296 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_295 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_148 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1176 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1175 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1174 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1173 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_294 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1176 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1175 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1174 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1173 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1172 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1171 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1170 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1169 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_293 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1172 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1171 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1170 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1169 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_147 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(sel), .ZN(n13) );
  INV_X1 U3 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U4 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U5 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U7 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_147 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_294 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_293 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_147 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1168 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1167 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1166 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1165 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_292 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1168 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1167 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1166 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1165 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1164 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1163 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1162 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1161 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_291 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1164 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1163 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1162 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1161 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_146 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_146 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_292 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_291 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_146 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1160 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1159 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1158 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1157 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_290 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1160 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1159 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1158 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1157 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1156 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1155 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1154 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1153 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_289 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1156 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1155 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1154 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1153 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_145 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_145 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_290 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_289 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_145 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_10 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_160 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_159 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_158 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_157 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_156 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_155 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_154 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_153 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_152 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_151 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_150 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), .S(S[43:40]) );
  carry_select_block_NPB4_149 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), .S(S[47:44]) );
  carry_select_block_NPB4_148 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), .S(S[51:48]) );
  carry_select_block_NPB4_147 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), .S(S[55:52]) );
  carry_select_block_NPB4_146 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), .S(S[59:56]) );
  carry_select_block_NPB4_145 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), .S(S[63:60]) );
endmodule


module P4_ADDER_N64_10 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_10 CGEN ( .A(A), .B({B[63:49], n3, B[47:37], n25, 
        B[35:33], n21, B[31:29], n17, B[27:25], n22, B[23:21], n16, B[19:17], 
        n24, B[15:0]}), .Cin(Cin), .Co(CoutCgen) );
  sum_generator_N64_NPB4_10 SGEN ( .A(A), .B({B[63:48], n13, B[46:44], n15, 
        B[42], n6, B[40], n19, n5, B[37:36], n20, B[34:32], n8, n14, B[29:28], 
        n23, n1, B[25:24], n4, n11, B[21:20], n10, B[18:16], n18, B[14:0]}), 
        .Ci({CoutCgen, Cin}), .S(S), .Co(Cout) );
  BUF_X1 U1 ( .A(B[22]), .Z(n11) );
  BUF_X1 U2 ( .A(B[30]), .Z(n14) );
  BUF_X1 U3 ( .A(B[41]), .Z(n6) );
  CLKBUF_X1 U4 ( .A(B[26]), .Z(n1) );
  CLKBUF_X1 U5 ( .A(B[47]), .Z(n2) );
  CLKBUF_X1 U6 ( .A(B[48]), .Z(n3) );
  CLKBUF_X1 U7 ( .A(B[23]), .Z(n4) );
  CLKBUF_X1 U8 ( .A(B[38]), .Z(n5) );
  INV_X1 U9 ( .A(B[31]), .ZN(n7) );
  INV_X1 U10 ( .A(n7), .ZN(n8) );
  INV_X1 U11 ( .A(B[19]), .ZN(n9) );
  INV_X1 U12 ( .A(n9), .ZN(n10) );
  CLKBUF_X1 U13 ( .A(B[15]), .Z(n18) );
  CLKBUF_X1 U14 ( .A(B[28]), .Z(n17) );
  CLKBUF_X1 U15 ( .A(B[36]), .Z(n25) );
  CLKBUF_X1 U16 ( .A(B[24]), .Z(n22) );
  INV_X1 U17 ( .A(n2), .ZN(n12) );
  INV_X1 U18 ( .A(n12), .ZN(n13) );
  CLKBUF_X1 U19 ( .A(B[43]), .Z(n15) );
  CLKBUF_X1 U20 ( .A(B[20]), .Z(n16) );
  CLKBUF_X1 U21 ( .A(B[39]), .Z(n19) );
  CLKBUF_X1 U22 ( .A(B[35]), .Z(n20) );
  CLKBUF_X1 U23 ( .A(B[32]), .Z(n21) );
  CLKBUF_X1 U24 ( .A(B[27]), .Z(n23) );
  CLKBUF_X1 U25 ( .A(B[16]), .Z(n24) );
endmodule


module Booth_Encoder_9 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_9 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306;

  NAND2_X1 U1 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  NAND2_X1 U2 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  NAND2_X1 U3 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  NAND2_X1 U4 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  NAND2_X1 U5 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  NOR3_X1 U6 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U7 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  NAND2_X2 U8 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  BUF_X1 U9 ( .A(n158), .Z(n159) );
  BUF_X1 U10 ( .A(n158), .Z(n162) );
  BUF_X1 U11 ( .A(n158), .Z(n161) );
  BUF_X1 U12 ( .A(n158), .Z(n160) );
  BUF_X1 U13 ( .A(n158), .Z(n163) );
  BUF_X1 U14 ( .A(n303), .Z(n158) );
  NOR4_X1 U15 ( .A1(n150), .A2(n144), .A3(n153), .A4(n167), .ZN(n303) );
  BUF_X1 U16 ( .A(n151), .Z(n154) );
  BUF_X1 U17 ( .A(n151), .Z(n155) );
  BUF_X1 U18 ( .A(n165), .Z(n168) );
  BUF_X1 U19 ( .A(n165), .Z(n169) );
  BUF_X1 U20 ( .A(n151), .Z(n153) );
  BUF_X1 U21 ( .A(n165), .Z(n167) );
  BUF_X1 U22 ( .A(n152), .Z(n156) );
  BUF_X1 U23 ( .A(n166), .Z(n170) );
  BUF_X1 U24 ( .A(n152), .Z(n157) );
  BUF_X1 U25 ( .A(n166), .Z(n171) );
  BUF_X1 U26 ( .A(n301), .Z(n148) );
  BUF_X1 U27 ( .A(n301), .Z(n149) );
  BUF_X1 U28 ( .A(n304), .Z(n165) );
  BUF_X1 U29 ( .A(n302), .Z(n151) );
  BUF_X1 U30 ( .A(n301), .Z(n146) );
  BUF_X1 U31 ( .A(n301), .Z(n147) );
  BUF_X1 U32 ( .A(n304), .Z(n166) );
  BUF_X1 U33 ( .A(n302), .Z(n152) );
  BUF_X1 U34 ( .A(n301), .Z(n145) );
  BUF_X1 U35 ( .A(n300), .Z(n142) );
  BUF_X1 U36 ( .A(n300), .Z(n139) );
  BUF_X1 U37 ( .A(n300), .Z(n140) );
  BUF_X1 U38 ( .A(n300), .Z(n143) );
  BUF_X1 U39 ( .A(n300), .Z(n141) );
  INV_X1 U40 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U41 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n304) );
  AND3_X1 U42 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U43 ( .A(sel[2]), .ZN(n173) );
  AOI222_X1 U44 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n153), .ZN(n184) );
  NAND2_X1 U45 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI22_X1 U46 ( .A1(C[17]), .A2(n149), .B1(A[17]), .B2(n143), .ZN(n191) );
  NAND2_X1 U47 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI22_X1 U48 ( .A1(C[19]), .A2(n149), .B1(A[19]), .B2(n143), .ZN(n195) );
  NAND2_X1 U49 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI22_X1 U50 ( .A1(C[22]), .A2(n149), .B1(A[22]), .B2(n143), .ZN(n203) );
  AOI222_X1 U51 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n154), .ZN(n202) );
  NAND2_X1 U52 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  AOI22_X1 U53 ( .A1(C[53]), .A2(n146), .B1(A[53]), .B2(n140), .ZN(n271) );
  AOI222_X1 U54 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n156), .ZN(n270) );
  NAND2_X1 U55 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI22_X1 U56 ( .A1(C[54]), .A2(n146), .B1(A[54]), .B2(n140), .ZN(n273) );
  AOI222_X1 U57 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n156), .ZN(n272) );
  NAND2_X1 U58 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI22_X1 U59 ( .A1(C[55]), .A2(n146), .B1(A[55]), .B2(n140), .ZN(n275) );
  AOI222_X1 U60 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n156), .ZN(n274) );
  NAND2_X1 U61 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI22_X1 U62 ( .A1(C[23]), .A2(n149), .B1(A[23]), .B2(n143), .ZN(n205) );
  AOI222_X1 U63 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n154), .ZN(n204) );
  NAND2_X1 U64 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI222_X1 U65 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n154), .ZN(n212) );
  AOI22_X1 U66 ( .A1(C[27]), .A2(n148), .B1(A[27]), .B2(n142), .ZN(n213) );
  NAND2_X1 U67 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI222_X1 U68 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n154), .ZN(n222) );
  AOI22_X1 U69 ( .A1(C[31]), .A2(n148), .B1(A[31]), .B2(n142), .ZN(n223) );
  NAND2_X1 U70 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI22_X1 U71 ( .A1(C[21]), .A2(n149), .B1(A[21]), .B2(n143), .ZN(n201) );
  AOI222_X1 U72 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n154), .ZN(n200) );
  NAND2_X1 U73 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI22_X1 U74 ( .A1(C[29]), .A2(n148), .B1(A[29]), .B2(n142), .ZN(n217) );
  AOI222_X1 U75 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n154), .ZN(n216) );
  NAND2_X1 U76 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI22_X1 U77 ( .A1(C[33]), .A2(n148), .B1(A[33]), .B2(n142), .ZN(n227) );
  AOI222_X1 U78 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n155), .ZN(n226) );
  NAND2_X1 U79 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  AOI22_X1 U80 ( .A1(C[16]), .A2(n149), .B1(A[16]), .B2(n143), .ZN(n189) );
  NAND2_X1 U81 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI222_X1 U82 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n155), .ZN(n234) );
  NAND2_X1 U83 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI222_X1 U84 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n155), .ZN(n244) );
  NAND2_X1 U85 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI22_X1 U86 ( .A1(C[38]), .A2(n147), .B1(A[38]), .B2(n141), .ZN(n237) );
  AOI222_X1 U87 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n155), .ZN(n236) );
  NAND2_X1 U88 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI22_X1 U89 ( .A1(C[18]), .A2(n149), .B1(A[18]), .B2(n143), .ZN(n193) );
  NAND2_X1 U90 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI22_X1 U91 ( .A1(C[26]), .A2(n148), .B1(A[26]), .B2(n142), .ZN(n211) );
  AOI222_X1 U92 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n154), .ZN(n210) );
  NAND2_X1 U93 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U94 ( .A1(C[30]), .A2(n148), .B1(A[30]), .B2(n142), .ZN(n221) );
  AOI222_X1 U95 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n154), .ZN(n220) );
  NAND2_X1 U96 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI22_X1 U97 ( .A1(C[34]), .A2(n148), .B1(A[34]), .B2(n142), .ZN(n229) );
  AOI222_X1 U98 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n155), .ZN(n228) );
  NAND2_X1 U99 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  AOI22_X1 U100 ( .A1(C[52]), .A2(n146), .B1(A[52]), .B2(n140), .ZN(n269) );
  AOI222_X1 U101 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n156), .ZN(n268) );
  NAND2_X1 U102 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI222_X1 U103 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n156), .ZN(n252) );
  NAND2_X1 U104 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI22_X1 U105 ( .A1(C[49]), .A2(n146), .B1(A[49]), .B2(n140), .ZN(n261) );
  AOI222_X1 U106 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n156), .ZN(n260) );
  NAND2_X1 U107 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI222_X1 U108 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n156), .ZN(n254) );
  AOI22_X1 U109 ( .A1(C[46]), .A2(n146), .B1(A[46]), .B2(n140), .ZN(n255) );
  NAND2_X1 U110 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI22_X1 U111 ( .A1(C[50]), .A2(n146), .B1(A[50]), .B2(n140), .ZN(n265) );
  AOI222_X1 U112 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n156), .ZN(n264) );
  NAND2_X1 U113 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  AOI22_X1 U114 ( .A1(C[51]), .A2(n146), .B1(A[51]), .B2(n140), .ZN(n267) );
  AOI222_X1 U115 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n156), .ZN(n266) );
  AOI22_X1 U116 ( .A1(C[24]), .A2(n149), .B1(A[24]), .B2(n143), .ZN(n207) );
  AOI222_X1 U117 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n154), .ZN(n206) );
  AOI22_X1 U118 ( .A1(C[28]), .A2(n148), .B1(A[28]), .B2(n142), .ZN(n215) );
  AOI222_X1 U119 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n154), .ZN(n214) );
  AOI22_X1 U120 ( .A1(C[32]), .A2(n148), .B1(A[32]), .B2(n142), .ZN(n225) );
  AOI222_X1 U121 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n155), .ZN(n224) );
  NAND2_X1 U122 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI222_X1 U123 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n155), .ZN(n246) );
  NAND2_X1 U124 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI222_X1 U125 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n155), .ZN(n230) );
  AOI22_X1 U126 ( .A1(C[35]), .A2(n148), .B1(A[35]), .B2(n142), .ZN(n231) );
  NAND2_X1 U127 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI222_X1 U128 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n155), .ZN(n238) );
  AOI22_X1 U129 ( .A1(C[39]), .A2(n147), .B1(A[39]), .B2(n141), .ZN(n239) );
  NAND2_X1 U130 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI22_X1 U131 ( .A1(C[25]), .A2(n148), .B1(A[25]), .B2(n142), .ZN(n209) );
  AOI222_X1 U132 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n154), .ZN(n208) );
  NAND2_X1 U133 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  AOI22_X1 U134 ( .A1(C[48]), .A2(n146), .B1(A[48]), .B2(n140), .ZN(n259) );
  AOI222_X1 U135 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n156), .ZN(n258) );
  NAND2_X1 U136 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI22_X1 U137 ( .A1(C[47]), .A2(n146), .B1(A[47]), .B2(n140), .ZN(n257) );
  AOI222_X1 U138 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n156), .ZN(n256) );
  AOI22_X1 U139 ( .A1(C[36]), .A2(n147), .B1(A[36]), .B2(n141), .ZN(n233) );
  AOI222_X1 U140 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n155), .ZN(n232) );
  AOI22_X1 U141 ( .A1(C[40]), .A2(n147), .B1(A[40]), .B2(n141), .ZN(n243) );
  AOI222_X1 U142 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n155), .ZN(n242) );
  AOI22_X1 U143 ( .A1(C[44]), .A2(n147), .B1(A[44]), .B2(n141), .ZN(n251) );
  AOI222_X1 U144 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n156), .ZN(n250) );
  NAND2_X1 U145 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  AOI22_X1 U146 ( .A1(C[20]), .A2(n149), .B1(A[20]), .B2(n143), .ZN(n199) );
  AOI222_X1 U147 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n154), .ZN(n198) );
  NAND2_X1 U148 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI222_X1 U149 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n155), .ZN(n248) );
  AOI22_X1 U150 ( .A1(C[43]), .A2(n147), .B1(A[43]), .B2(n141), .ZN(n249) );
  NAND2_X1 U151 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  AOI22_X1 U152 ( .A1(C[56]), .A2(n146), .B1(A[56]), .B2(n140), .ZN(n277) );
  AOI222_X1 U153 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n157), .ZN(n276) );
  NAND2_X1 U154 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U155 ( .A1(C[60]), .A2(n145), .B1(A[60]), .B2(n139), .ZN(n287) );
  AOI222_X1 U156 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n157), .ZN(n286) );
  NAND2_X1 U157 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  AOI22_X1 U158 ( .A1(C[57]), .A2(n145), .B1(A[57]), .B2(n139), .ZN(n279) );
  AOI222_X1 U159 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n157), .ZN(n278) );
  NAND2_X1 U160 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI22_X1 U161 ( .A1(C[58]), .A2(n145), .B1(A[58]), .B2(n139), .ZN(n281) );
  AOI222_X1 U162 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n157), .ZN(n280) );
  NAND2_X1 U163 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U164 ( .A1(C[59]), .A2(n145), .B1(A[59]), .B2(n139), .ZN(n283) );
  AOI222_X1 U165 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n157), .ZN(n282) );
  NAND2_X1 U166 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U167 ( .A1(C[61]), .A2(n145), .B1(A[61]), .B2(n139), .ZN(n289) );
  AOI222_X1 U168 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n157), .ZN(n288) );
  NAND2_X1 U169 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U170 ( .A1(C[62]), .A2(n145), .B1(A[62]), .B2(n139), .ZN(n291) );
  AOI222_X1 U171 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n157), .ZN(n290) );
  NAND2_X1 U172 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U173 ( .A1(C[63]), .A2(n145), .B1(A[63]), .B2(n139), .ZN(n293) );
  AOI222_X1 U174 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n157), .ZN(n292) );
  NAND2_X1 U175 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U176 ( .A1(C[0]), .A2(n145), .B1(A[0]), .B2(n139), .ZN(n175) );
  AOI222_X1 U177 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n153), .ZN(n174) );
  NAND2_X1 U178 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U179 ( .A1(C[4]), .A2(n146), .B1(A[4]), .B2(n140), .ZN(n263) );
  AOI222_X1 U180 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n156), .ZN(n262) );
  NAND2_X1 U181 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI22_X1 U182 ( .A1(C[8]), .A2(n145), .B1(A[8]), .B2(n139), .ZN(n299) );
  AOI222_X1 U183 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n157), .ZN(n298) );
  NAND2_X1 U184 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  AOI22_X1 U185 ( .A1(C[12]), .A2(n150), .B1(A[12]), .B2(n144), .ZN(n181) );
  AOI222_X1 U186 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n153), .ZN(n180) );
  NAND2_X1 U187 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U188 ( .A1(C[1]), .A2(n149), .B1(A[1]), .B2(n143), .ZN(n197) );
  AOI222_X1 U189 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n153), .ZN(n196) );
  NAND2_X1 U190 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U191 ( .A1(C[5]), .A2(n145), .B1(A[5]), .B2(n139), .ZN(n285) );
  AOI222_X1 U192 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n157), .ZN(n284) );
  NAND2_X1 U193 ( .A1(n306), .A2(n305), .ZN(Y[9]) );
  AOI22_X1 U194 ( .A1(C[9]), .A2(n147), .B1(A[9]), .B2(n141), .ZN(n306) );
  AOI222_X1 U195 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n157), .ZN(n305) );
  NAND2_X1 U196 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U197 ( .A1(C[13]), .A2(n150), .B1(A[13]), .B2(n144), .ZN(n183) );
  AOI222_X1 U198 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n153), .ZN(n182) );
  NAND2_X1 U199 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U200 ( .A1(C[2]), .A2(n148), .B1(A[2]), .B2(n142), .ZN(n219) );
  AOI222_X1 U201 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n154), .ZN(n218) );
  NAND2_X1 U202 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U203 ( .A1(C[6]), .A2(n145), .B1(A[6]), .B2(n139), .ZN(n295) );
  AOI222_X1 U204 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n157), .ZN(n294) );
  NAND2_X1 U205 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U206 ( .A1(C[10]), .A2(n150), .B1(A[10]), .B2(n144), .ZN(n177) );
  AOI222_X1 U207 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n153), .ZN(n176) );
  NAND2_X1 U208 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U209 ( .A1(C[3]), .A2(n147), .B1(A[3]), .B2(n141), .ZN(n241) );
  AOI222_X1 U210 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n155), .ZN(n240) );
  NAND2_X1 U211 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U212 ( .A1(C[7]), .A2(n145), .B1(A[7]), .B2(n139), .ZN(n297) );
  AOI222_X1 U213 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n157), .ZN(n296) );
  NAND2_X1 U214 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U215 ( .A1(C[11]), .A2(n150), .B1(A[11]), .B2(n144), .ZN(n179) );
  AOI222_X1 U216 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n153), .ZN(n178) );
  AOI22_X1 U217 ( .A1(C[42]), .A2(n147), .B1(A[42]), .B2(n141), .ZN(n247) );
  AOI22_X1 U218 ( .A1(C[41]), .A2(n147), .B1(A[41]), .B2(n141), .ZN(n245) );
  AOI22_X1 U219 ( .A1(C[14]), .A2(n149), .B1(A[14]), .B2(n143), .ZN(n185) );
  AOI22_X1 U220 ( .A1(C[15]), .A2(n149), .B1(A[15]), .B2(n143), .ZN(n187) );
  NAND2_X1 U221 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  NAND2_X1 U222 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI222_X1 U223 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n153), .ZN(n194) );
  AOI222_X1 U224 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n153), .ZN(n192) );
  AOI22_X1 U225 ( .A1(C[37]), .A2(n147), .B1(A[37]), .B2(n141), .ZN(n235) );
  AOI222_X1 U226 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n153), .ZN(n186) );
  AOI22_X1 U227 ( .A1(C[45]), .A2(n147), .B1(A[45]), .B2(n141), .ZN(n253) );
  AOI222_X1 U228 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n153), .ZN(n190) );
  AOI222_X1 U229 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n153), .ZN(n188) );
  CLKBUF_X1 U230 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U231 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U232 ( .A(n158), .Z(n164) );
endmodule


module G_153 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_567 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_566 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_565 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_564 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_563 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_562 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_561 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_560 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_559 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_558 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_557 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_556 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_555 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_554 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_553 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_552 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_551 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_550 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_549 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_548 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_547 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_546 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_545 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_544 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_543 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_542 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_541 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_540 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_539 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_538 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_537 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_152 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_536 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_535 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_534 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3, n5;

  AND2_X1 U1 ( .A1(P_IK), .A2(G_K_1), .ZN(n3) );
  NOR2_X1 U2 ( .A1(n3), .A2(G_IK), .ZN(n5) );
  INV_X1 U3 ( .A(n5), .ZN(Gx) );
  AND2_X1 U4 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_533 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_532 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_531 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_530 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_529 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_528 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_527 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_526 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_525 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_524 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_523 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_522 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_151 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_521 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_520 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_519 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_518 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_517 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_516 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_515 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_150 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_149 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_514 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_513 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_512 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  OR2_X1 U2 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_511 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_510 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_509 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_148 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_147 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_146 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_145 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_508 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_507 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_506 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_505 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_144 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_143 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_142 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_141 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_140 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_139 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_138 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_137 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module carry_generator_N64_NPB4_9 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U77 ( .A(B[59]), .B(A[59]), .Z(\PG_Network[0][0][59] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U81 ( .A(B[55]), .B(A[55]), .Z(\PG_Network[0][0][55] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U85 ( .A(B[51]), .B(A[51]), .Z(\PG_Network[0][0][51] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U88 ( .A(B[49]), .B(A[49]), .Z(\PG_Network[0][0][49] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U91 ( .A(B[46]), .B(A[46]), .Z(\PG_Network[0][0][46] ) );
  XOR2_X1 U92 ( .A(B[45]), .B(A[45]), .Z(\PG_Network[0][0][45] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U101 ( .A(B[37]), .B(A[37]), .Z(\PG_Network[0][0][37] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U125 ( .A(B[15]), .B(A[15]), .Z(\PG_Network[0][0][15] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_153 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n25), .Gx(\PG_Network[1][1][1] ) );
  PG_567 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_566 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_565 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_564 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_563 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_562 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_561 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_560 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_559 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_558 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_557 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_556 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_555 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_554 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_553 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_552 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_551 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_550 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_549 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_548 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_547 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_546 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_545 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_544 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_543 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_542 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_541 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_540 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_539 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_538 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_537 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_152 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_536 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_535 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_534 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_533 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_532 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_531 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_530 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_529 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_528 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_527 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_526 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_525 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_524 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_523 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_522 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_151 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_521 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_520 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_519 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_518 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_517 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_516 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(n6), .P_K_1(\PG_Network[2][0][51] ), 
        .Gx(\PG_Network[3][1][55] ), .Px(\PG_Network[3][0][55] ) );
  PG_515 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_150 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), .G_K_1(Co[1]), .Gx(Co[3]) );
  G_149 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_514 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_513 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_512 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(n17), 
        .Gx(\PG_Network[4][1][47] ), .Px(\PG_Network[4][0][47] ) );
  PG_511 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(n17), 
        .Gx(\PG_Network[4][1][43] ), .Px(\PG_Network[4][0][43] ) );
  PG_510 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][63] ), .Px(
        \PG_Network[4][0][63] ) );
  PG_509 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][59] ), .Px(
        \PG_Network[4][0][59] ) );
  G_148 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), .G_K_1(n5), .Gx(Co[7]) );
  G_147 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), .G_K_1(n5), .Gx(Co[6]) );
  G_146 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), .G_K_1(n5), .Gx(Co[5]) );
  G_145 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), .G_K_1(Co[3]), .Gx(Co[4]) );
  PG_508 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(n23), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][63] ), .Px(\PG_Network[5][0][63] ) );
  PG_507 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(n23), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][59] ), .Px(\PG_Network[5][0][59] ) );
  PG_506 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(n23), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][55] ), .Px(\PG_Network[5][0][55] ) );
  PG_505 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(n23), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][51] ), .Px(\PG_Network[5][0][51] ) );
  G_144 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), .G_K_1(n15), .Gx(Co[15]) );
  G_143 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), .G_K_1(n15), .Gx(Co[14]) );
  G_142 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), .G_K_1(n15), .Gx(Co[13]) );
  G_141 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), .G_K_1(Co[7]), .Gx(Co[12]) );
  G_140 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), .G_K_1(Co[7]), .Gx(Co[11]) );
  G_139 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), .G_K_1(Co[7]), .Gx(Co[10]) );
  G_138 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), .G_K_1(Co[7]), .Gx(Co[9]) );
  G_137 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), .G_K_1(Co[7]), .Gx(Co[8]) );
  CLKBUF_X1 U1 ( .A(Co[3]), .Z(n5) );
  BUF_X1 U2 ( .A(\PG_Network[3][0][39] ), .Z(n17) );
  CLKBUF_X1 U3 ( .A(\PG_Network[2][1][51] ), .Z(n6) );
  INV_X1 U4 ( .A(A[19]), .ZN(n8) );
  INV_X1 U5 ( .A(A[30]), .ZN(n7) );
  INV_X1 U6 ( .A(A[23]), .ZN(n21) );
  INV_X1 U7 ( .A(A[31]), .ZN(n19) );
  INV_X1 U8 ( .A(A[39]), .ZN(n14) );
  INV_X1 U9 ( .A(A[47]), .ZN(n24) );
  INV_X1 U10 ( .A(A[43]), .ZN(n22) );
  INV_X1 U11 ( .A(A[25]), .ZN(n18) );
  INV_X1 U12 ( .A(A[29]), .ZN(n9) );
  INV_X1 U13 ( .A(A[27]), .ZN(n20) );
  INV_X1 U14 ( .A(A[38]), .ZN(n10) );
  XNOR2_X1 U15 ( .A(B[30]), .B(n7), .ZN(\PG_Network[0][0][30] ) );
  XNOR2_X1 U16 ( .A(B[19]), .B(n8), .ZN(\PG_Network[0][0][19] ) );
  XNOR2_X1 U17 ( .A(B[29]), .B(n9), .ZN(\PG_Network[0][0][29] ) );
  XNOR2_X1 U18 ( .A(B[38]), .B(n10), .ZN(\PG_Network[0][0][38] ) );
  NAND2_X1 U19 ( .A1(B[35]), .A2(n16), .ZN(n12) );
  NAND2_X1 U20 ( .A1(n11), .A2(A[35]), .ZN(n13) );
  NAND2_X1 U21 ( .A1(n12), .A2(n13), .ZN(\PG_Network[0][0][35] ) );
  INV_X1 U22 ( .A(B[35]), .ZN(n11) );
  INV_X1 U23 ( .A(A[35]), .ZN(n16) );
  XNOR2_X1 U24 ( .A(B[39]), .B(n14), .ZN(\PG_Network[0][0][39] ) );
  CLKBUF_X1 U25 ( .A(Co[7]), .Z(n15) );
  XNOR2_X1 U26 ( .A(B[25]), .B(n18), .ZN(\PG_Network[0][0][25] ) );
  XNOR2_X1 U27 ( .A(B[31]), .B(n19), .ZN(\PG_Network[0][0][31] ) );
  XNOR2_X1 U28 ( .A(B[27]), .B(n20), .ZN(\PG_Network[0][0][27] ) );
  XNOR2_X1 U29 ( .A(B[23]), .B(n21), .ZN(\PG_Network[0][0][23] ) );
  XNOR2_X1 U30 ( .A(B[43]), .B(n22), .ZN(\PG_Network[0][0][43] ) );
  CLKBUF_X1 U31 ( .A(\PG_Network[4][1][47] ), .Z(n23) );
  XNOR2_X1 U32 ( .A(B[47]), .B(n24), .ZN(\PG_Network[0][0][47] ) );
  AND2_X1 U33 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U34 ( .A1(B[27]), .A2(A[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U35 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U36 ( .A1(B[35]), .A2(A[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U37 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U38 ( .A1(A[51]), .A2(B[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U39 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U40 ( .A1(B[46]), .A2(A[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U41 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U42 ( .A1(B[25]), .A2(A[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U43 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U44 ( .A1(A[19]), .A2(B[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U45 ( .A1(A[21]), .A2(B[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U46 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U47 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U48 ( .A1(A[41]), .A2(B[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U49 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U50 ( .A1(B[31]), .A2(A[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U51 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U52 ( .A1(A[15]), .A2(B[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U53 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U54 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U55 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U56 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U57 ( .A1(A[45]), .A2(B[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U58 ( .A1(A[49]), .A2(B[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U59 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U60 ( .A1(A[55]), .A2(B[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U61 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U62 ( .A1(A[59]), .A2(B[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U63 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U64 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
  AND2_X1 U65 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U66 ( .A1(B[29]), .A2(A[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U67 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U90 ( .A1(A[53]), .A2(B[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U94 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AND2_X1 U99 ( .A1(B[23]), .A2(A[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U100 ( .A1(A[37]), .A2(B[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U103 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U107 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U108 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U110 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U112 ( .A1(A[11]), .A2(B[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U114 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U116 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U121 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U131 ( .A(n28), .ZN(n25) );
  AND2_X1 U132 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U133 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U134 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AND2_X1 U135 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U136 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U137 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U138 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U139 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U140 ( .A1(A[7]), .A2(B[7]), .ZN(\PG_Network[0][1][7] ) );
  AOI21_X1 U141 ( .B1(A[0]), .B2(B[0]), .A(n26), .ZN(n28) );
  INV_X1 U142 ( .A(n27), .ZN(n26) );
  OAI21_X1 U143 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n27) );
  AND2_X1 U144 ( .A1(B[47]), .A2(A[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U145 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U146 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U147 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U148 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U149 ( .A1(B[43]), .A2(A[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U150 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
endmodule


module FA_1152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_288 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1152 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1151 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1150 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1149 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1148 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1147 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1146 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1145 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_287 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1148 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1147 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1146 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1145 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_144 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U2 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_144 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_288 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_287 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_144 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_286 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1144 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1143 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1142 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1141 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1140 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1139 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1138 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1137 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_285 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1140 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1139 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1138 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1137 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_143 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_143 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_286 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_285 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_143 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_284 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1136 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1135 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1134 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1133 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1132 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1131 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1130 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1129 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_283 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1132 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1131 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1130 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1129 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_142 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_142 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_284 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_283 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_142 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_282 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1128 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1127 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1126 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1125 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1123 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1122 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1121 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_281 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1124 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1123 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1122 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1121 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_141 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_141 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_282 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_281 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_141 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_280 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1120 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1119 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1118 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1117 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_279 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1116 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1115 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1114 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1113 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_140 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(sel), .ZN(n13) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
endmodule


module carry_select_block_NPB4_140 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_280 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_279 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_140 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n5), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_278 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1112 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1111 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1110 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1109 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_277 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1108 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1107 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1106 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1105 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_139 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n18), .ZN(Y[2]) );
  BUF_X1 U3 ( .A(n15), .Z(n5) );
  CLKBUF_X1 U4 ( .A(sel), .Z(n10) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U6 ( .A(sel), .ZN(n15) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U11 ( .A(n19), .ZN(Y[3]) );
endmodule


module carry_select_block_NPB4_139 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_278 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_277 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_139 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(n5), .B(B), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_1102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_276 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1104 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1103 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1102 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1101 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1099 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1098 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1097 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_275 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1100 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1099 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1098 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1097 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_138 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19, n20;

  INV_X1 U1 ( .A(n17), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n20), .ZN(Y[3]) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n11) );
  CLKBUF_X1 U4 ( .A(n5), .Z(n10) );
  INV_X1 U5 ( .A(sel), .ZN(n5) );
  INV_X1 U6 ( .A(n19), .ZN(Y[2]) );
  INV_X1 U7 ( .A(n18), .ZN(Y[1]) );
  INV_X1 U8 ( .A(sel), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n11), .B1(B[3]), .B2(n10), .ZN(n20) );
  AOI22_X1 U10 ( .A1(A[2]), .A2(n11), .B1(B[2]), .B2(n10), .ZN(n19) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n5), .ZN(n18) );
  AOI22_X1 U12 ( .A1(sel), .A2(A[0]), .B1(n16), .B2(B[0]), .ZN(n17) );
endmodule


module carry_select_block_NPB4_138 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_276 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_275 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_138 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1096 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1095 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68719, n4, n5, n6;
  assign Co = net68719;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n6) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  OAI21_X1 U5 ( .B1(n4), .B2(n5), .A(n6), .ZN(net68719) );
endmodule


module FA_1094 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_1093 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_274 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1096 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1095 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1094 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1093 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1092 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1091 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1090 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1089 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_273 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1092 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1091 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1090 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1089 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_137 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U2 ( .A(n17), .ZN(Y[1]) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n5) );
  INV_X1 U4 ( .A(sel), .ZN(n10) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[2]), .B1(n15), .B2(B[2]), .ZN(n18) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[1]), .B1(n10), .B2(B[1]), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n15), .ZN(n19) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n10), .B2(B[0]), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_137 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_274 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_273 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_137 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1088 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_1087 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1086 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1085 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_272 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1088 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1087 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1086 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1085 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1084 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1083 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1082 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1081 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_271 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1084 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1083 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1082 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1081 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_136 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n16), .ZN(Y[1]) );
  BUF_X1 U2 ( .A(n14), .Z(n5) );
  INV_X1 U3 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U4 ( .A(sel), .ZN(n14) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U6 ( .A(n17), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n17) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n5), .ZN(n18) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
endmodule


module carry_select_block_NPB4_136 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_272 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_271 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_136 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1080 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_1079 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1078 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68702, n4, n5, n6;
  assign Co = net68702;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n6) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  OAI21_X1 U5 ( .B1(n5), .B2(n4), .A(n6), .ZN(net68702) );
endmodule


module FA_1077 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(n4), .ZN(n7) );
endmodule


module RCA_N4_270 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1080 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1079 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1078 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1077 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1076 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1075 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1074 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1073 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_269 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1076 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1075 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1074 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1073 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_135 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(sel), .Z(n11) );
  INV_X1 U2 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U4 ( .A(sel), .ZN(n5) );
  INV_X1 U5 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U6 ( .A(n11), .ZN(n10) );
  INV_X1 U7 ( .A(n16), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n11), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U9 ( .A1(n11), .A2(A[1]), .B1(n5), .B2(B[1]), .ZN(n17) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n5), .B2(B[0]), .ZN(n16) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n11), .B1(B[3]), .B2(n10), .ZN(n19) );
endmodule


module carry_select_block_NPB4_135 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_270 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_269 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_135 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1072 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n4), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_1071 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1070 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1069 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_268 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1072 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1071 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1070 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1069 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1068 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1067 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1066 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1065 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_267 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1068 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1067 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1066 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1065 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_134 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n10), .ZN(n5) );
  BUF_X2 U3 ( .A(sel), .Z(n10) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U6 ( .A(sel), .ZN(n15) );
  AOI22_X1 U7 ( .A1(n10), .A2(A[1]), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U10 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U11 ( .A1(n10), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n19) );
endmodule


module carry_select_block_NPB4_134 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_268 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_267 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_134 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1064 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8, n9;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n5) );
  CLKBUF_X1 U2 ( .A(n9), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n8), .A2(n7), .ZN(Co) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(n7) );
  NAND2_X1 U7 ( .A1(n9), .A2(Ci), .ZN(n8) );
endmodule


module FA_1063 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1062 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_1061 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_266 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1064 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1063 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1062 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1061 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1060 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1059 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1058 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1057 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_265 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1060 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1059 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1058 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1057 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_133 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(sel), .ZN(n10) );
  INV_X1 U3 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  AOI22_X1 U6 ( .A1(n5), .A2(A[2]), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n10), .ZN(n17) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
  INV_X1 U9 ( .A(sel), .ZN(n15) );
  INV_X1 U10 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n10), .ZN(n19) );
endmodule


module carry_select_block_NPB4_133 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_266 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_265 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_133 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1056 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_1055 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1054 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1053 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(n4), .ZN(n7) );
endmodule


module RCA_N4_264 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1056 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1055 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1054 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1053 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1052 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1051 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1050 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1049 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_263 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1052 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1051 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1050 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1049 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_132 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19, n20;

  BUF_X1 U1 ( .A(n16), .Z(n10) );
  BUF_X1 U2 ( .A(n11), .Z(n5) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n11) );
  INV_X2 U4 ( .A(n17), .ZN(Y[0]) );
  INV_X1 U5 ( .A(n20), .ZN(Y[3]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[2]) );
  INV_X1 U7 ( .A(n18), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n10), .ZN(n19) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(n11), .B1(B[1]), .B2(n16), .ZN(n18) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n10), .ZN(n20) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n16), .ZN(n17) );
  INV_X1 U12 ( .A(sel), .ZN(n16) );
endmodule


module carry_select_block_NPB4_132 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_264 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_263 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_132 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1048 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1047 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1046 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1045 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_262 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1048 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1047 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1046 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1045 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1044 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1043 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1042 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1041 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_261 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1044 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1043 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1042 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1041 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_131 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  BUF_X1 U1 ( .A(n14), .Z(n5) );
  INV_X1 U2 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n17) );
  INV_X1 U6 ( .A(n16), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n18) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
  INV_X1 U10 ( .A(sel), .ZN(n14) );
endmodule


module carry_select_block_NPB4_131 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_262 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_261 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_131 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1040 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1039 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1038 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1037 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_260 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1040 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1039 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1038 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1037 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1036 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1035 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1034 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1033 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_259 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1036 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1035 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1034 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1033 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_130 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_130 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_260 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_259 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_130 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1032 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1031 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1030 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1029 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_258 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1032 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1031 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1030 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1029 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1028 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1027 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1026 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1025 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_257 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1028 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1027 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1026 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1025 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_129 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_129 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_258 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_257 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_129 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_9 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_144 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_143 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_142 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_141 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_140 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_139 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_138 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_137 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_136 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_135 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_134 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), .S(S[43:40]) );
  carry_select_block_NPB4_133 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), .S(S[47:44]) );
  carry_select_block_NPB4_132 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), .S(S[51:48]) );
  carry_select_block_NPB4_131 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), .S(S[55:52]) );
  carry_select_block_NPB4_130 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), .S(S[59:56]) );
  carry_select_block_NPB4_129 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), .S(S[63:60]) );
endmodule


module P4_ADDER_N64_9 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_9 CGEN ( .A(A), .B({B[63:49], n4, B[47:45], n18, 
        B[43:41], n17, B[39:33], n1, B[31:21], n19, B[19:0]}), .Cin(Cin), .Co(
        CoutCgen) );
  sum_generator_N64_NPB4_9 SGEN ( .A(A), .B({B[63:48], n10, B[46:44], n3, 
        B[42:40], n14, n13, n6, B[36], n5, B[34:32], n7, n9, B[29:28], n11, 
        B[26:24], n2, B[22:20], n16, B[18:0]}), .Ci({CoutCgen, Cin}), .S(S), 
        .Co(Cout) );
  BUF_X2 U1 ( .A(B[37]), .Z(n6) );
  CLKBUF_X1 U2 ( .A(B[32]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(B[23]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(B[43]), .Z(n3) );
  CLKBUF_X1 U5 ( .A(B[48]), .Z(n4) );
  CLKBUF_X1 U6 ( .A(B[35]), .Z(n5) );
  CLKBUF_X1 U7 ( .A(B[31]), .Z(n7) );
  INV_X1 U8 ( .A(B[30]), .ZN(n8) );
  INV_X1 U9 ( .A(n8), .ZN(n9) );
  CLKBUF_X1 U10 ( .A(B[47]), .Z(n10) );
  CLKBUF_X1 U11 ( .A(B[27]), .Z(n11) );
  INV_X1 U12 ( .A(B[38]), .ZN(n12) );
  INV_X1 U13 ( .A(n12), .ZN(n13) );
  CLKBUF_X1 U14 ( .A(B[39]), .Z(n14) );
  INV_X1 U15 ( .A(B[19]), .ZN(n15) );
  INV_X1 U16 ( .A(n15), .ZN(n16) );
  CLKBUF_X1 U17 ( .A(B[40]), .Z(n17) );
  CLKBUF_X1 U18 ( .A(B[20]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(B[44]), .Z(n18) );
endmodule


module Booth_Encoder_8 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_8 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306;

  NAND2_X1 U1 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  NAND2_X1 U2 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  NAND2_X1 U3 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  NAND2_X1 U4 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  NAND2_X1 U5 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  NAND2_X1 U6 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  NAND2_X2 U7 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  NOR3_X1 U8 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U9 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  BUF_X1 U10 ( .A(n158), .Z(n161) );
  BUF_X1 U11 ( .A(n158), .Z(n160) );
  BUF_X1 U12 ( .A(n158), .Z(n159) );
  BUF_X1 U13 ( .A(n158), .Z(n162) );
  BUF_X1 U14 ( .A(n158), .Z(n163) );
  BUF_X1 U15 ( .A(n151), .Z(n154) );
  BUF_X1 U16 ( .A(n165), .Z(n168) );
  BUF_X1 U17 ( .A(n151), .Z(n153) );
  BUF_X1 U18 ( .A(n165), .Z(n167) );
  BUF_X1 U19 ( .A(n303), .Z(n158) );
  NOR4_X1 U20 ( .A1(n150), .A2(n144), .A3(n153), .A4(n167), .ZN(n303) );
  BUF_X1 U21 ( .A(n151), .Z(n155) );
  BUF_X1 U22 ( .A(n152), .Z(n156) );
  BUF_X1 U23 ( .A(n165), .Z(n169) );
  BUF_X1 U24 ( .A(n166), .Z(n170) );
  BUF_X1 U25 ( .A(n152), .Z(n157) );
  BUF_X1 U26 ( .A(n166), .Z(n171) );
  BUF_X1 U27 ( .A(n301), .Z(n149) );
  BUF_X1 U28 ( .A(n304), .Z(n165) );
  BUF_X1 U29 ( .A(n302), .Z(n151) );
  BUF_X1 U30 ( .A(n301), .Z(n148) );
  BUF_X1 U31 ( .A(n301), .Z(n146) );
  BUF_X1 U32 ( .A(n301), .Z(n147) );
  BUF_X1 U33 ( .A(n304), .Z(n166) );
  BUF_X1 U34 ( .A(n302), .Z(n152) );
  BUF_X1 U35 ( .A(n301), .Z(n145) );
  BUF_X1 U36 ( .A(n300), .Z(n142) );
  BUF_X1 U37 ( .A(n300), .Z(n139) );
  BUF_X1 U38 ( .A(n300), .Z(n140) );
  BUF_X1 U39 ( .A(n300), .Z(n143) );
  BUF_X1 U40 ( .A(n300), .Z(n141) );
  INV_X1 U41 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U42 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n304) );
  AND3_X1 U43 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U44 ( .A(sel[2]), .ZN(n173) );
  AOI22_X1 U45 ( .A1(C[24]), .A2(n149), .B1(A[24]), .B2(n143), .ZN(n207) );
  AOI222_X1 U46 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n154), .ZN(n206) );
  AOI22_X1 U47 ( .A1(C[28]), .A2(n148), .B1(A[28]), .B2(n142), .ZN(n215) );
  AOI222_X1 U48 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n154), .ZN(n214) );
  NAND2_X1 U49 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI22_X1 U50 ( .A1(C[25]), .A2(n148), .B1(A[25]), .B2(n142), .ZN(n209) );
  AOI222_X1 U51 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n154), .ZN(n208) );
  NAND2_X1 U52 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI22_X1 U53 ( .A1(C[22]), .A2(n149), .B1(A[22]), .B2(n143), .ZN(n203) );
  AOI222_X1 U54 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n154), .ZN(n202) );
  NAND2_X1 U55 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI22_X1 U56 ( .A1(C[26]), .A2(n148), .B1(A[26]), .B2(n142), .ZN(n211) );
  AOI222_X1 U57 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n154), .ZN(n210) );
  NAND2_X1 U58 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U59 ( .A1(C[30]), .A2(n148), .B1(A[30]), .B2(n142), .ZN(n221) );
  AOI222_X1 U60 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n154), .ZN(n220) );
  NAND2_X1 U61 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI22_X1 U62 ( .A1(C[23]), .A2(n149), .B1(A[23]), .B2(n143), .ZN(n205) );
  AOI222_X1 U63 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n154), .ZN(n204) );
  AOI222_X1 U64 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n153), .ZN(n188) );
  NAND2_X1 U65 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI22_X1 U66 ( .A1(C[18]), .A2(n149), .B1(A[18]), .B2(n143), .ZN(n193) );
  NAND2_X1 U67 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI22_X1 U68 ( .A1(C[19]), .A2(n149), .B1(A[19]), .B2(n143), .ZN(n195) );
  NAND2_X1 U69 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI22_X1 U70 ( .A1(C[21]), .A2(n149), .B1(A[21]), .B2(n143), .ZN(n201) );
  NAND2_X1 U71 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI22_X1 U72 ( .A1(C[34]), .A2(n148), .B1(A[34]), .B2(n142), .ZN(n229) );
  AOI222_X1 U73 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n155), .ZN(n228) );
  NAND2_X1 U74 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI22_X1 U75 ( .A1(C[27]), .A2(n148), .B1(A[27]), .B2(n142), .ZN(n213) );
  AOI222_X1 U76 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n154), .ZN(n212) );
  NAND2_X1 U77 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI22_X1 U78 ( .A1(C[35]), .A2(n148), .B1(A[35]), .B2(n142), .ZN(n231) );
  AOI222_X1 U79 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n155), .ZN(n230) );
  NAND2_X1 U80 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  AOI22_X1 U81 ( .A1(C[20]), .A2(n149), .B1(A[20]), .B2(n143), .ZN(n199) );
  AOI22_X1 U82 ( .A1(C[32]), .A2(n148), .B1(A[32]), .B2(n142), .ZN(n225) );
  AOI222_X1 U83 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n155), .ZN(n224) );
  NAND2_X1 U84 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI22_X1 U85 ( .A1(C[49]), .A2(n146), .B1(A[49]), .B2(n140), .ZN(n261) );
  AOI222_X1 U86 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n156), .ZN(n260) );
  NAND2_X1 U87 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI22_X1 U88 ( .A1(C[50]), .A2(n146), .B1(A[50]), .B2(n140), .ZN(n265) );
  AOI222_X1 U89 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n156), .ZN(n264) );
  NAND2_X1 U90 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  AOI22_X1 U91 ( .A1(C[51]), .A2(n146), .B1(A[51]), .B2(n140), .ZN(n267) );
  AOI222_X1 U92 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n156), .ZN(n266) );
  NAND2_X1 U93 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI22_X1 U94 ( .A1(C[38]), .A2(n147), .B1(A[38]), .B2(n141), .ZN(n237) );
  AOI222_X1 U95 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n155), .ZN(n236) );
  NAND2_X1 U96 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI22_X1 U97 ( .A1(C[42]), .A2(n147), .B1(A[42]), .B2(n141), .ZN(n247) );
  AOI222_X1 U98 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n155), .ZN(n246) );
  NAND2_X1 U99 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI22_X1 U100 ( .A1(C[46]), .A2(n146), .B1(A[46]), .B2(n140), .ZN(n255) );
  AOI222_X1 U101 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n156), .ZN(n254) );
  NAND2_X1 U102 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI222_X1 U103 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n154), .ZN(n216) );
  AOI22_X1 U104 ( .A1(C[29]), .A2(n148), .B1(A[29]), .B2(n142), .ZN(n217) );
  NAND2_X1 U105 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI222_X1 U106 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n155), .ZN(n226) );
  AOI22_X1 U107 ( .A1(C[33]), .A2(n148), .B1(A[33]), .B2(n142), .ZN(n227) );
  NAND2_X1 U108 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI222_X1 U109 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n155), .ZN(n234) );
  AOI22_X1 U110 ( .A1(C[37]), .A2(n147), .B1(A[37]), .B2(n141), .ZN(n235) );
  NAND2_X1 U111 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI222_X1 U112 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n155), .ZN(n244) );
  AOI22_X1 U113 ( .A1(C[41]), .A2(n147), .B1(A[41]), .B2(n141), .ZN(n245) );
  NAND2_X1 U114 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI222_X1 U115 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n156), .ZN(n252) );
  AOI22_X1 U116 ( .A1(C[45]), .A2(n147), .B1(A[45]), .B2(n141), .ZN(n253) );
  AOI22_X1 U117 ( .A1(C[40]), .A2(n147), .B1(A[40]), .B2(n141), .ZN(n243) );
  AOI222_X1 U118 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n155), .ZN(n242) );
  NAND2_X1 U119 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI222_X1 U120 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n155), .ZN(n238) );
  NAND2_X1 U121 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI222_X1 U122 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n155), .ZN(n248) );
  NAND2_X1 U123 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI222_X1 U124 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n156), .ZN(n256) );
  AOI22_X1 U125 ( .A1(C[36]), .A2(n147), .B1(A[36]), .B2(n141), .ZN(n233) );
  AOI222_X1 U126 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n155), .ZN(n232) );
  AOI222_X1 U127 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n156), .ZN(n258) );
  AOI22_X1 U128 ( .A1(C[48]), .A2(n146), .B1(A[48]), .B2(n140), .ZN(n259) );
  AOI222_X1 U129 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n156), .ZN(n250) );
  NAND2_X1 U130 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI22_X1 U131 ( .A1(C[31]), .A2(n148), .B1(A[31]), .B2(n142), .ZN(n223) );
  AOI222_X1 U132 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n154), .ZN(n222) );
  NAND2_X1 U133 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  AOI22_X1 U134 ( .A1(C[56]), .A2(n146), .B1(A[56]), .B2(n140), .ZN(n277) );
  AOI222_X1 U135 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n157), .ZN(n276) );
  NAND2_X1 U136 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  AOI22_X1 U137 ( .A1(C[53]), .A2(n146), .B1(A[53]), .B2(n140), .ZN(n271) );
  AOI222_X1 U138 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n156), .ZN(n270) );
  NAND2_X1 U139 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  AOI22_X1 U140 ( .A1(C[57]), .A2(n145), .B1(A[57]), .B2(n139), .ZN(n279) );
  AOI222_X1 U141 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n157), .ZN(n278) );
  NAND2_X1 U142 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI22_X1 U143 ( .A1(C[54]), .A2(n146), .B1(A[54]), .B2(n140), .ZN(n273) );
  AOI222_X1 U144 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n156), .ZN(n272) );
  NAND2_X1 U145 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI22_X1 U146 ( .A1(C[58]), .A2(n145), .B1(A[58]), .B2(n139), .ZN(n281) );
  AOI222_X1 U147 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n157), .ZN(n280) );
  NAND2_X1 U148 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI22_X1 U149 ( .A1(C[55]), .A2(n146), .B1(A[55]), .B2(n140), .ZN(n275) );
  AOI222_X1 U150 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n156), .ZN(n274) );
  NAND2_X1 U151 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U152 ( .A1(C[59]), .A2(n145), .B1(A[59]), .B2(n139), .ZN(n283) );
  AOI222_X1 U153 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n157), .ZN(n282) );
  NAND2_X1 U154 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  AOI22_X1 U155 ( .A1(C[52]), .A2(n146), .B1(A[52]), .B2(n140), .ZN(n269) );
  AOI222_X1 U156 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n156), .ZN(n268) );
  NAND2_X1 U157 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U158 ( .A1(C[60]), .A2(n145), .B1(A[60]), .B2(n139), .ZN(n287) );
  AOI222_X1 U159 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n157), .ZN(n286) );
  NAND2_X1 U160 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U161 ( .A1(C[61]), .A2(n145), .B1(A[61]), .B2(n139), .ZN(n289) );
  AOI222_X1 U162 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n157), .ZN(n288) );
  NAND2_X1 U163 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U164 ( .A1(C[62]), .A2(n145), .B1(A[62]), .B2(n139), .ZN(n291) );
  AOI222_X1 U165 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n157), .ZN(n290) );
  NAND2_X1 U166 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U167 ( .A1(C[63]), .A2(n145), .B1(A[63]), .B2(n139), .ZN(n293) );
  AOI222_X1 U168 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n157), .ZN(n292) );
  NAND2_X1 U169 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U170 ( .A1(C[0]), .A2(n145), .B1(A[0]), .B2(n139), .ZN(n175) );
  AOI222_X1 U171 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n153), .ZN(n174) );
  NAND2_X1 U172 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U173 ( .A1(C[4]), .A2(n146), .B1(A[4]), .B2(n140), .ZN(n263) );
  AOI222_X1 U174 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n156), .ZN(n262) );
  NAND2_X1 U175 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI22_X1 U176 ( .A1(C[8]), .A2(n145), .B1(A[8]), .B2(n139), .ZN(n299) );
  AOI222_X1 U177 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n157), .ZN(n298) );
  NAND2_X1 U178 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  AOI22_X1 U179 ( .A1(C[12]), .A2(n150), .B1(A[12]), .B2(n144), .ZN(n181) );
  AOI222_X1 U180 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n153), .ZN(n180) );
  NAND2_X1 U181 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U182 ( .A1(C[1]), .A2(n149), .B1(A[1]), .B2(n143), .ZN(n197) );
  AOI222_X1 U183 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n153), .ZN(n196) );
  NAND2_X1 U184 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U185 ( .A1(C[5]), .A2(n145), .B1(A[5]), .B2(n139), .ZN(n285) );
  AOI222_X1 U186 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n157), .ZN(n284) );
  NAND2_X1 U187 ( .A1(n306), .A2(n305), .ZN(Y[9]) );
  AOI22_X1 U188 ( .A1(C[9]), .A2(n147), .B1(A[9]), .B2(n141), .ZN(n306) );
  AOI222_X1 U189 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n157), .ZN(n305) );
  NAND2_X1 U190 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U191 ( .A1(C[13]), .A2(n150), .B1(A[13]), .B2(n144), .ZN(n183) );
  AOI222_X1 U192 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n153), .ZN(n182) );
  NAND2_X1 U193 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U194 ( .A1(C[2]), .A2(n148), .B1(A[2]), .B2(n142), .ZN(n219) );
  AOI222_X1 U195 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n154), .ZN(n218) );
  NAND2_X1 U196 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U197 ( .A1(C[6]), .A2(n145), .B1(A[6]), .B2(n139), .ZN(n295) );
  AOI222_X1 U198 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n157), .ZN(n294) );
  NAND2_X1 U199 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U200 ( .A1(C[10]), .A2(n150), .B1(A[10]), .B2(n144), .ZN(n177) );
  AOI222_X1 U201 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n153), .ZN(n176) );
  NAND2_X1 U202 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U203 ( .A1(C[14]), .A2(n149), .B1(A[14]), .B2(n143), .ZN(n185) );
  AOI222_X1 U204 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n153), .ZN(n184) );
  NAND2_X1 U205 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U206 ( .A1(C[3]), .A2(n147), .B1(A[3]), .B2(n141), .ZN(n241) );
  AOI222_X1 U207 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n155), .ZN(n240) );
  NAND2_X1 U208 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U209 ( .A1(C[7]), .A2(n145), .B1(A[7]), .B2(n139), .ZN(n297) );
  AOI222_X1 U210 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n157), .ZN(n296) );
  NAND2_X1 U211 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U212 ( .A1(C[11]), .A2(n150), .B1(A[11]), .B2(n144), .ZN(n179) );
  AOI222_X1 U213 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n153), .ZN(n178) );
  NAND2_X1 U214 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U215 ( .A1(C[15]), .A2(n149), .B1(A[15]), .B2(n143), .ZN(n187) );
  AOI222_X1 U216 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n153), .ZN(n186) );
  AOI22_X1 U217 ( .A1(C[44]), .A2(n147), .B1(A[44]), .B2(n141), .ZN(n251) );
  AOI22_X1 U218 ( .A1(C[43]), .A2(n147), .B1(A[43]), .B2(n141), .ZN(n249) );
  AOI22_X1 U219 ( .A1(C[16]), .A2(n149), .B1(A[16]), .B2(n143), .ZN(n189) );
  AOI22_X1 U220 ( .A1(C[17]), .A2(n149), .B1(A[17]), .B2(n143), .ZN(n191) );
  NAND2_X1 U221 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  NAND2_X1 U222 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI222_X1 U223 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n154), .ZN(n200) );
  AOI222_X1 U224 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n154), .ZN(n198) );
  AOI22_X1 U225 ( .A1(C[39]), .A2(n147), .B1(A[39]), .B2(n141), .ZN(n239) );
  AOI222_X1 U226 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n153), .ZN(n190) );
  AOI22_X1 U227 ( .A1(C[47]), .A2(n146), .B1(A[47]), .B2(n140), .ZN(n257) );
  AOI222_X1 U228 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n153), .ZN(n192) );
  AOI222_X1 U229 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n153), .ZN(n194) );
  CLKBUF_X1 U230 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U231 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U232 ( .A(n158), .Z(n164) );
endmodule


module G_136 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_504 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_503 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_502 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_501 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_500 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_499 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_498 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_497 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_496 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_495 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_494 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_493 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_492 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_491 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_490 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_489 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_488 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_487 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_486 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_485 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_484 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_483 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_482 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_481 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_480 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_479 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_478 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_477 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_476 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_475 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_474 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_135 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_473 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_472 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_471 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_470 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_469 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_468 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_467 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_466 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_465 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_464 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_463 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_462 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_461 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_460 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_459 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_134 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_458 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_457 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_456 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_455 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AND2_X1 U3 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
endmodule


module PG_454 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_453 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_452 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_133 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_132 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_451 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_450 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_449 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  OR2_X1 U2 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_448 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_447 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_446 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_131 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_130 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_129 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_128 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module PG_445 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_444 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_443 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_442 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_127 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_126 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_125 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module G_124 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_123 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_122 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_121 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n3;

  OR2_X2 U1 ( .A1(G_IK), .A2(n3), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n3) );
endmodule


module G_120 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module carry_generator_N64_NPB4_8 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U77 ( .A(B[59]), .B(A[59]), .Z(\PG_Network[0][0][59] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U88 ( .A(B[49]), .B(A[49]), .Z(\PG_Network[0][0][49] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U91 ( .A(B[46]), .B(A[46]), .Z(\PG_Network[0][0][46] ) );
  XOR2_X1 U92 ( .A(B[45]), .B(A[45]), .Z(\PG_Network[0][0][45] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U100 ( .A(B[38]), .B(A[38]), .Z(\PG_Network[0][0][38] ) );
  XOR2_X1 U101 ( .A(B[37]), .B(A[37]), .Z(\PG_Network[0][0][37] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U108 ( .A(B[30]), .B(A[30]), .Z(\PG_Network[0][0][30] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U110 ( .A(B[29]), .B(A[29]), .Z(\PG_Network[0][0][29] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U114 ( .A(B[25]), .B(A[25]), .Z(\PG_Network[0][0][25] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U125 ( .A(B[15]), .B(A[15]), .Z(\PG_Network[0][0][15] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_136 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n23), .Gx(\PG_Network[1][1][1] ) );
  PG_504 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_503 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_502 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_501 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_500 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_499 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_498 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_497 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_496 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_495 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_494 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_493 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_492 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_491 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_490 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_489 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_488 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_487 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_486 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_485 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_484 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_483 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_482 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_481 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_480 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_479 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_478 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_477 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_476 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_475 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_474 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_135 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_473 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_472 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_471 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_470 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_469 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_468 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_467 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_466 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_465 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_464 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_463 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_462 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_461 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_460 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_459 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_134 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_458 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_457 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_456 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_455 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_454 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_453 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(n5), .P_K_1(\PG_Network[2][0][51] ), 
        .Gx(\PG_Network[3][1][55] ), .Px(\PG_Network[3][0][55] ) );
  PG_452 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_133 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), .G_K_1(Co[1]), .Gx(Co[3]) );
  G_132 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_451 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_450 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_449 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][47] ), .Px(
        \PG_Network[4][0][47] ) );
  PG_448 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][43] ), .Px(
        \PG_Network[4][0][43] ) );
  PG_447 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][63] ), .Px(
        \PG_Network[4][0][63] ) );
  PG_446 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][59] ), .Px(
        \PG_Network[4][0][59] ) );
  G_131 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), .G_K_1(Co[3]), .Gx(Co[7]) );
  G_130 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), .G_K_1(Co[3]), .Gx(Co[6]) );
  G_129 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), .G_K_1(Co[3]), .Gx(Co[5]) );
  G_128 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), .G_K_1(Co[3]), .Gx(Co[4]) );
  PG_445 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(n7), .P_K_1(n9), .Gx(
        \PG_Network[5][1][63] ), .Px(\PG_Network[5][0][63] ) );
  PG_444 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(n7), .P_K_1(n9), .Gx(
        \PG_Network[5][1][59] ), .Px(\PG_Network[5][0][59] ) );
  PG_443 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(n22), .P_K_1(n9), .Gx(
        \PG_Network[5][1][55] ), .Px(\PG_Network[5][0][55] ) );
  PG_442 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(n22), .P_K_1(n9), .Gx(
        \PG_Network[5][1][51] ), .Px(\PG_Network[5][0][51] ) );
  G_127 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), .G_K_1(n19), .Gx(Co[15]) );
  G_126 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), .G_K_1(n19), .Gx(Co[14]) );
  G_125 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), .G_K_1(n19), .Gx(Co[13]) );
  G_124 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), .G_K_1(n19), .Gx(Co[12]) );
  G_123 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), .G_K_1(n19), .Gx(Co[11]) );
  G_122 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), .G_K_1(n19), .Gx(Co[10]) );
  G_121 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), .G_K_1(n11), .Gx(Co[9]) );
  G_120 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), .G_K_1(Co[7]), .Gx(Co[8]) );
  CLKBUF_X1 U1 ( .A(\PG_Network[2][1][51] ), .Z(n5) );
  INV_X1 U2 ( .A(A[43]), .ZN(n14) );
  INV_X1 U3 ( .A(A[55]), .ZN(n6) );
  INV_X1 U4 ( .A(A[23]), .ZN(n16) );
  INV_X1 U5 ( .A(A[19]), .ZN(n12) );
  INV_X1 U6 ( .A(A[27]), .ZN(n17) );
  INV_X1 U7 ( .A(A[35]), .ZN(n15) );
  INV_X1 U8 ( .A(A[51]), .ZN(n13) );
  INV_X1 U9 ( .A(A[39]), .ZN(n21) );
  INV_X1 U10 ( .A(A[47]), .ZN(n18) );
  INV_X1 U11 ( .A(A[31]), .ZN(n20) );
  INV_X1 U12 ( .A(A[24]), .ZN(n8) );
  INV_X1 U13 ( .A(A[44]), .ZN(n10) );
  XNOR2_X1 U14 ( .A(B[55]), .B(n6), .ZN(\PG_Network[0][0][55] ) );
  CLKBUF_X1 U15 ( .A(\PG_Network[4][1][47] ), .Z(n22) );
  CLKBUF_X1 U16 ( .A(n22), .Z(n7) );
  XNOR2_X1 U17 ( .A(B[24]), .B(n8), .ZN(\PG_Network[0][0][24] ) );
  CLKBUF_X1 U18 ( .A(\PG_Network[4][0][47] ), .Z(n9) );
  XNOR2_X1 U19 ( .A(B[44]), .B(n10), .ZN(\PG_Network[0][0][44] ) );
  CLKBUF_X1 U20 ( .A(Co[7]), .Z(n11) );
  CLKBUF_X1 U21 ( .A(n11), .Z(n19) );
  XNOR2_X1 U22 ( .A(B[19]), .B(n12), .ZN(\PG_Network[0][0][19] ) );
  XNOR2_X1 U23 ( .A(B[51]), .B(n13), .ZN(\PG_Network[0][0][51] ) );
  XNOR2_X1 U24 ( .A(B[43]), .B(n14), .ZN(\PG_Network[0][0][43] ) );
  XNOR2_X1 U25 ( .A(B[35]), .B(n15), .ZN(\PG_Network[0][0][35] ) );
  XNOR2_X1 U26 ( .A(B[23]), .B(n16), .ZN(\PG_Network[0][0][23] ) );
  XNOR2_X1 U27 ( .A(B[27]), .B(n17), .ZN(\PG_Network[0][0][27] ) );
  XNOR2_X1 U28 ( .A(B[47]), .B(n18), .ZN(\PG_Network[0][0][47] ) );
  XNOR2_X1 U29 ( .A(B[31]), .B(n20), .ZN(\PG_Network[0][0][31] ) );
  XNOR2_X1 U30 ( .A(B[39]), .B(n21), .ZN(\PG_Network[0][0][39] ) );
  AND2_X1 U31 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U32 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AND2_X1 U33 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U34 ( .A1(A[46]), .A2(B[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U35 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U36 ( .A1(A[55]), .A2(B[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U37 ( .A1(B[37]), .A2(A[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U38 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U39 ( .A1(B[45]), .A2(A[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U40 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U41 ( .A1(B[19]), .A2(A[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U42 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U43 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U44 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U45 ( .A1(B[25]), .A2(A[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U46 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U47 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U48 ( .A1(A[49]), .A2(B[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U49 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U50 ( .A1(A[59]), .A2(B[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U51 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
  AND2_X1 U52 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U53 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U54 ( .A1(B[27]), .A2(A[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U55 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U56 ( .A1(B[35]), .A2(A[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U57 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U58 ( .A1(B[51]), .A2(A[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U59 ( .A1(A[41]), .A2(B[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U60 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U61 ( .A1(B[29]), .A2(A[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U62 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U63 ( .A1(A[21]), .A2(B[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U64 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U65 ( .A1(A[53]), .A2(B[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U66 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U67 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U81 ( .A1(A[11]), .A2(B[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U85 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U90 ( .A1(A[15]), .A2(B[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U93 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U94 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U99 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U103 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U107 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U112 ( .A(n26), .ZN(n23) );
  AND2_X1 U115 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U116 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U121 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U131 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U132 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U133 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U134 ( .A1(A[7]), .A2(B[7]), .ZN(\PG_Network[0][1][7] ) );
  AND2_X1 U135 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U136 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AOI21_X1 U137 ( .B1(A[0]), .B2(B[0]), .A(n24), .ZN(n26) );
  INV_X1 U138 ( .A(n25), .ZN(n24) );
  OAI21_X1 U139 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n25) );
  AND2_X1 U140 ( .A1(B[23]), .A2(A[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U141 ( .A1(B[44]), .A2(A[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U142 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U143 ( .A1(A[43]), .A2(B[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U144 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U145 ( .A1(B[31]), .A2(A[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U146 ( .A1(B[47]), .A2(A[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U147 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U148 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
endmodule


module FA_1024 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1023 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1022 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1021 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_256 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1024 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1023 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1022 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1021 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1020 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1019 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1018 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1017 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_255 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1020 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1019 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1018 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1017 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_128 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U2 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_128 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_256 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_255 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_128 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1016 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1015 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1014 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1013 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_254 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1016 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1015 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1014 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1013 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1012 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1011 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1010 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1009 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_253 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1012 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1011 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1010 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1009 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_127 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_127 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_254 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_253 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_127 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1008 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1007 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1006 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1005 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_252 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1008 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1007 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1006 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1005 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_1004 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1003 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1002 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1001 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_251 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1004 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1003 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1002 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1001 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_126 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_126 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_252 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_251 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_126 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_1000 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_999 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_998 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_997 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_250 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1000 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_999 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_998 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_997 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_996 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_995 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_994 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_993 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_249 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_996 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_995 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_994 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_993 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_125 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_125 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_250 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_249 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_125 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_992 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_991 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_990 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_989 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_248 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_992 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_991 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_990 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_989 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_988 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_987 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_986 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_985 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_247 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_988 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_987 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_986 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_985 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_124 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_124 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_248 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_247 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_124 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_984 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_983 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_982 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_981 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_246 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_984 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_983 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_982 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_981 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_980 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_979 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_978 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_977 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_245 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_980 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_979 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_978 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_977 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_123 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U6 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U7 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U8 ( .A(sel), .ZN(n13) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
endmodule


module carry_select_block_NPB4_123 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_246 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_245 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_123 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_976 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_975 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_974 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_973 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  OR2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_244 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_976 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_975 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_974 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_973 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_972 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_971 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_970 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_969 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_243 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_972 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_971 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_970 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_969 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_122 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  CLKBUF_X1 U1 ( .A(sel), .Z(n10) );
  INV_X2 U2 ( .A(n16), .ZN(Y[0]) );
  BUF_X1 U3 ( .A(n15), .Z(n5) );
  INV_X1 U4 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U5 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n10), .B1(B[1]), .B2(n5), .ZN(n17) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U9 ( .A(sel), .ZN(n15) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n15), .ZN(n19) );
  INV_X2 U11 ( .A(n18), .ZN(Y[2]) );
endmodule


module carry_select_block_NPB4_122 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_244 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_243 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_122 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_968 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(n4), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_967 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_966 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_965 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  OR2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_242 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_968 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_967 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_966 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_965 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_964 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_963 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_962 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_961 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_241 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_964 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_963 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_962 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_961 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_121 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U4 ( .A(sel), .ZN(n10) );
  INV_X1 U5 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[0]), .B1(n10), .B2(B[0]), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(n15), .B2(B[1]), .ZN(n17) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n15), .ZN(n19) );
endmodule


module carry_select_block_NPB4_121 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_242 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_241 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_121 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_960 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_959 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_958 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_957 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n8, n10, n11;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n10) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n4), .A2(n10), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n10), .ZN(n5) );
  CLKBUF_X1 U7 ( .A(Ci), .Z(n8) );
  INV_X1 U8 ( .A(n11), .ZN(Co) );
  AOI22_X1 U9 ( .A1(B), .A2(A), .B1(n10), .B2(n8), .ZN(n11) );
endmodule


module RCA_N4_240 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_960 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_959 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_958 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_957 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_956 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_955 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_954 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_953 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_239 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_956 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_955 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_954 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_953 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_120 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(n15), .Z(n5) );
  INV_X1 U2 ( .A(n16), .ZN(Y[0]) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n10) );
  INV_X1 U4 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(n10), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_120 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_240 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_239 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_120 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_952 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n8), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_951 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_950 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_949 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n8, n10, n11;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n5), .ZN(n4) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n5), .A2(n10), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n7), .A2(n8), .ZN(S) );
  INV_X1 U6 ( .A(Ci), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(n6) );
  INV_X1 U8 ( .A(n11), .ZN(Co) );
  AOI22_X1 U9 ( .A1(B), .A2(A), .B1(n10), .B2(n4), .ZN(n11) );
endmodule


module RCA_N4_238 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_952 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_951 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_950 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_949 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_948 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_947 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_946 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_945 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_237 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_948 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_947 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_946 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_945 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_119 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n17), .ZN(Y[1]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n10) );
  BUF_X1 U3 ( .A(n15), .Z(n5) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(n10), .A2(A[2]), .B1(n5), .B2(B[2]), .ZN(n18) );
  AOI22_X1 U8 ( .A1(n10), .A2(A[1]), .B1(n5), .B2(B[1]), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n10), .B1(n5), .B2(B[3]), .ZN(n19) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_119 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_238 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_237 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_119 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_944 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n6) );
  XNOR2_X1 U4 ( .A(n6), .B(n4), .ZN(n5) );
  XNOR2_X1 U5 ( .A(n6), .B(B), .ZN(n8) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_943 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_942 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_941 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_236 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_944 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_943 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_942 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_941 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_940 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_939 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_938 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_937 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_235 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_940 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_939 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_938 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_937 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_118 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  CLKBUF_X1 U1 ( .A(sel), .Z(n10) );
  INV_X1 U2 ( .A(sel), .ZN(n5) );
  INV_X1 U3 ( .A(sel), .ZN(n15) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(n10), .B1(n15), .B2(B[2]), .ZN(n18) );
  INV_X1 U6 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U7 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(n10), .B1(n15), .B2(B[3]), .ZN(n19) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n15), .ZN(n17) );
  INV_X1 U10 ( .A(n16), .ZN(Y[0]) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n5), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_118 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_236 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_235 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_118 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_936 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_935 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_934 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_933 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_234 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_936 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_935 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_934 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_933 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_932 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_931 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_930 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_929 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_233 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_932 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_931 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_930 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_929 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_117 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  CLKBUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X2 U2 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U3 ( .A(sel), .ZN(n10) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U6 ( .A1(n5), .A2(A[2]), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[1]), .B1(n10), .B2(B[1]), .ZN(n17) );
  INV_X1 U8 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n10), .ZN(n19) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_117 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_234 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_233 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_117 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_928 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n9), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(n5), .B(B), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n8), .A2(n7), .ZN(Co) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(n7) );
  NAND2_X1 U7 ( .A1(n9), .A2(Ci), .ZN(n8) );
endmodule


module FA_927 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_926 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_925 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_232 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_928 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_927 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_926 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_925 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_924 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_923 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_922 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_921 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_231 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_924 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_923 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_922 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_921 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_116 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U2 ( .A(sel), .ZN(n5) );
  INV_X1 U3 ( .A(n11), .ZN(n10) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[1]) );
  CLKBUF_X1 U6 ( .A(sel), .Z(n11) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(n11), .B1(B[3]), .B2(n10), .ZN(n19) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n11), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n5), .ZN(n17) );
  INV_X1 U10 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n5), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_116 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_232 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_231 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_116 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_920 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_919 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_918 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_917 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_230 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_920 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_919 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_918 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_917 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_916 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_915 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_914 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_913 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_229 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_916 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_915 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_914 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_913 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_115 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18;

  CLKBUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(sel), .ZN(n10) );
  INV_X1 U3 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U6 ( .A(n15), .ZN(Y[0]) );
  AOI22_X1 U7 ( .A1(n5), .A2(A[3]), .B1(B[3]), .B2(n10), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n10), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n10), .ZN(n16) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n10), .ZN(n15) );
endmodule


module carry_select_block_NPB4_115 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_230 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_229 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_115 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_912 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_911 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_910 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_909 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_228 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_912 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_911 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_910 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_909 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_908 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_907 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_906 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_905 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_227 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_908 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_907 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_906 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_905 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_114 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X2 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(sel), .ZN(n13) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_114 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_228 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_227 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_114 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_904 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_903 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_902 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_901 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_226 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_904 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_903 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_902 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_901 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_900 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_899 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_898 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_897 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_225 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_900 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_899 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_898 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_897 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_113 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_113 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_226 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_225 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_113 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_8 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_128 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_127 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_126 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_125 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_124 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_123 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_122 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_121 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_120 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_119 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_118 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), .S(S[43:40]) );
  carry_select_block_NPB4_117 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), .S(S[47:44]) );
  carry_select_block_NPB4_116 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), .S(S[51:48]) );
  carry_select_block_NPB4_115 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), .S(S[55:52]) );
  carry_select_block_NPB4_114 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), .S(S[59:56]) );
  carry_select_block_NPB4_113 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), .S(S[63:60]) );
endmodule


module P4_ADDER_N64_8 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_8 CGEN ( .A(A), .B({B[63:45], n21, B[43:41], n12, 
        B[39:37], n18, B[35:33], n10, B[31:29], n5, B[27:21], n22, B[19:0]}), 
        .Cin(Cin), .Co(CoutCgen) );
  sum_generator_N64_NPB4_8 SGEN ( .A(A), .B({B[63:48], n17, n9, n11, B[44], 
        n20, B[42:40], n6, n3, B[37:36], n15, B[34:32], n13, B[30:28], n1, 
        B[26:24], n4, B[22:20], n7, B[18:0]}), .Ci({CoutCgen, Cin}), .S(S), 
        .Co(Cout) );
  BUF_X1 U1 ( .A(B[45]), .Z(n11) );
  BUF_X1 U2 ( .A(B[27]), .Z(n1) );
  INV_X1 U3 ( .A(B[38]), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  CLKBUF_X1 U5 ( .A(B[44]), .Z(n21) );
  CLKBUF_X1 U6 ( .A(B[28]), .Z(n5) );
  CLKBUF_X1 U7 ( .A(B[23]), .Z(n4) );
  CLKBUF_X1 U8 ( .A(B[39]), .Z(n6) );
  CLKBUF_X1 U9 ( .A(B[20]), .Z(n22) );
  CLKBUF_X1 U10 ( .A(B[19]), .Z(n7) );
  INV_X1 U11 ( .A(B[46]), .ZN(n8) );
  INV_X1 U12 ( .A(n8), .ZN(n9) );
  CLKBUF_X1 U13 ( .A(B[32]), .Z(n10) );
  CLKBUF_X1 U14 ( .A(B[40]), .Z(n12) );
  CLKBUF_X1 U15 ( .A(B[31]), .Z(n13) );
  INV_X1 U16 ( .A(B[35]), .ZN(n14) );
  INV_X1 U17 ( .A(n14), .ZN(n15) );
  INV_X1 U18 ( .A(B[47]), .ZN(n16) );
  INV_X1 U19 ( .A(n16), .ZN(n17) );
  CLKBUF_X1 U20 ( .A(B[36]), .Z(n18) );
  INV_X1 U21 ( .A(B[43]), .ZN(n19) );
  INV_X1 U22 ( .A(n19), .ZN(n20) );
endmodule


module Booth_Encoder_7 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_7 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306;

  NAND2_X2 U1 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  NAND2_X1 U2 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  NAND2_X1 U3 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  NAND2_X1 U4 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  NAND2_X1 U5 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  NAND2_X1 U6 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  NOR3_X1 U7 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U8 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  BUF_X1 U9 ( .A(n158), .Z(n162) );
  BUF_X1 U10 ( .A(n158), .Z(n161) );
  BUF_X1 U11 ( .A(n158), .Z(n159) );
  BUF_X1 U12 ( .A(n158), .Z(n160) );
  BUF_X1 U13 ( .A(n158), .Z(n163) );
  BUF_X1 U14 ( .A(n151), .Z(n155) );
  BUF_X1 U15 ( .A(n165), .Z(n169) );
  BUF_X1 U16 ( .A(n151), .Z(n153) );
  BUF_X1 U17 ( .A(n165), .Z(n167) );
  BUF_X1 U18 ( .A(n151), .Z(n154) );
  BUF_X1 U19 ( .A(n165), .Z(n168) );
  BUF_X1 U20 ( .A(n303), .Z(n158) );
  NOR4_X1 U21 ( .A1(n150), .A2(n144), .A3(n153), .A4(n167), .ZN(n303) );
  BUF_X1 U22 ( .A(n152), .Z(n156) );
  BUF_X1 U23 ( .A(n166), .Z(n170) );
  BUF_X1 U24 ( .A(n152), .Z(n157) );
  BUF_X1 U25 ( .A(n166), .Z(n171) );
  BUF_X1 U26 ( .A(n301), .Z(n148) );
  BUF_X1 U27 ( .A(n301), .Z(n147) );
  BUF_X1 U28 ( .A(n301), .Z(n149) );
  BUF_X1 U29 ( .A(n304), .Z(n165) );
  BUF_X1 U30 ( .A(n302), .Z(n151) );
  BUF_X1 U31 ( .A(n301), .Z(n146) );
  BUF_X1 U32 ( .A(n304), .Z(n166) );
  BUF_X1 U33 ( .A(n302), .Z(n152) );
  BUF_X1 U34 ( .A(n301), .Z(n145) );
  BUF_X1 U35 ( .A(n300), .Z(n142) );
  BUF_X1 U36 ( .A(n300), .Z(n139) );
  BUF_X1 U37 ( .A(n300), .Z(n141) );
  BUF_X1 U38 ( .A(n300), .Z(n140) );
  BUF_X1 U39 ( .A(n300), .Z(n143) );
  INV_X1 U40 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U41 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n304) );
  AND3_X1 U42 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U43 ( .A(sel[2]), .ZN(n173) );
  NAND2_X1 U44 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI22_X1 U45 ( .A1(C[22]), .A2(n149), .B1(A[22]), .B2(n143), .ZN(n203) );
  AOI22_X1 U46 ( .A1(C[24]), .A2(n149), .B1(A[24]), .B2(n143), .ZN(n207) );
  AOI222_X1 U47 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n154), .ZN(n206) );
  AOI22_X1 U48 ( .A1(C[28]), .A2(n148), .B1(A[28]), .B2(n142), .ZN(n215) );
  AOI222_X1 U49 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n154), .ZN(n214) );
  NAND2_X1 U50 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI22_X1 U51 ( .A1(C[25]), .A2(n148), .B1(A[25]), .B2(n142), .ZN(n209) );
  AOI222_X1 U52 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n154), .ZN(n208) );
  AOI222_X1 U53 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n153), .ZN(n192) );
  NAND2_X1 U54 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  AOI22_X1 U55 ( .A1(C[20]), .A2(n149), .B1(A[20]), .B2(n143), .ZN(n199) );
  NAND2_X1 U56 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI222_X1 U57 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n155), .ZN(n244) );
  NAND2_X1 U58 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI22_X1 U59 ( .A1(C[42]), .A2(n147), .B1(A[42]), .B2(n141), .ZN(n247) );
  AOI222_X1 U60 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n155), .ZN(n246) );
  NAND2_X1 U61 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI22_X1 U62 ( .A1(C[21]), .A2(n149), .B1(A[21]), .B2(n143), .ZN(n201) );
  NAND2_X1 U63 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI22_X1 U64 ( .A1(C[23]), .A2(n149), .B1(A[23]), .B2(n143), .ZN(n205) );
  NAND2_X1 U65 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI22_X1 U66 ( .A1(C[26]), .A2(n148), .B1(A[26]), .B2(n142), .ZN(n211) );
  AOI222_X1 U67 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n154), .ZN(n210) );
  NAND2_X1 U68 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI22_X1 U69 ( .A1(C[34]), .A2(n148), .B1(A[34]), .B2(n142), .ZN(n229) );
  AOI222_X1 U70 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n155), .ZN(n228) );
  NAND2_X1 U71 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  AOI22_X1 U72 ( .A1(C[56]), .A2(n146), .B1(A[56]), .B2(n140), .ZN(n277) );
  AOI222_X1 U73 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n157), .ZN(n276) );
  NAND2_X1 U74 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  AOI22_X1 U75 ( .A1(C[53]), .A2(n146), .B1(A[53]), .B2(n140), .ZN(n271) );
  AOI222_X1 U76 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n156), .ZN(n270) );
  NAND2_X1 U77 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  AOI22_X1 U78 ( .A1(C[57]), .A2(n145), .B1(A[57]), .B2(n139), .ZN(n279) );
  AOI222_X1 U79 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n157), .ZN(n278) );
  NAND2_X1 U80 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI22_X1 U81 ( .A1(C[55]), .A2(n146), .B1(A[55]), .B2(n140), .ZN(n275) );
  AOI222_X1 U82 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n156), .ZN(n274) );
  NAND2_X1 U83 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI22_X1 U84 ( .A1(C[33]), .A2(n148), .B1(A[33]), .B2(n142), .ZN(n227) );
  AOI222_X1 U85 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n155), .ZN(n226) );
  NAND2_X1 U86 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI22_X1 U87 ( .A1(C[27]), .A2(n148), .B1(A[27]), .B2(n142), .ZN(n213) );
  AOI222_X1 U88 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n154), .ZN(n212) );
  NAND2_X1 U89 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI222_X1 U90 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n154), .ZN(n222) );
  AOI22_X1 U91 ( .A1(C[31]), .A2(n148), .B1(A[31]), .B2(n142), .ZN(n223) );
  NAND2_X1 U92 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI222_X1 U93 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n155), .ZN(n230) );
  AOI22_X1 U94 ( .A1(C[35]), .A2(n148), .B1(A[35]), .B2(n142), .ZN(n231) );
  AOI22_X1 U95 ( .A1(C[32]), .A2(n148), .B1(A[32]), .B2(n142), .ZN(n225) );
  AOI222_X1 U96 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n155), .ZN(n224) );
  NAND2_X1 U97 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI22_X1 U98 ( .A1(C[37]), .A2(n147), .B1(A[37]), .B2(n141), .ZN(n235) );
  AOI222_X1 U99 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n155), .ZN(n234) );
  NAND2_X1 U100 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U101 ( .A1(C[30]), .A2(n148), .B1(A[30]), .B2(n142), .ZN(n221) );
  AOI222_X1 U102 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n154), .ZN(n220) );
  NAND2_X1 U103 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI22_X1 U104 ( .A1(C[38]), .A2(n147), .B1(A[38]), .B2(n141), .ZN(n237) );
  AOI222_X1 U105 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n155), .ZN(n236) );
  NAND2_X1 U106 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI222_X1 U107 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n156), .ZN(n264) );
  AOI22_X1 U108 ( .A1(C[50]), .A2(n146), .B1(A[50]), .B2(n140), .ZN(n265) );
  NAND2_X1 U109 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI22_X1 U110 ( .A1(C[54]), .A2(n146), .B1(A[54]), .B2(n140), .ZN(n273) );
  AOI222_X1 U111 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n156), .ZN(n272) );
  NAND2_X1 U112 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI222_X1 U113 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n156), .ZN(n254) );
  NAND2_X1 U114 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI22_X1 U115 ( .A1(C[29]), .A2(n148), .B1(A[29]), .B2(n142), .ZN(n217) );
  AOI222_X1 U116 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n154), .ZN(n216) );
  AOI22_X1 U117 ( .A1(C[36]), .A2(n147), .B1(A[36]), .B2(n141), .ZN(n233) );
  AOI222_X1 U118 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n155), .ZN(n232) );
  AOI22_X1 U119 ( .A1(C[40]), .A2(n147), .B1(A[40]), .B2(n141), .ZN(n243) );
  AOI222_X1 U120 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n155), .ZN(n242) );
  NAND2_X1 U121 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI222_X1 U122 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n156), .ZN(n260) );
  NAND2_X1 U123 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI222_X1 U124 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n156), .ZN(n252) );
  NAND2_X1 U125 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  AOI22_X1 U126 ( .A1(C[52]), .A2(n146), .B1(A[52]), .B2(n140), .ZN(n269) );
  AOI222_X1 U127 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n156), .ZN(n268) );
  NAND2_X1 U128 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  AOI22_X1 U129 ( .A1(C[51]), .A2(n146), .B1(A[51]), .B2(n140), .ZN(n267) );
  AOI222_X1 U130 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n156), .ZN(n266) );
  NAND2_X1 U131 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI222_X1 U132 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n155), .ZN(n238) );
  AOI22_X1 U133 ( .A1(C[39]), .A2(n147), .B1(A[39]), .B2(n141), .ZN(n239) );
  NAND2_X1 U134 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI222_X1 U135 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n155), .ZN(n248) );
  AOI22_X1 U136 ( .A1(C[43]), .A2(n147), .B1(A[43]), .B2(n141), .ZN(n249) );
  NAND2_X1 U137 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI222_X1 U138 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n156), .ZN(n256) );
  AOI22_X1 U139 ( .A1(C[47]), .A2(n146), .B1(A[47]), .B2(n140), .ZN(n257) );
  NAND2_X1 U140 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  AOI22_X1 U141 ( .A1(C[44]), .A2(n147), .B1(A[44]), .B2(n141), .ZN(n251) );
  AOI222_X1 U142 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n156), .ZN(n250) );
  AOI22_X1 U143 ( .A1(C[48]), .A2(n146), .B1(A[48]), .B2(n140), .ZN(n259) );
  AOI222_X1 U144 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n156), .ZN(n258) );
  NAND2_X1 U145 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U146 ( .A1(C[60]), .A2(n145), .B1(A[60]), .B2(n139), .ZN(n287) );
  AOI222_X1 U147 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n157), .ZN(n286) );
  NAND2_X1 U148 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U149 ( .A1(C[61]), .A2(n145), .B1(A[61]), .B2(n139), .ZN(n289) );
  AOI222_X1 U150 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n157), .ZN(n288) );
  NAND2_X1 U151 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI22_X1 U152 ( .A1(C[58]), .A2(n145), .B1(A[58]), .B2(n139), .ZN(n281) );
  AOI222_X1 U153 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n157), .ZN(n280) );
  NAND2_X1 U154 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U155 ( .A1(C[62]), .A2(n145), .B1(A[62]), .B2(n139), .ZN(n291) );
  AOI222_X1 U156 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n157), .ZN(n290) );
  NAND2_X1 U157 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U158 ( .A1(C[59]), .A2(n145), .B1(A[59]), .B2(n139), .ZN(n283) );
  AOI222_X1 U159 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n157), .ZN(n282) );
  NAND2_X1 U160 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U161 ( .A1(C[63]), .A2(n145), .B1(A[63]), .B2(n139), .ZN(n293) );
  AOI222_X1 U162 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n157), .ZN(n292) );
  NAND2_X1 U163 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U164 ( .A1(C[0]), .A2(n145), .B1(A[0]), .B2(n139), .ZN(n175) );
  AOI222_X1 U165 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n153), .ZN(n174) );
  NAND2_X1 U166 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U167 ( .A1(C[4]), .A2(n146), .B1(A[4]), .B2(n140), .ZN(n263) );
  AOI222_X1 U168 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n156), .ZN(n262) );
  NAND2_X1 U169 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI22_X1 U170 ( .A1(C[8]), .A2(n145), .B1(A[8]), .B2(n139), .ZN(n299) );
  AOI222_X1 U171 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n157), .ZN(n298) );
  NAND2_X1 U172 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  AOI22_X1 U173 ( .A1(C[12]), .A2(n150), .B1(A[12]), .B2(n144), .ZN(n181) );
  AOI222_X1 U174 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n153), .ZN(n180) );
  NAND2_X1 U175 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  AOI22_X1 U176 ( .A1(C[16]), .A2(n149), .B1(A[16]), .B2(n143), .ZN(n189) );
  AOI222_X1 U177 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n153), .ZN(n188) );
  NAND2_X1 U178 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U179 ( .A1(C[1]), .A2(n149), .B1(A[1]), .B2(n143), .ZN(n197) );
  AOI222_X1 U180 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n153), .ZN(n196) );
  NAND2_X1 U181 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U182 ( .A1(C[5]), .A2(n145), .B1(A[5]), .B2(n139), .ZN(n285) );
  AOI222_X1 U183 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n157), .ZN(n284) );
  NAND2_X1 U184 ( .A1(n306), .A2(n305), .ZN(Y[9]) );
  AOI22_X1 U185 ( .A1(C[9]), .A2(n147), .B1(A[9]), .B2(n141), .ZN(n306) );
  AOI222_X1 U186 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n157), .ZN(n305) );
  NAND2_X1 U187 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U188 ( .A1(C[13]), .A2(n150), .B1(A[13]), .B2(n144), .ZN(n183) );
  AOI222_X1 U189 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n153), .ZN(n182) );
  NAND2_X1 U190 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI22_X1 U191 ( .A1(C[17]), .A2(n149), .B1(A[17]), .B2(n143), .ZN(n191) );
  AOI222_X1 U192 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n153), .ZN(n190) );
  NAND2_X1 U193 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U194 ( .A1(C[2]), .A2(n148), .B1(A[2]), .B2(n142), .ZN(n219) );
  AOI222_X1 U195 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n154), .ZN(n218) );
  NAND2_X1 U196 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U197 ( .A1(C[6]), .A2(n145), .B1(A[6]), .B2(n139), .ZN(n295) );
  AOI222_X1 U198 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n157), .ZN(n294) );
  NAND2_X1 U199 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U200 ( .A1(C[10]), .A2(n150), .B1(A[10]), .B2(n144), .ZN(n177) );
  AOI222_X1 U201 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n153), .ZN(n176) );
  NAND2_X1 U202 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U203 ( .A1(C[14]), .A2(n149), .B1(A[14]), .B2(n143), .ZN(n185) );
  AOI222_X1 U204 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n153), .ZN(n184) );
  NAND2_X1 U205 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U206 ( .A1(C[3]), .A2(n147), .B1(A[3]), .B2(n141), .ZN(n241) );
  AOI222_X1 U207 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n155), .ZN(n240) );
  NAND2_X1 U208 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U209 ( .A1(C[7]), .A2(n145), .B1(A[7]), .B2(n139), .ZN(n297) );
  AOI222_X1 U210 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n157), .ZN(n296) );
  NAND2_X1 U211 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U212 ( .A1(C[11]), .A2(n150), .B1(A[11]), .B2(n144), .ZN(n179) );
  AOI222_X1 U213 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n153), .ZN(n178) );
  NAND2_X1 U214 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U215 ( .A1(C[15]), .A2(n149), .B1(A[15]), .B2(n143), .ZN(n187) );
  AOI222_X1 U216 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n153), .ZN(n186) );
  AOI22_X1 U217 ( .A1(C[46]), .A2(n146), .B1(A[46]), .B2(n140), .ZN(n255) );
  AOI22_X1 U218 ( .A1(C[45]), .A2(n147), .B1(A[45]), .B2(n141), .ZN(n253) );
  AOI22_X1 U219 ( .A1(C[18]), .A2(n149), .B1(A[18]), .B2(n143), .ZN(n193) );
  AOI22_X1 U220 ( .A1(C[19]), .A2(n149), .B1(A[19]), .B2(n143), .ZN(n195) );
  NAND2_X1 U221 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  NAND2_X1 U222 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI222_X1 U223 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n154), .ZN(n204) );
  AOI222_X1 U224 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n154), .ZN(n202) );
  AOI22_X1 U225 ( .A1(C[41]), .A2(n147), .B1(A[41]), .B2(n141), .ZN(n245) );
  AOI222_X1 U226 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n153), .ZN(n194) );
  AOI22_X1 U227 ( .A1(C[49]), .A2(n146), .B1(A[49]), .B2(n140), .ZN(n261) );
  AOI222_X1 U228 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n154), .ZN(n200) );
  AOI222_X1 U229 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n154), .ZN(n198) );
  CLKBUF_X1 U230 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U231 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U232 ( .A(n158), .Z(n164) );
endmodule


module G_119 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_441 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_440 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_439 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_438 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_437 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_436 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_435 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_434 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_433 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_432 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_431 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_430 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_429 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_428 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_427 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_426 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_425 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_424 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_423 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_422 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_421 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_420 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_419 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_418 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_417 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_416 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_415 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_414 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_413 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_412 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_411 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_118 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_410 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_409 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_408 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_407 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_406 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_405 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_404 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AND2_X1 U3 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
endmodule


module PG_403 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_402 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_401 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  OR2_X1 U2 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_400 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_399 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_398 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_397 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_396 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_117 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_395 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_394 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_393 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_392 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AND2_X1 U3 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
endmodule


module PG_391 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_390 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_389 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_116 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_115 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_388 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_387 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_386 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_385 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_384 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_383 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_114 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_113 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_112 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_111 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_382 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_381 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_380 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_379 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_110 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_109 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_108 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_107 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_106 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_105 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_104 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_103 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module carry_generator_N64_NPB4_7 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U77 ( .A(B[59]), .B(A[59]), .Z(\PG_Network[0][0][59] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U88 ( .A(B[49]), .B(A[49]), .Z(\PG_Network[0][0][49] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U92 ( .A(B[45]), .B(A[45]), .Z(\PG_Network[0][0][45] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U100 ( .A(B[38]), .B(A[38]), .Z(\PG_Network[0][0][38] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U108 ( .A(B[30]), .B(A[30]), .Z(\PG_Network[0][0][30] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U110 ( .A(B[29]), .B(A[29]), .Z(\PG_Network[0][0][29] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U121 ( .A(B[19]), .B(A[19]), .Z(\PG_Network[0][0][19] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U125 ( .A(B[15]), .B(A[15]), .Z(\PG_Network[0][0][15] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_119 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n21), .Gx(\PG_Network[1][1][1] ) );
  PG_441 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_440 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_439 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_438 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_437 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_436 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_435 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_434 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_433 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_432 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_431 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_430 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_429 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_428 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_427 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_426 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_425 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_424 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_423 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_422 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_421 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_420 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_419 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_418 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_417 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_416 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_415 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_414 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_413 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_412 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_411 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_118 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_410 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_409 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_408 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_407 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_406 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_405 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_404 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_403 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_402 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_401 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_400 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_399 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_398 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_397 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_396 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_117 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_395 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_394 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_393 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_392 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_391 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(n17), .P_K_1(\PG_Network[2][0][43] ), 
        .Gx(\PG_Network[3][1][47] ), .Px(\PG_Network[3][0][47] ) );
  PG_390 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_389 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_116 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), .G_K_1(Co[1]), .Gx(Co[3]) );
  G_115 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_388 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_387 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_386 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][47] ), .Px(
        \PG_Network[4][0][47] ) );
  PG_385 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][43] ), .Px(
        \PG_Network[4][0][43] ) );
  PG_384 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][63] ), .Px(
        \PG_Network[4][0][63] ) );
  PG_383 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][59] ), .Px(
        \PG_Network[4][0][59] ) );
  G_114 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), .G_K_1(Co[3]), .Gx(Co[7]) );
  G_113 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), .G_K_1(Co[3]), .Gx(Co[6]) );
  G_112 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), .G_K_1(Co[3]), .Gx(Co[5]) );
  G_111 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), .G_K_1(Co[3]), .Gx(Co[4]) );
  PG_382 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(n20), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][63] ), .Px(\PG_Network[5][0][63] ) );
  PG_381 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(n20), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][59] ), .Px(\PG_Network[5][0][59] ) );
  PG_380 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(n20), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][55] ), .Px(\PG_Network[5][0][55] ) );
  PG_379 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][51] ), .Px(
        \PG_Network[5][0][51] ) );
  G_110 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), .G_K_1(n12), .Gx(Co[15]) );
  G_109 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), .G_K_1(n12), .Gx(Co[14]) );
  G_108 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), .G_K_1(n12), .Gx(Co[13]) );
  G_107 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), .G_K_1(n12), .Gx(Co[12]) );
  G_106 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), .G_K_1(Co[7]), .Gx(Co[11]) );
  G_105 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), .G_K_1(Co[7]), .Gx(Co[10]) );
  G_104 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), .G_K_1(Co[7]), .Gx(Co[9]) );
  G_103 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), .G_K_1(Co[7]), .Gx(Co[8]) );
  INV_X1 U1 ( .A(A[23]), .ZN(n10) );
  INV_X1 U2 ( .A(A[55]), .ZN(n6) );
  INV_X1 U3 ( .A(A[46]), .ZN(n9) );
  INV_X1 U4 ( .A(A[43]), .ZN(n8) );
  INV_X1 U5 ( .A(A[25]), .ZN(n5) );
  INV_X1 U6 ( .A(A[27]), .ZN(n13) );
  INV_X1 U7 ( .A(A[31]), .ZN(n16) );
  INV_X1 U8 ( .A(A[35]), .ZN(n11) );
  INV_X1 U9 ( .A(A[51]), .ZN(n19) );
  INV_X1 U10 ( .A(A[39]), .ZN(n15) );
  INV_X1 U11 ( .A(A[47]), .ZN(n18) );
  INV_X1 U12 ( .A(A[37]), .ZN(n14) );
  INV_X1 U13 ( .A(A[40]), .ZN(n7) );
  XNOR2_X1 U14 ( .A(B[25]), .B(n5), .ZN(\PG_Network[0][0][25] ) );
  XNOR2_X1 U15 ( .A(B[55]), .B(n6), .ZN(\PG_Network[0][0][55] ) );
  XNOR2_X1 U16 ( .A(B[40]), .B(n7), .ZN(\PG_Network[0][0][40] ) );
  XNOR2_X1 U17 ( .A(B[43]), .B(n8), .ZN(\PG_Network[0][0][43] ) );
  XNOR2_X1 U18 ( .A(B[46]), .B(n9), .ZN(\PG_Network[0][0][46] ) );
  XNOR2_X1 U19 ( .A(B[23]), .B(n10), .ZN(\PG_Network[0][0][23] ) );
  CLKBUF_X1 U20 ( .A(\PG_Network[4][1][47] ), .Z(n20) );
  XNOR2_X1 U21 ( .A(B[35]), .B(n11), .ZN(\PG_Network[0][0][35] ) );
  CLKBUF_X1 U22 ( .A(Co[7]), .Z(n12) );
  XNOR2_X1 U23 ( .A(B[27]), .B(n13), .ZN(\PG_Network[0][0][27] ) );
  XNOR2_X1 U24 ( .A(B[37]), .B(n14), .ZN(\PG_Network[0][0][37] ) );
  XNOR2_X1 U25 ( .A(B[39]), .B(n15), .ZN(\PG_Network[0][0][39] ) );
  XNOR2_X1 U26 ( .A(B[31]), .B(n16), .ZN(\PG_Network[0][0][31] ) );
  CLKBUF_X1 U27 ( .A(\PG_Network[2][1][43] ), .Z(n17) );
  XNOR2_X1 U28 ( .A(B[47]), .B(n18), .ZN(\PG_Network[0][0][47] ) );
  XNOR2_X1 U29 ( .A(B[51]), .B(n19), .ZN(\PG_Network[0][0][51] ) );
  AND2_X1 U30 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U31 ( .A1(B[27]), .A2(A[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U32 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U33 ( .A1(B[31]), .A2(A[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U34 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U35 ( .A1(A[46]), .A2(B[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U36 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U37 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U38 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AND2_X1 U39 ( .A1(A[23]), .A2(B[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U40 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U41 ( .A1(A[55]), .A2(B[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U42 ( .A1(B[41]), .A2(A[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U43 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U44 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U45 ( .A1(A[19]), .A2(B[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U46 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U47 ( .A1(B[35]), .A2(A[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U48 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U49 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U50 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U51 ( .A1(A[59]), .A2(B[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U52 ( .A1(A[49]), .A2(B[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U53 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
  AND2_X1 U54 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U55 ( .A1(A[21]), .A2(B[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U56 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U57 ( .A1(B[37]), .A2(A[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U58 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U59 ( .A1(A[53]), .A2(B[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U60 ( .A1(B[29]), .A2(A[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U61 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U62 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U63 ( .A1(A[11]), .A2(B[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U64 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U65 ( .A1(A[15]), .A2(B[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U66 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U67 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U81 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U85 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U90 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U91 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U94 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U97 ( .A(n24), .ZN(n21) );
  AND2_X1 U99 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U101 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U103 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U107 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U112 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U114 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U116 ( .A1(A[7]), .A2(B[7]), .ZN(\PG_Network[0][1][7] ) );
  AND2_X1 U131 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U132 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AOI21_X1 U133 ( .B1(A[0]), .B2(B[0]), .A(n22), .ZN(n24) );
  INV_X1 U134 ( .A(n23), .ZN(n22) );
  OAI21_X1 U135 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n23) );
  AND2_X1 U136 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U137 ( .A1(A[43]), .A2(B[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U138 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U139 ( .A1(B[25]), .A2(A[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U140 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U141 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U142 ( .A1(B[47]), .A2(A[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U143 ( .A1(A[45]), .A2(B[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U144 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U145 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U146 ( .A1(B[51]), .A2(A[51]), .ZN(\PG_Network[0][1][51] ) );
endmodule


module FA_896 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_895 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_894 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_893 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_224 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_896 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_895 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_894 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_893 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_892 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_891 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_890 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_889 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_223 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_892 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_891 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_890 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_889 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_112 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U2 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_112 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_224 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_223 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_112 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_888 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_887 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_886 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_885 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_222 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_888 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_887 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_886 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_885 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_884 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_883 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_882 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_881 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_221 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_884 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_883 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_882 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_881 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_111 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_111 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_222 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_221 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_111 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_880 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_879 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_878 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_877 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_220 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_880 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_879 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_878 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_877 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_876 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_875 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_874 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_873 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_219 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_876 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_875 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_874 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_873 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_110 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_110 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_220 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_219 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_110 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_872 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_871 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_870 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_869 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_218 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_872 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_871 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_870 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_869 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_868 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_867 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_866 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_865 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_217 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_868 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_867 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_866 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_865 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_109 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_109 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_218 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_217 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_109 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_864 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_863 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_862 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_861 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_216 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_864 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_863 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_862 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_861 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_860 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_859 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_858 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_857 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_215 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_860 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_859 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_858 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_857 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_108 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_108 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_216 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_215 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_108 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_856 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_855 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_854 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_853 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_214 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_856 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_855 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_854 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_853 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_852 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_851 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_850 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_849 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_213 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_852 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_851 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_850 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_849 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_107 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(sel), .ZN(n13) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n13), .ZN(n17) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_107 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_214 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_213 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_107 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_848 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n8) );
  CLKBUF_X1 U4 ( .A(B), .Z(n5) );
  CLKBUF_X1 U5 ( .A(n8), .Z(n6) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_847 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_846 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_845 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_212 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_848 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_847 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_846 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_845 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_844 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_843 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_842 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_841 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_211 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_844 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_843 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_842 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_841 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_106 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U2 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U3 ( .A(sel), .ZN(n5) );
  CLKBUF_X1 U4 ( .A(sel), .Z(n10) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  INV_X1 U7 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n15), .ZN(n17) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
endmodule


module carry_select_block_NPB4_106 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_212 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_211 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_106 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_840 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n8), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  AOI22_X1 U6 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_839 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_838 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_837 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_210 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_840 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_839 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_838 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_837 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_836 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_835 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_834 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_833 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_209 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_836 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_835 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_834 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_833 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_105 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n17), .ZN(Y[2]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n5) );
  INV_X1 U3 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n14), .ZN(n18) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[2]), .B1(n14), .B2(B[2]), .ZN(n17) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[1]), .B1(n14), .B2(B[1]), .ZN(n16) );
  INV_X1 U8 ( .A(sel), .ZN(n14) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[0]), .B1(n14), .B2(B[0]), .ZN(n15) );
  INV_X2 U10 ( .A(n15), .ZN(Y[0]) );
endmodule


module carry_select_block_NPB4_105 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_210 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_209 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_105 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_832 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n4), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_831 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_830 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_829 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_208 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_832 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_831 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_830 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_829 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_828 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_827 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_826 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_825 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_207 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_828 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_827 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_826 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_825 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_104 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n18), .ZN(Y[2]) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n5) );
  INV_X1 U4 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U5 ( .A(sel), .ZN(n10) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U7 ( .A(sel), .ZN(n15) );
  AOI22_X1 U8 ( .A1(n5), .A2(A[3]), .B1(B[3]), .B2(n15), .ZN(n19) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U10 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n10), .ZN(n16) );
endmodule


module carry_select_block_NPB4_104 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_208 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_207 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_104 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_824 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n4), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_823 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68447, n4, n5, n6, n7;
  assign Co = net68447;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  AOI22_X1 U2 ( .A1(n7), .A2(A), .B1(Ci), .B2(n6), .ZN(n5) );
  INV_X1 U5 ( .A(n5), .ZN(net68447) );
  CLKBUF_X1 U6 ( .A(B), .Z(n7) );
endmodule


module FA_822 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_821 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_206 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_824 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_823 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_822 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_821 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_820 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_819 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(n4), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_818 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_817 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_205 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_820 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_819 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_818 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_817 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_103 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n17), .ZN(Y[2]) );
  INV_X2 U2 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U5 ( .A(sel), .ZN(n5) );
  AOI22_X1 U6 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n5), .ZN(n18) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[2]), .B1(n5), .B2(B[2]), .ZN(n17) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[1]), .B1(n5), .B2(B[1]), .ZN(n16) );
  INV_X1 U9 ( .A(sel), .ZN(n14) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n14), .B2(B[0]), .ZN(n15) );
endmodule


module carry_select_block_NPB4_103 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_206 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_205 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_103 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_816 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n8), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_815 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(n7), .Z(S) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(n5), .B(B), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(Ci), .B2(n7), .ZN(n8) );
endmodule


module FA_814 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_813 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_204 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_816 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_815 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_814 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_813 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_812 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_811 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n5) );
  XNOR2_X1 U2 ( .A(n5), .B(B), .ZN(n4) );
  XNOR2_X1 U4 ( .A(n5), .B(B), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_810 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_809 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_203 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_812 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_811 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_810 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_809 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_102 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(sel), .Z(n11) );
  INV_X1 U2 ( .A(sel), .ZN(n5) );
  INV_X1 U3 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U4 ( .A(sel), .ZN(n10) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U7 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n11), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n11), .B1(B[3]), .B2(n10), .ZN(n19) );
  AOI22_X1 U10 ( .A1(A[1]), .A2(n11), .B1(B[1]), .B2(n10), .ZN(n17) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n5), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_102 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_204 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_203 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_102 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_808 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68432, n4, n5, n6, n7;
  assign Co = net68432;

  INV_X1 U1 ( .A(Ci), .ZN(n6) );
  CLKBUF_X1 U2 ( .A(n5), .Z(n4) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n7) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n5) );
  XNOR2_X1 U5 ( .A(Ci), .B(n4), .ZN(S) );
  OAI21_X1 U6 ( .B1(n5), .B2(n6), .A(n7), .ZN(net68432) );
endmodule


module FA_807 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n5), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n8) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n5) );
  CLKBUF_X1 U5 ( .A(n8), .Z(n6) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(Ci), .B2(n8), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_806 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68430, n4, n5;
  assign Co = net68430;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(net68430) );
endmodule


module FA_805 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_202 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_808 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_807 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_806 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_805 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_804 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_803 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_802 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_801 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_201 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_804 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_803 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_802 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_801 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_101 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n17), .ZN(Y[1]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n5) );
  INV_X1 U3 ( .A(sel), .ZN(n10) );
  INV_X1 U4 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U7 ( .A(sel), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n15), .ZN(n19) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n10), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_101 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_202 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_201 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_101 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_800 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(n4), .ZN(n8) );
  CLKBUF_X1 U4 ( .A(B), .Z(n5) );
  XOR2_X1 U5 ( .A(A), .B(n5), .Z(n6) );
  AOI22_X1 U6 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_799 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_798 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_797 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_200 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_800 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_799 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_798 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_797 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_796 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_795 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_794 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_793 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_199 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_796 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_795 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_794 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_793 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_100 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n17), .ZN(Y[1]) );
  BUF_X1 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U4 ( .A(sel), .ZN(n5) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(n10), .A2(A[2]), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n5), .ZN(n17) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
  INV_X1 U9 ( .A(sel), .ZN(n15) );
  INV_X1 U10 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
endmodule


module carry_select_block_NPB4_100 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_200 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_199 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_100 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_792 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_791 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_790 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_789 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_198 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_792 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_791 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_790 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_789 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_788 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_787 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_786 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_785 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_197 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_788 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_787 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_786 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_785 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_99 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  CLKBUF_X1 U1 ( .A(n15), .Z(n5) );
  INV_X1 U2 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(n10) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U6 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(n10), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(n10), .B1(B[1]), .B2(n5), .ZN(n17) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_99 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_198 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_197 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_99 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_784 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_783 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_782 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_781 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_196 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_784 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_783 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_782 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_781 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_780 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_779 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_778 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_777 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_195 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_780 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_779 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_778 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_777 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_98 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X2 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U6 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_98 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_196 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_195 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_98 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_776 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_775 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_774 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_773 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_194 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_776 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_775 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_774 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_773 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_772 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_771 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_770 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_769 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_193 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_772 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_771 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_770 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_769 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_97 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(sel), .ZN(n13) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_97 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_194 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_193 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_97 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_7 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_112 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_111 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_110 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_109 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_108 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_107 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_106 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_105 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_104 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_103 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_102 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), .S(S[43:40]) );
  carry_select_block_NPB4_101 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), .S(S[47:44]) );
  carry_select_block_NPB4_100 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), .S(S[51:48]) );
  carry_select_block_NPB4_99 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), 
        .S(S[55:52]) );
  carry_select_block_NPB4_98 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), 
        .S(S[59:56]) );
  carry_select_block_NPB4_97 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), 
        .S(S[63:60]) );
endmodule


module P4_ADDER_N64_7 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_7 CGEN ( .A(A), .B({B[63:53], n5, B[51:49], n24, 
        B[47:41], n20, B[39:37], n22, B[35:33], n21, B[31:29], n6, B[27:0]}), 
        .Cin(Cin), .Co(CoutCgen) );
  sum_generator_N64_NPB4_7 SGEN ( .A(A), .B({B[63:52], n23, B[50:48], n4, n16, 
        n15, B[44], n7, n9, n11, B[40], n12, n10, B[37:36], n19, B[34:32], n8, 
        n2, B[29:28], n17, B[26:24], n14, B[22:0]}), .Ci({CoutCgen, Cin}), .S(
        S), .Co(Cout) );
  BUF_X1 U1 ( .A(B[41]), .Z(n11) );
  CLKBUF_X1 U2 ( .A(B[23]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(B[30]), .Z(n2) );
  INV_X1 U4 ( .A(B[47]), .ZN(n3) );
  INV_X1 U5 ( .A(n3), .ZN(n4) );
  CLKBUF_X1 U6 ( .A(B[52]), .Z(n5) );
  BUF_X2 U7 ( .A(B[45]), .Z(n15) );
  CLKBUF_X1 U8 ( .A(B[28]), .Z(n6) );
  CLKBUF_X1 U9 ( .A(B[43]), .Z(n7) );
  CLKBUF_X1 U10 ( .A(B[31]), .Z(n8) );
  BUF_X1 U11 ( .A(B[42]), .Z(n9) );
  CLKBUF_X1 U12 ( .A(B[38]), .Z(n10) );
  CLKBUF_X1 U13 ( .A(B[39]), .Z(n12) );
  INV_X1 U14 ( .A(n1), .ZN(n13) );
  INV_X1 U15 ( .A(n13), .ZN(n14) );
  BUF_X1 U16 ( .A(B[46]), .Z(n16) );
  CLKBUF_X1 U17 ( .A(B[27]), .Z(n17) );
  INV_X1 U18 ( .A(B[35]), .ZN(n18) );
  INV_X1 U19 ( .A(n18), .ZN(n19) );
  CLKBUF_X1 U20 ( .A(B[51]), .Z(n23) );
  CLKBUF_X1 U21 ( .A(B[40]), .Z(n20) );
  CLKBUF_X1 U22 ( .A(B[32]), .Z(n21) );
  CLKBUF_X1 U23 ( .A(B[36]), .Z(n22) );
  CLKBUF_X1 U24 ( .A(B[48]), .Z(n24) );
endmodule


module Booth_Encoder_6 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_6 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306;

  NAND2_X1 U1 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  NAND2_X1 U2 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  NAND2_X1 U3 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  NAND2_X1 U4 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  NAND2_X1 U5 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  NAND2_X1 U6 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  NOR3_X1 U7 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U8 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  NAND2_X2 U9 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  BUF_X1 U10 ( .A(n158), .Z(n161) );
  BUF_X1 U11 ( .A(n158), .Z(n160) );
  BUF_X1 U12 ( .A(n158), .Z(n162) );
  BUF_X1 U13 ( .A(n158), .Z(n163) );
  BUF_X1 U14 ( .A(n158), .Z(n159) );
  BUF_X1 U15 ( .A(n151), .Z(n153) );
  BUF_X1 U16 ( .A(n165), .Z(n167) );
  BUF_X1 U17 ( .A(n151), .Z(n154) );
  BUF_X1 U18 ( .A(n303), .Z(n158) );
  NOR4_X1 U19 ( .A1(n150), .A2(n144), .A3(n153), .A4(n167), .ZN(n303) );
  BUF_X1 U20 ( .A(n151), .Z(n155) );
  BUF_X1 U21 ( .A(n152), .Z(n156) );
  BUF_X1 U22 ( .A(n165), .Z(n169) );
  BUF_X1 U23 ( .A(n166), .Z(n170) );
  BUF_X1 U24 ( .A(n165), .Z(n168) );
  BUF_X1 U25 ( .A(n152), .Z(n157) );
  BUF_X1 U26 ( .A(n166), .Z(n171) );
  BUF_X1 U27 ( .A(n304), .Z(n165) );
  BUF_X1 U28 ( .A(n302), .Z(n151) );
  BUF_X1 U29 ( .A(n301), .Z(n148) );
  BUF_X1 U30 ( .A(n301), .Z(n147) );
  BUF_X1 U31 ( .A(n301), .Z(n149) );
  BUF_X1 U32 ( .A(n301), .Z(n146) );
  BUF_X1 U33 ( .A(n304), .Z(n166) );
  BUF_X1 U34 ( .A(n302), .Z(n152) );
  BUF_X1 U35 ( .A(n301), .Z(n145) );
  BUF_X1 U36 ( .A(n300), .Z(n142) );
  BUF_X1 U37 ( .A(n300), .Z(n139) );
  BUF_X1 U38 ( .A(n300), .Z(n141) );
  BUF_X1 U39 ( .A(n300), .Z(n143) );
  BUF_X1 U40 ( .A(n300), .Z(n140) );
  INV_X1 U41 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U42 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n304) );
  AND3_X1 U43 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U44 ( .A(sel[2]), .ZN(n173) );
  NAND2_X1 U45 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI22_X1 U46 ( .A1(C[22]), .A2(n149), .B1(A[22]), .B2(n143), .ZN(n203) );
  NAND2_X1 U47 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI22_X1 U48 ( .A1(C[23]), .A2(n149), .B1(A[23]), .B2(n143), .ZN(n205) );
  NAND2_X1 U49 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI22_X1 U50 ( .A1(C[25]), .A2(n148), .B1(A[25]), .B2(n142), .ZN(n209) );
  AOI22_X1 U51 ( .A1(C[24]), .A2(n149), .B1(A[24]), .B2(n143), .ZN(n207) );
  NAND2_X1 U52 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI22_X1 U53 ( .A1(C[54]), .A2(n146), .B1(A[54]), .B2(n140), .ZN(n273) );
  AOI222_X1 U54 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n156), .ZN(n272) );
  NAND2_X1 U55 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI22_X1 U56 ( .A1(C[27]), .A2(n148), .B1(A[27]), .B2(n142), .ZN(n213) );
  AOI222_X1 U57 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n154), .ZN(n212) );
  NAND2_X1 U58 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI22_X1 U59 ( .A1(C[31]), .A2(n148), .B1(A[31]), .B2(n142), .ZN(n223) );
  AOI222_X1 U60 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n154), .ZN(n222) );
  NAND2_X1 U61 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI22_X1 U62 ( .A1(C[26]), .A2(n148), .B1(A[26]), .B2(n142), .ZN(n211) );
  AOI222_X1 U63 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n154), .ZN(n210) );
  NAND2_X1 U64 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI22_X1 U65 ( .A1(C[39]), .A2(n147), .B1(A[39]), .B2(n141), .ZN(n239) );
  AOI222_X1 U66 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n155), .ZN(n238) );
  AOI22_X1 U67 ( .A1(C[44]), .A2(n147), .B1(A[44]), .B2(n141), .ZN(n251) );
  AOI222_X1 U68 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n156), .ZN(n250) );
  AOI22_X1 U69 ( .A1(C[40]), .A2(n147), .B1(A[40]), .B2(n141), .ZN(n243) );
  AOI222_X1 U70 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n155), .ZN(n242) );
  NAND2_X1 U71 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  AOI22_X1 U72 ( .A1(C[36]), .A2(n147), .B1(A[36]), .B2(n141), .ZN(n233) );
  AOI222_X1 U73 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n155), .ZN(n232) );
  NAND2_X1 U74 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  AOI22_X1 U75 ( .A1(C[53]), .A2(n146), .B1(A[53]), .B2(n140), .ZN(n271) );
  AOI222_X1 U76 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n156), .ZN(n270) );
  AOI222_X1 U77 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n156), .ZN(n258) );
  NAND2_X1 U78 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI22_X1 U79 ( .A1(C[29]), .A2(n148), .B1(A[29]), .B2(n142), .ZN(n217) );
  AOI222_X1 U80 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n154), .ZN(n216) );
  NAND2_X1 U81 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI222_X1 U82 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n156), .ZN(n252) );
  AOI22_X1 U83 ( .A1(C[45]), .A2(n147), .B1(A[45]), .B2(n141), .ZN(n253) );
  NAND2_X1 U84 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI222_X1 U85 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n156), .ZN(n260) );
  AOI22_X1 U86 ( .A1(C[49]), .A2(n146), .B1(A[49]), .B2(n140), .ZN(n261) );
  NAND2_X1 U87 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U88 ( .A1(C[30]), .A2(n148), .B1(A[30]), .B2(n142), .ZN(n221) );
  AOI222_X1 U89 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n154), .ZN(n220) );
  NAND2_X1 U90 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI22_X1 U91 ( .A1(C[38]), .A2(n147), .B1(A[38]), .B2(n141), .ZN(n237) );
  AOI222_X1 U92 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n155), .ZN(n236) );
  NAND2_X1 U93 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI22_X1 U94 ( .A1(C[42]), .A2(n147), .B1(A[42]), .B2(n141), .ZN(n247) );
  AOI222_X1 U95 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n155), .ZN(n246) );
  NAND2_X1 U96 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI22_X1 U97 ( .A1(C[46]), .A2(n146), .B1(A[46]), .B2(n140), .ZN(n255) );
  AOI222_X1 U98 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n156), .ZN(n254) );
  NAND2_X1 U99 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI22_X1 U100 ( .A1(C[50]), .A2(n146), .B1(A[50]), .B2(n140), .ZN(n265) );
  AOI222_X1 U101 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n156), .ZN(n264) );
  NAND2_X1 U102 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI222_X1 U103 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n155), .ZN(n248) );
  NAND2_X1 U104 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI222_X1 U105 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n156), .ZN(n256) );
  NAND2_X1 U106 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI222_X1 U107 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n155), .ZN(n244) );
  AOI22_X1 U108 ( .A1(C[41]), .A2(n147), .B1(A[41]), .B2(n141), .ZN(n245) );
  AOI22_X1 U109 ( .A1(C[28]), .A2(n148), .B1(A[28]), .B2(n142), .ZN(n215) );
  AOI222_X1 U110 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n154), .ZN(n214) );
  NAND2_X1 U111 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  AOI222_X1 U112 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n156), .ZN(n266) );
  NAND2_X1 U113 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI22_X1 U114 ( .A1(C[55]), .A2(n146), .B1(A[55]), .B2(n140), .ZN(n275) );
  AOI222_X1 U115 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n156), .ZN(n274) );
  NAND2_X1 U116 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  AOI222_X1 U117 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n156), .ZN(n268) );
  AOI22_X1 U118 ( .A1(C[52]), .A2(n146), .B1(A[52]), .B2(n140), .ZN(n269) );
  AOI222_X1 U119 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n154), .ZN(n198) );
  AOI22_X1 U120 ( .A1(C[32]), .A2(n148), .B1(A[32]), .B2(n142), .ZN(n225) );
  AOI222_X1 U121 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n155), .ZN(n224) );
  NAND2_X1 U122 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U123 ( .A1(C[60]), .A2(n145), .B1(A[60]), .B2(n139), .ZN(n287) );
  AOI222_X1 U124 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n157), .ZN(n286) );
  NAND2_X1 U125 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  AOI22_X1 U126 ( .A1(C[57]), .A2(n145), .B1(A[57]), .B2(n139), .ZN(n279) );
  AOI222_X1 U127 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n157), .ZN(n278) );
  NAND2_X1 U128 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U129 ( .A1(C[61]), .A2(n145), .B1(A[61]), .B2(n139), .ZN(n289) );
  AOI222_X1 U130 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n157), .ZN(n288) );
  NAND2_X1 U131 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U132 ( .A1(C[59]), .A2(n145), .B1(A[59]), .B2(n139), .ZN(n283) );
  AOI222_X1 U133 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n157), .ZN(n282) );
  NAND2_X1 U134 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI22_X1 U135 ( .A1(C[35]), .A2(n148), .B1(A[35]), .B2(n142), .ZN(n231) );
  AOI222_X1 U136 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n155), .ZN(n230) );
  NAND2_X1 U137 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI222_X1 U138 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n155), .ZN(n226) );
  AOI22_X1 U139 ( .A1(C[33]), .A2(n148), .B1(A[33]), .B2(n142), .ZN(n227) );
  NAND2_X1 U140 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI22_X1 U141 ( .A1(C[34]), .A2(n148), .B1(A[34]), .B2(n142), .ZN(n229) );
  AOI222_X1 U142 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n155), .ZN(n228) );
  AOI22_X1 U143 ( .A1(C[56]), .A2(n146), .B1(A[56]), .B2(n140), .ZN(n277) );
  AOI222_X1 U144 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n157), .ZN(n276) );
  NAND2_X1 U145 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI22_X1 U146 ( .A1(C[58]), .A2(n145), .B1(A[58]), .B2(n139), .ZN(n281) );
  AOI222_X1 U147 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n157), .ZN(n280) );
  NAND2_X1 U148 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI222_X1 U149 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n155), .ZN(n234) );
  AOI22_X1 U150 ( .A1(C[37]), .A2(n147), .B1(A[37]), .B2(n141), .ZN(n235) );
  NAND2_X1 U151 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U152 ( .A1(C[62]), .A2(n145), .B1(A[62]), .B2(n139), .ZN(n291) );
  AOI222_X1 U153 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n157), .ZN(n290) );
  NAND2_X1 U154 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U155 ( .A1(C[63]), .A2(n145), .B1(A[63]), .B2(n139), .ZN(n293) );
  AOI222_X1 U156 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n157), .ZN(n292) );
  NAND2_X1 U157 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U158 ( .A1(C[0]), .A2(n145), .B1(A[0]), .B2(n139), .ZN(n175) );
  AOI222_X1 U159 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n153), .ZN(n174) );
  NAND2_X1 U160 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U161 ( .A1(C[4]), .A2(n146), .B1(A[4]), .B2(n140), .ZN(n263) );
  AOI222_X1 U162 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n156), .ZN(n262) );
  NAND2_X1 U163 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI22_X1 U164 ( .A1(C[8]), .A2(n145), .B1(A[8]), .B2(n139), .ZN(n299) );
  AOI222_X1 U165 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n157), .ZN(n298) );
  NAND2_X1 U166 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  AOI22_X1 U167 ( .A1(C[12]), .A2(n150), .B1(A[12]), .B2(n144), .ZN(n181) );
  AOI222_X1 U168 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n153), .ZN(n180) );
  NAND2_X1 U169 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  AOI22_X1 U170 ( .A1(C[16]), .A2(n149), .B1(A[16]), .B2(n143), .ZN(n189) );
  AOI222_X1 U171 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n153), .ZN(n188) );
  NAND2_X1 U172 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U173 ( .A1(C[1]), .A2(n149), .B1(A[1]), .B2(n143), .ZN(n197) );
  AOI222_X1 U174 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n153), .ZN(n196) );
  NAND2_X1 U175 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U176 ( .A1(C[5]), .A2(n145), .B1(A[5]), .B2(n139), .ZN(n285) );
  AOI222_X1 U177 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n157), .ZN(n284) );
  NAND2_X1 U178 ( .A1(n306), .A2(n305), .ZN(Y[9]) );
  AOI22_X1 U179 ( .A1(C[9]), .A2(n147), .B1(A[9]), .B2(n141), .ZN(n306) );
  AOI222_X1 U180 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n157), .ZN(n305) );
  NAND2_X1 U181 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U182 ( .A1(C[13]), .A2(n150), .B1(A[13]), .B2(n144), .ZN(n183) );
  AOI222_X1 U183 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n153), .ZN(n182) );
  NAND2_X1 U184 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI22_X1 U185 ( .A1(C[17]), .A2(n149), .B1(A[17]), .B2(n143), .ZN(n191) );
  AOI222_X1 U186 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n153), .ZN(n190) );
  NAND2_X1 U187 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U188 ( .A1(C[2]), .A2(n148), .B1(A[2]), .B2(n142), .ZN(n219) );
  AOI222_X1 U189 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n154), .ZN(n218) );
  NAND2_X1 U190 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U191 ( .A1(C[6]), .A2(n145), .B1(A[6]), .B2(n139), .ZN(n295) );
  AOI222_X1 U192 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n157), .ZN(n294) );
  NAND2_X1 U193 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U194 ( .A1(C[10]), .A2(n150), .B1(A[10]), .B2(n144), .ZN(n177) );
  AOI222_X1 U195 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n153), .ZN(n176) );
  NAND2_X1 U196 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U197 ( .A1(C[14]), .A2(n149), .B1(A[14]), .B2(n143), .ZN(n185) );
  AOI222_X1 U198 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n153), .ZN(n184) );
  NAND2_X1 U199 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI22_X1 U200 ( .A1(C[18]), .A2(n149), .B1(A[18]), .B2(n143), .ZN(n193) );
  AOI222_X1 U201 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n153), .ZN(n192) );
  NAND2_X1 U202 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U203 ( .A1(C[3]), .A2(n147), .B1(A[3]), .B2(n141), .ZN(n241) );
  AOI222_X1 U204 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n155), .ZN(n240) );
  NAND2_X1 U205 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U206 ( .A1(C[7]), .A2(n145), .B1(A[7]), .B2(n139), .ZN(n297) );
  AOI222_X1 U207 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n157), .ZN(n296) );
  NAND2_X1 U208 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U209 ( .A1(C[11]), .A2(n150), .B1(A[11]), .B2(n144), .ZN(n179) );
  AOI222_X1 U210 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n153), .ZN(n178) );
  NAND2_X1 U211 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U212 ( .A1(C[15]), .A2(n149), .B1(A[15]), .B2(n143), .ZN(n187) );
  AOI222_X1 U213 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n153), .ZN(n186) );
  NAND2_X1 U214 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI22_X1 U215 ( .A1(C[19]), .A2(n149), .B1(A[19]), .B2(n143), .ZN(n195) );
  AOI222_X1 U216 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n153), .ZN(n194) );
  AOI22_X1 U217 ( .A1(C[48]), .A2(n146), .B1(A[48]), .B2(n140), .ZN(n259) );
  AOI22_X1 U218 ( .A1(C[47]), .A2(n146), .B1(A[47]), .B2(n140), .ZN(n257) );
  AOI22_X1 U219 ( .A1(C[20]), .A2(n149), .B1(A[20]), .B2(n143), .ZN(n199) );
  AOI22_X1 U220 ( .A1(C[21]), .A2(n149), .B1(A[21]), .B2(n143), .ZN(n201) );
  NAND2_X1 U221 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  NAND2_X1 U222 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI222_X1 U223 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n154), .ZN(n208) );
  AOI222_X1 U224 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n154), .ZN(n206) );
  AOI22_X1 U225 ( .A1(C[43]), .A2(n147), .B1(A[43]), .B2(n141), .ZN(n249) );
  AOI222_X1 U226 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n154), .ZN(n200) );
  AOI22_X1 U227 ( .A1(C[51]), .A2(n146), .B1(A[51]), .B2(n140), .ZN(n267) );
  AOI222_X1 U228 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n154), .ZN(n202) );
  AOI222_X1 U229 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n154), .ZN(n204) );
  CLKBUF_X1 U230 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U231 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U232 ( .A(n158), .Z(n164) );
endmodule


module G_102 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_378 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_377 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_376 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_375 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_374 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_373 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_372 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_371 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_370 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_369 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_368 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3, n5;

  CLKBUF_X1 U1 ( .A(P_IK), .Z(n3) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n5) );
  AND2_X1 U3 ( .A1(n3), .A2(P_K_1), .ZN(Px) );
  INV_X1 U4 ( .A(n5), .ZN(Gx) );
endmodule


module PG_367 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_366 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_365 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_364 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_363 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_362 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_361 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_360 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_359 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_358 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_357 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_356 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_355 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_354 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_353 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_352 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_351 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_350 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_349 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_348 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_101 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_347 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_346 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_345 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_344 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_343 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_342 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_341 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_340 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_339 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_338 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_337 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_336 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_335 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_334 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_333 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_100 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_332 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_331 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_330 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_329 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_328 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_327 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_326 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_99 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_98 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_325 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_324 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_323 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  OR2_X2 U2 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_322 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_321 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_320 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_97 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_96 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_95 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n3, n5;

  AND2_X1 U1 ( .A1(P_IK), .A2(G_K_1), .ZN(n3) );
  NOR2_X1 U2 ( .A1(n3), .A2(G_IK), .ZN(n5) );
  INV_X1 U3 ( .A(n5), .ZN(Gx) );
endmodule


module G_94 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_319 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_318 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_317 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_316 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module G_93 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_92 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_91 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_90 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_89 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_88 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n3;

  AND2_X1 U1 ( .A1(P_IK), .A2(G_K_1), .ZN(n3) );
  OR2_X2 U2 ( .A1(G_IK), .A2(n3), .ZN(Gx) );
endmodule


module G_87 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_86 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module carry_generator_N64_NPB4_6 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U88 ( .A(B[49]), .B(A[49]), .Z(\PG_Network[0][0][49] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U91 ( .A(B[46]), .B(A[46]), .Z(\PG_Network[0][0][46] ) );
  XOR2_X1 U92 ( .A(B[45]), .B(A[45]), .Z(\PG_Network[0][0][45] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U101 ( .A(B[37]), .B(A[37]), .Z(\PG_Network[0][0][37] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U108 ( .A(B[30]), .B(A[30]), .Z(\PG_Network[0][0][30] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U114 ( .A(B[25]), .B(A[25]), .Z(\PG_Network[0][0][25] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U121 ( .A(B[19]), .B(A[19]), .Z(\PG_Network[0][0][19] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U125 ( .A(B[15]), .B(A[15]), .Z(\PG_Network[0][0][15] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_102 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n25), .Gx(\PG_Network[1][1][1] ) );
  PG_378 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_377 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_376 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_375 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_374 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_373 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_372 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_371 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_370 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_369 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_368 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_367 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_366 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_365 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_364 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_363 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_362 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_361 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_360 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_359 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_358 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_357 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_356 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_355 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_354 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_353 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_352 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_351 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_350 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_349 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_348 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_101 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_347 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_346 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_345 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_344 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_343 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_342 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_341 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_340 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_339 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_338 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_337 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_336 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_335 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_334 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_333 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_100 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_332 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_331 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_330 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_329 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_328 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_327 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_326 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_99 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), 
        .G_K_1(Co[1]), .Gx(Co[3]) );
  G_98 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), 
        .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_325 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_324 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_323 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][47] ), .Px(
        \PG_Network[4][0][47] ) );
  PG_322 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][43] ), .Px(
        \PG_Network[4][0][43] ) );
  PG_321 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(n15), .P_K_1(\PG_Network[3][0][55] ), 
        .Gx(\PG_Network[4][1][63] ), .Px(\PG_Network[4][0][63] ) );
  PG_320 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(n15), .P_K_1(\PG_Network[3][0][55] ), 
        .Gx(\PG_Network[4][1][59] ), .Px(\PG_Network[4][0][59] ) );
  G_97 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), 
        .G_K_1(Co[3]), .Gx(Co[7]) );
  G_96 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), 
        .G_K_1(Co[3]), .Gx(Co[6]) );
  G_95 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), 
        .G_K_1(Co[3]), .Gx(Co[5]) );
  G_94 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), 
        .G_K_1(Co[3]), .Gx(Co[4]) );
  PG_319 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(n24), .P_K_1(n9), .Gx(
        \PG_Network[5][1][63] ), .Px(\PG_Network[5][0][63] ) );
  PG_318 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(n24), .P_K_1(n9), .Gx(
        \PG_Network[5][1][59] ), .Px(\PG_Network[5][0][59] ) );
  PG_317 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(n24), .P_K_1(n11), .Gx(
        \PG_Network[5][1][55] ), .Px(\PG_Network[5][0][55] ) );
  PG_316 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(n11), 
        .Gx(\PG_Network[5][1][51] ), .Px(\PG_Network[5][0][51] ) );
  G_93 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), 
        .G_K_1(n13), .Gx(Co[15]) );
  G_92 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), 
        .G_K_1(n13), .Gx(Co[14]) );
  G_91 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), 
        .G_K_1(n13), .Gx(Co[13]) );
  G_90 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), 
        .G_K_1(n8), .Gx(Co[12]) );
  G_89 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), 
        .G_K_1(n13), .Gx(Co[11]) );
  G_88 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), 
        .G_K_1(n8), .Gx(Co[10]) );
  G_87 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), 
        .G_K_1(n12), .Gx(Co[9]) );
  G_86 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), 
        .G_K_1(Co[7]), .Gx(Co[8]) );
  CLKBUF_X1 U1 ( .A(B[46]), .Z(n5) );
  INV_X1 U2 ( .A(A[29]), .ZN(n7) );
  INV_X1 U3 ( .A(A[38]), .ZN(n6) );
  INV_X1 U4 ( .A(A[59]), .ZN(n10) );
  INV_X1 U5 ( .A(A[23]), .ZN(n14) );
  INV_X1 U6 ( .A(A[27]), .ZN(n16) );
  INV_X1 U7 ( .A(A[31]), .ZN(n20) );
  INV_X1 U8 ( .A(A[39]), .ZN(n21) );
  INV_X1 U9 ( .A(A[43]), .ZN(n19) );
  INV_X1 U10 ( .A(A[47]), .ZN(n22) );
  INV_X1 U11 ( .A(A[51]), .ZN(n23) );
  INV_X1 U12 ( .A(A[35]), .ZN(n18) );
  INV_X1 U13 ( .A(A[55]), .ZN(n17) );
  XNOR2_X1 U14 ( .A(B[38]), .B(n6), .ZN(\PG_Network[0][0][38] ) );
  XNOR2_X1 U15 ( .A(B[29]), .B(n7), .ZN(\PG_Network[0][0][29] ) );
  CLKBUF_X1 U16 ( .A(Co[7]), .Z(n8) );
  CLKBUF_X1 U17 ( .A(n11), .Z(n9) );
  XNOR2_X1 U18 ( .A(B[59]), .B(n10), .ZN(\PG_Network[0][0][59] ) );
  BUF_X1 U19 ( .A(\PG_Network[4][0][47] ), .Z(n11) );
  CLKBUF_X1 U20 ( .A(Co[7]), .Z(n13) );
  CLKBUF_X1 U21 ( .A(Co[7]), .Z(n12) );
  XNOR2_X1 U22 ( .A(B[23]), .B(n14), .ZN(\PG_Network[0][0][23] ) );
  CLKBUF_X1 U23 ( .A(\PG_Network[3][1][55] ), .Z(n15) );
  XNOR2_X1 U24 ( .A(B[27]), .B(n16), .ZN(\PG_Network[0][0][27] ) );
  XNOR2_X1 U25 ( .A(B[55]), .B(n17), .ZN(\PG_Network[0][0][55] ) );
  XNOR2_X1 U26 ( .A(B[35]), .B(n18), .ZN(\PG_Network[0][0][35] ) );
  XNOR2_X1 U27 ( .A(B[43]), .B(n19), .ZN(\PG_Network[0][0][43] ) );
  XNOR2_X1 U28 ( .A(B[31]), .B(n20), .ZN(\PG_Network[0][0][31] ) );
  XNOR2_X1 U29 ( .A(B[39]), .B(n21), .ZN(\PG_Network[0][0][39] ) );
  XNOR2_X1 U30 ( .A(B[47]), .B(n22), .ZN(\PG_Network[0][0][47] ) );
  XNOR2_X1 U31 ( .A(B[51]), .B(n23), .ZN(\PG_Network[0][0][51] ) );
  CLKBUF_X1 U32 ( .A(\PG_Network[4][1][47] ), .Z(n24) );
  AND2_X1 U33 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U34 ( .A1(A[59]), .A2(B[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U35 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U36 ( .A1(A[46]), .A2(n5), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U37 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U38 ( .A1(A[49]), .A2(B[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U39 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U40 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U41 ( .A1(B[31]), .A2(A[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U42 ( .A1(A[25]), .A2(B[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U43 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U44 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U45 ( .A1(B[27]), .A2(A[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U46 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U47 ( .A1(B[35]), .A2(A[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U48 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U49 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U50 ( .A1(A[41]), .A2(B[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U51 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U52 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U53 ( .A1(A[45]), .A2(B[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U54 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
  AND2_X1 U55 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U56 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AND2_X1 U57 ( .A1(B[23]), .A2(A[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U58 ( .A1(A[53]), .A2(B[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U59 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U60 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U61 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U62 ( .A1(B[37]), .A2(A[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U63 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U64 ( .A1(A[29]), .A2(B[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U65 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U66 ( .A1(A[21]), .A2(B[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U67 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U77 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U81 ( .A1(A[11]), .A2(B[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U85 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U90 ( .A1(A[15]), .A2(B[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U94 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U99 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U100 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U103 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U107 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U110 ( .A1(A[19]), .A2(B[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U112 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U116 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U131 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U132 ( .A(n28), .ZN(n25) );
  AND2_X1 U133 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U134 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U135 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U136 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U137 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U138 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U139 ( .A1(A[7]), .A2(B[7]), .ZN(\PG_Network[0][1][7] ) );
  AND2_X1 U140 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U141 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AOI21_X1 U142 ( .B1(A[0]), .B2(B[0]), .A(n26), .ZN(n28) );
  INV_X1 U143 ( .A(n27), .ZN(n26) );
  OAI21_X1 U144 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n27) );
  AND2_X1 U145 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U146 ( .A1(B[43]), .A2(A[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U147 ( .A1(B[47]), .A2(A[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U148 ( .A1(B[51]), .A2(A[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U149 ( .A1(A[55]), .A2(B[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U150 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
endmodule


module FA_768 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_767 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_766 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_765 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_192 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_768 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_767 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_766 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_765 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_764 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_763 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_762 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_761 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_191 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_764 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_763 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_762 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_761 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_96 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U2 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_96 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_192 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_191 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_96 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_760 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_759 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_758 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_757 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_190 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_760 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_759 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_758 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_757 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_756 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_755 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_754 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_753 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_189 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_756 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_755 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_754 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_753 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_95 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_95 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_190 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_189 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_95 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_752 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_751 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_750 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_749 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_188 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_752 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_751 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_750 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_749 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_748 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_747 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_746 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_745 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_187 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_748 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_747 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_746 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_745 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_94 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_94 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_188 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_187 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_94 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_744 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_743 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_742 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_741 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_186 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_744 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_743 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_742 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_741 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_740 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_739 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_738 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_737 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_185 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_740 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_739 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_738 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_737 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_93 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_93 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_186 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_185 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_93 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_736 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_735 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_734 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_733 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_184 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_736 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_735 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_734 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_733 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_732 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_731 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_730 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_729 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_183 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_732 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_731 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_730 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_729 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_92 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_92 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_184 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_183 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_92 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_728 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_727 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_726 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_725 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_182 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_728 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_727 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_726 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_725 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_724 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_723 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_722 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_721 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_181 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_724 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_723 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_722 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_721 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_91 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_91 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_182 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_181 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_91 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_720 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6, n7, n8;

  XOR2_X1 U3 ( .A(n8), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n5) );
  OR2_X1 U2 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n8) );
  AND2_X1 U5 ( .A1(B), .A2(A), .ZN(n6) );
  AND2_X1 U6 ( .A1(n8), .A2(Ci), .ZN(n7) );
endmodule


module FA_719 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_718 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_717 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_180 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_720 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_719 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_718 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_717 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_716 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_715 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_714 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_713 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_179 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_716 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_715 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_714 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_713 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_90 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[0]) );
  CLKBUF_X1 U4 ( .A(sel), .Z(n5) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U6 ( .A(sel), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n14), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n14), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
endmodule


module carry_select_block_NPB4_90 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_180 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_179 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_90 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_712 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_711 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_710 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_709 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_178 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_712 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_711 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_710 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_709 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_708 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_707 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_706 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_705 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_177 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_708 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_707 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_706 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_705 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_89 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U5 ( .A(sel), .ZN(n5) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n16) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n5), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n5), .ZN(n14) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n5), .ZN(n17) );
endmodule


module carry_select_block_NPB4_89 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_178 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_177 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_89 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_704 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_703 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_702 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_701 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_176 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_704 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_703 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_702 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_701 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_700 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_699 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_698 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_697 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_175 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_700 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_699 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_698 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_697 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_88 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U6 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n13), .ZN(n17) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_88 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_176 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_175 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_88 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_696 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68320, n4, n5, n6, n7;
  assign Co = net68320;

  INV_X1 U1 ( .A(Ci), .ZN(n6) );
  CLKBUF_X1 U2 ( .A(n5), .Z(n4) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n7) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n5) );
  XNOR2_X1 U5 ( .A(Ci), .B(n4), .ZN(S) );
  OAI21_X1 U6 ( .B1(n5), .B2(n6), .A(n7), .ZN(net68320) );
endmodule


module FA_695 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n4) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n4), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_694 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68318, n4, n5;
  assign Co = net68318;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(net68318) );
endmodule


module FA_693 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_174 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_696 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_695 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_694 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_693 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_692 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_691 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  BUF_X1 U1 ( .A(B), .Z(n4) );
  XOR2_X1 U2 ( .A(A), .B(n4), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_690 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_689 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_173 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_692 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_691 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_690 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_689 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_87 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[0]) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n5) );
  INV_X1 U4 ( .A(sel), .ZN(n10) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U6 ( .A(n17), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n10), .ZN(n17) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n10), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n10), .ZN(n18) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n10), .B2(B[0]), .ZN(n15) );
endmodule


module carry_select_block_NPB4_87 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_174 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_173 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_87 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_688 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n8), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_687 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_686 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_685 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n8, n10, n11;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n5), .ZN(n4) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n5), .A2(n10), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n7), .A2(n8), .ZN(S) );
  INV_X1 U6 ( .A(Ci), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(n6) );
  INV_X1 U8 ( .A(n11), .ZN(Co) );
  AOI22_X1 U9 ( .A1(B), .A2(A), .B1(n10), .B2(n4), .ZN(n11) );
endmodule


module RCA_N4_172 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_688 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_687 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_686 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_685 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_684 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_683 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  XOR2_X1 U2 ( .A(A), .B(n4), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_682 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_681 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_171 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_684 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_683 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_682 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_681 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_86 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19, n20;

  INV_X1 U1 ( .A(n17), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n11), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n10) );
  CLKBUF_X1 U4 ( .A(sel), .Z(n11) );
  INV_X1 U5 ( .A(n18), .ZN(Y[1]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[2]) );
  INV_X1 U7 ( .A(n20), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n16), .ZN(n20) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(n11), .B1(n5), .B2(B[2]), .ZN(n19) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[1]), .B1(n16), .B2(B[1]), .ZN(n18) );
  INV_X1 U11 ( .A(sel), .ZN(n16) );
  AOI22_X1 U12 ( .A1(sel), .A2(A[0]), .B1(n16), .B2(B[0]), .ZN(n17) );
endmodule


module carry_select_block_NPB4_86 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_172 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_171 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_86 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_680 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(n4), .ZN(n8) );
  CLKBUF_X1 U4 ( .A(B), .Z(n5) );
  XOR2_X1 U5 ( .A(A), .B(n5), .Z(n6) );
  AOI22_X1 U6 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_679 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_678 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_677 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  OR2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n7) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n7), .A2(n6), .ZN(S) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(n4), .ZN(n10) );
endmodule


module RCA_N4_170 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_680 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_679 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_678 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_677 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_676 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_675 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_674 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_673 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_169 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_676 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_675 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_674 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_673 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_85 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n12, n17, n18, n19, n20, n21;

  BUF_X1 U1 ( .A(n12), .Z(n5) );
  BUF_X1 U2 ( .A(sel), .Z(n11) );
  INV_X1 U3 ( .A(n18), .ZN(Y[0]) );
  CLKBUF_X1 U4 ( .A(sel), .Z(n10) );
  INV_X1 U5 ( .A(n20), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[1]) );
  INV_X1 U7 ( .A(sel), .ZN(n12) );
  INV_X1 U8 ( .A(n21), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(n10), .A2(A[2]), .B1(n5), .B2(B[2]), .ZN(n20) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n11), .B1(n12), .B2(B[3]), .ZN(n21) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[1]), .B1(n12), .B2(B[1]), .ZN(n19) );
  AOI22_X1 U12 ( .A1(sel), .A2(A[0]), .B1(n17), .B2(B[0]), .ZN(n18) );
  INV_X1 U13 ( .A(sel), .ZN(n17) );
endmodule


module carry_select_block_NPB4_85 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_170 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_169 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_85 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_672 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n8), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_671 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_670 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_669 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_168 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_672 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_671 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_670 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_669 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_668 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_667 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_666 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_665 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_167 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_668 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_667 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_666 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_665 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_84 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19, n20;

  INV_X1 U1 ( .A(n16), .ZN(n5) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n11) );
  INV_X1 U3 ( .A(n17), .ZN(Y[0]) );
  INV_X1 U4 ( .A(sel), .ZN(n10) );
  INV_X1 U5 ( .A(n19), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n11), .B1(B[2]), .B2(n16), .ZN(n19) );
  INV_X1 U7 ( .A(n18), .ZN(Y[1]) );
  INV_X1 U8 ( .A(n20), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n16), .ZN(n20) );
  AOI22_X1 U10 ( .A1(n11), .A2(A[1]), .B1(B[1]), .B2(n16), .ZN(n18) );
  INV_X1 U11 ( .A(sel), .ZN(n16) );
  AOI22_X1 U12 ( .A1(sel), .A2(A[0]), .B1(n10), .B2(B[0]), .ZN(n17) );
endmodule


module carry_select_block_NPB4_84 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_168 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_167 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_84 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_664 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_663 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_662 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_661 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_166 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_664 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_663 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_662 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_661 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_660 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_659 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_658 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_657 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module RCA_N4_165 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_660 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_659 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_658 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_657 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_83 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n12, n13, n18, n19, n20, n21;

  INV_X1 U1 ( .A(n20), .ZN(Y[2]) );
  BUF_X1 U2 ( .A(n5), .Z(n10) );
  INV_X2 U3 ( .A(n18), .ZN(Y[0]) );
  BUF_X1 U4 ( .A(sel), .Z(n11) );
  INV_X1 U5 ( .A(sel), .ZN(n5) );
  BUF_X1 U6 ( .A(n10), .Z(n13) );
  CLKBUF_X1 U7 ( .A(n11), .Z(n12) );
  INV_X1 U8 ( .A(n19), .ZN(Y[1]) );
  INV_X1 U9 ( .A(n21), .ZN(Y[3]) );
  AOI22_X1 U10 ( .A1(A[2]), .A2(n12), .B1(B[2]), .B2(n13), .ZN(n20) );
  AOI22_X1 U11 ( .A1(n11), .A2(A[1]), .B1(n10), .B2(B[1]), .ZN(n19) );
  AOI22_X1 U12 ( .A1(A[3]), .A2(n12), .B1(B[3]), .B2(n13), .ZN(n21) );
  AOI22_X1 U13 ( .A1(sel), .A2(A[0]), .B1(n5), .B2(B[0]), .ZN(n18) );
endmodule


module carry_select_block_NPB4_83 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_166 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_165 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_83 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_656 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(n4) );
  NAND2_X1 U2 ( .A1(n8), .A2(Ci), .ZN(n5) );
  AND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(n9) );
  XOR2_X1 U6 ( .A(A), .B(B), .Z(n6) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_655 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_654 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_653 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_164 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_656 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_655 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_654 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_653 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_652 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_651 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_650 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_649 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_163 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_652 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_651 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_650 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_649 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_82 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X2 U1 ( .A(n15), .ZN(Y[0]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n5) );
  INV_X1 U3 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(n5), .A2(A[3]), .B1(B[3]), .B2(n14), .ZN(n18) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n14), .ZN(n17) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(n5), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[0]), .B1(n14), .B2(B[0]), .ZN(n15) );
  INV_X1 U10 ( .A(sel), .ZN(n14) );
endmodule


module carry_select_block_NPB4_82 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_164 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_163 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_82 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_648 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_647 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_646 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_645 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_162 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_648 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_647 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_646 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_645 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_644 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_643 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_642 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_641 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_161 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_644 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_643 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_642 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_641 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_81 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_81 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_162 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_161 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_81 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_6 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_96 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_95 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_94 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_93 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_92 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_91 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_90 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_89 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_88 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_87 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_86 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), 
        .S(S[43:40]) );
  carry_select_block_NPB4_85 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), 
        .S(S[47:44]) );
  carry_select_block_NPB4_84 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), 
        .S(S[51:48]) );
  carry_select_block_NPB4_83 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), 
        .S(S[55:52]) );
  carry_select_block_NPB4_82 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), 
        .S(S[59:56]) );
  carry_select_block_NPB4_81 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), 
        .S(S[63:60]) );
endmodule


module P4_ADDER_N64_6 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_6 CGEN ( .A(A), .B({B[63:53], n18, B[51:49], n15, 
        B[47:45], n4, B[43:41], n17, B[39:33], n8, B[31:25], n9, B[23:0]}), 
        .Cin(Cin), .Co(CoutCgen) );
  sum_generator_N64_NPB4_6 SGEN ( .A(A), .B({B[63:56], n3, B[54:52], n16, 
        B[50:48], n13, n1, B[45:44], n2, B[42:40], n14, n7, n10, B[36], n11, 
        B[34:32], n5, B[30:28], n6, B[26:24], n12, B[22:0]}), .Ci({CoutCgen, 
        Cin}), .S(S), .Co(Cout) );
  BUF_X1 U1 ( .A(B[37]), .Z(n10) );
  BUF_X1 U2 ( .A(B[46]), .Z(n1) );
  BUF_X1 U3 ( .A(B[55]), .Z(n3) );
  CLKBUF_X1 U4 ( .A(B[43]), .Z(n2) );
  CLKBUF_X1 U5 ( .A(B[44]), .Z(n4) );
  CLKBUF_X1 U6 ( .A(B[31]), .Z(n5) );
  CLKBUF_X1 U7 ( .A(B[27]), .Z(n6) );
  CLKBUF_X1 U8 ( .A(B[48]), .Z(n15) );
  CLKBUF_X1 U9 ( .A(B[38]), .Z(n7) );
  CLKBUF_X1 U10 ( .A(B[32]), .Z(n8) );
  CLKBUF_X1 U11 ( .A(B[24]), .Z(n9) );
  CLKBUF_X1 U12 ( .A(B[35]), .Z(n11) );
  CLKBUF_X1 U13 ( .A(B[23]), .Z(n12) );
  CLKBUF_X1 U14 ( .A(B[47]), .Z(n13) );
  CLKBUF_X1 U15 ( .A(B[39]), .Z(n14) );
  CLKBUF_X1 U16 ( .A(B[51]), .Z(n16) );
  CLKBUF_X1 U17 ( .A(B[40]), .Z(n17) );
  CLKBUF_X1 U18 ( .A(B[52]), .Z(n18) );
endmodule


module Booth_Encoder_5 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_5 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306;

  NAND2_X1 U1 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  NAND2_X1 U2 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  NAND2_X1 U3 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  NAND2_X2 U4 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  NOR3_X1 U5 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U6 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  NAND2_X2 U7 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  BUF_X1 U8 ( .A(n158), .Z(n162) );
  BUF_X1 U9 ( .A(n158), .Z(n161) );
  BUF_X1 U10 ( .A(n158), .Z(n160) );
  BUF_X1 U11 ( .A(n158), .Z(n163) );
  BUF_X1 U12 ( .A(n158), .Z(n159) );
  BUF_X1 U13 ( .A(n151), .Z(n153) );
  BUF_X1 U14 ( .A(n151), .Z(n155) );
  BUF_X1 U15 ( .A(n165), .Z(n167) );
  BUF_X1 U16 ( .A(n165), .Z(n169) );
  BUF_X1 U17 ( .A(n151), .Z(n154) );
  BUF_X1 U18 ( .A(n165), .Z(n168) );
  BUF_X1 U19 ( .A(n303), .Z(n158) );
  NOR4_X1 U20 ( .A1(n150), .A2(n144), .A3(n153), .A4(n167), .ZN(n303) );
  BUF_X1 U21 ( .A(n152), .Z(n157) );
  BUF_X1 U22 ( .A(n152), .Z(n156) );
  BUF_X1 U23 ( .A(n166), .Z(n171) );
  BUF_X1 U24 ( .A(n166), .Z(n170) );
  BUF_X1 U25 ( .A(n301), .Z(n148) );
  BUF_X1 U26 ( .A(n301), .Z(n147) );
  BUF_X1 U27 ( .A(n301), .Z(n149) );
  BUF_X1 U28 ( .A(n304), .Z(n165) );
  BUF_X1 U29 ( .A(n302), .Z(n151) );
  BUF_X1 U30 ( .A(n301), .Z(n145) );
  BUF_X1 U31 ( .A(n301), .Z(n146) );
  BUF_X1 U32 ( .A(n304), .Z(n166) );
  BUF_X1 U33 ( .A(n302), .Z(n152) );
  BUF_X1 U34 ( .A(n300), .Z(n142) );
  BUF_X1 U35 ( .A(n300), .Z(n139) );
  BUF_X1 U36 ( .A(n300), .Z(n141) );
  BUF_X1 U37 ( .A(n300), .Z(n143) );
  BUF_X1 U38 ( .A(n300), .Z(n140) );
  INV_X1 U39 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U40 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n304) );
  AND3_X1 U41 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U42 ( .A(sel[2]), .ZN(n173) );
  NAND2_X1 U43 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI22_X1 U44 ( .A1(C[29]), .A2(n148), .B1(A[29]), .B2(n142), .ZN(n217) );
  AOI222_X1 U45 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n154), .ZN(n216) );
  NAND2_X1 U46 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U47 ( .A1(C[30]), .A2(n148), .B1(A[30]), .B2(n142), .ZN(n221) );
  AOI222_X1 U48 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n154), .ZN(n220) );
  AOI222_X1 U49 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n154), .ZN(n204) );
  AOI222_X1 U50 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n154), .ZN(n202) );
  NAND2_X1 U51 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  AOI22_X1 U52 ( .A1(C[24]), .A2(n149), .B1(A[24]), .B2(n143), .ZN(n207) );
  NAND2_X1 U53 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI22_X1 U54 ( .A1(C[25]), .A2(n148), .B1(A[25]), .B2(n142), .ZN(n209) );
  NAND2_X1 U55 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI22_X1 U56 ( .A1(C[26]), .A2(n148), .B1(A[26]), .B2(n142), .ZN(n211) );
  NAND2_X1 U57 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI22_X1 U58 ( .A1(C[27]), .A2(n148), .B1(A[27]), .B2(n142), .ZN(n213) );
  NAND2_X1 U59 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI22_X1 U60 ( .A1(C[34]), .A2(n148), .B1(A[34]), .B2(n142), .ZN(n229) );
  AOI222_X1 U61 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n155), .ZN(n228) );
  NAND2_X1 U62 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  AOI22_X1 U63 ( .A1(C[57]), .A2(n145), .B1(A[57]), .B2(n139), .ZN(n279) );
  AOI222_X1 U64 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n157), .ZN(n278) );
  NAND2_X1 U65 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI22_X1 U66 ( .A1(C[33]), .A2(n148), .B1(A[33]), .B2(n142), .ZN(n227) );
  AOI222_X1 U67 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n155), .ZN(n226) );
  NAND2_X1 U68 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI22_X1 U69 ( .A1(C[37]), .A2(n147), .B1(A[37]), .B2(n141), .ZN(n235) );
  AOI222_X1 U70 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n155), .ZN(n234) );
  NAND2_X1 U71 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI22_X1 U72 ( .A1(C[31]), .A2(n148), .B1(A[31]), .B2(n142), .ZN(n223) );
  AOI222_X1 U73 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n154), .ZN(n222) );
  NAND2_X1 U74 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI222_X1 U75 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n155), .ZN(n238) );
  AOI22_X1 U76 ( .A1(C[39]), .A2(n147), .B1(A[39]), .B2(n141), .ZN(n239) );
  AOI22_X1 U77 ( .A1(C[28]), .A2(n148), .B1(A[28]), .B2(n142), .ZN(n215) );
  AOI222_X1 U78 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n154), .ZN(n214) );
  NAND2_X1 U79 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  AOI22_X1 U80 ( .A1(C[32]), .A2(n148), .B1(A[32]), .B2(n142), .ZN(n225) );
  AOI222_X1 U81 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n155), .ZN(n224) );
  AOI22_X1 U82 ( .A1(C[36]), .A2(n147), .B1(A[36]), .B2(n141), .ZN(n233) );
  AOI222_X1 U83 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n155), .ZN(n232) );
  NAND2_X1 U84 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI222_X1 U85 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n156), .ZN(n252) );
  NAND2_X1 U86 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI222_X1 U87 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n156), .ZN(n260) );
  NAND2_X1 U88 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI22_X1 U89 ( .A1(C[46]), .A2(n146), .B1(A[46]), .B2(n140), .ZN(n255) );
  AOI222_X1 U90 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n156), .ZN(n254) );
  NAND2_X1 U91 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI22_X1 U92 ( .A1(C[38]), .A2(n147), .B1(A[38]), .B2(n141), .ZN(n237) );
  AOI222_X1 U93 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n155), .ZN(n236) );
  NAND2_X1 U94 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI22_X1 U95 ( .A1(C[42]), .A2(n147), .B1(A[42]), .B2(n141), .ZN(n247) );
  AOI222_X1 U96 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n155), .ZN(n246) );
  NAND2_X1 U97 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI222_X1 U98 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n156), .ZN(n272) );
  AOI22_X1 U99 ( .A1(C[54]), .A2(n146), .B1(A[54]), .B2(n140), .ZN(n273) );
  NAND2_X1 U100 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI22_X1 U101 ( .A1(C[58]), .A2(n145), .B1(A[58]), .B2(n139), .ZN(n281) );
  AOI222_X1 U102 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n157), .ZN(n280) );
  NAND2_X1 U103 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U104 ( .A1(C[59]), .A2(n145), .B1(A[59]), .B2(n139), .ZN(n283) );
  AOI222_X1 U105 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n157), .ZN(n282) );
  NAND2_X1 U106 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI222_X1 U107 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n156), .ZN(n264) );
  AOI22_X1 U108 ( .A1(C[40]), .A2(n147), .B1(A[40]), .B2(n141), .ZN(n243) );
  AOI222_X1 U109 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n155), .ZN(n242) );
  AOI22_X1 U110 ( .A1(C[44]), .A2(n147), .B1(A[44]), .B2(n141), .ZN(n251) );
  AOI222_X1 U111 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n156), .ZN(n250) );
  AOI22_X1 U112 ( .A1(C[48]), .A2(n146), .B1(A[48]), .B2(n140), .ZN(n259) );
  AOI222_X1 U113 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n156), .ZN(n258) );
  NAND2_X1 U114 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI22_X1 U115 ( .A1(C[41]), .A2(n147), .B1(A[41]), .B2(n141), .ZN(n245) );
  AOI222_X1 U116 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n155), .ZN(n244) );
  NAND2_X1 U117 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  AOI222_X1 U118 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n156), .ZN(n270) );
  NAND2_X1 U119 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI222_X1 U120 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n155), .ZN(n230) );
  AOI22_X1 U121 ( .A1(C[35]), .A2(n148), .B1(A[35]), .B2(n142), .ZN(n231) );
  NAND2_X1 U122 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI222_X1 U123 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n155), .ZN(n248) );
  AOI22_X1 U124 ( .A1(C[43]), .A2(n147), .B1(A[43]), .B2(n141), .ZN(n249) );
  NAND2_X1 U125 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  AOI22_X1 U126 ( .A1(C[56]), .A2(n146), .B1(A[56]), .B2(n140), .ZN(n277) );
  AOI222_X1 U127 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n157), .ZN(n276) );
  NAND2_X1 U128 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI22_X1 U129 ( .A1(C[55]), .A2(n146), .B1(A[55]), .B2(n140), .ZN(n275) );
  AOI222_X1 U130 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n156), .ZN(n274) );
  NAND2_X1 U131 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI222_X1 U132 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n156), .ZN(n256) );
  AOI22_X1 U133 ( .A1(C[47]), .A2(n146), .B1(A[47]), .B2(n140), .ZN(n257) );
  NAND2_X1 U134 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  AOI222_X1 U135 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n156), .ZN(n266) );
  AOI22_X1 U136 ( .A1(C[51]), .A2(n146), .B1(A[51]), .B2(n140), .ZN(n267) );
  NAND2_X1 U137 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  AOI22_X1 U138 ( .A1(C[52]), .A2(n146), .B1(A[52]), .B2(n140), .ZN(n269) );
  AOI222_X1 U139 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n156), .ZN(n268) );
  NAND2_X1 U140 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U141 ( .A1(C[60]), .A2(n145), .B1(A[60]), .B2(n139), .ZN(n287) );
  AOI222_X1 U142 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n157), .ZN(n286) );
  NAND2_X1 U143 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U144 ( .A1(C[61]), .A2(n145), .B1(A[61]), .B2(n139), .ZN(n289) );
  AOI222_X1 U145 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n157), .ZN(n288) );
  NAND2_X1 U146 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U147 ( .A1(C[62]), .A2(n145), .B1(A[62]), .B2(n139), .ZN(n291) );
  AOI222_X1 U148 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n157), .ZN(n290) );
  NAND2_X1 U149 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U150 ( .A1(C[63]), .A2(n145), .B1(A[63]), .B2(n139), .ZN(n293) );
  AOI222_X1 U151 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n157), .ZN(n292) );
  NAND2_X1 U152 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U153 ( .A1(C[0]), .A2(n145), .B1(A[0]), .B2(n139), .ZN(n175) );
  AOI222_X1 U154 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n153), .ZN(n174) );
  NAND2_X1 U155 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U156 ( .A1(C[4]), .A2(n146), .B1(A[4]), .B2(n140), .ZN(n263) );
  AOI222_X1 U157 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n156), .ZN(n262) );
  NAND2_X1 U158 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI22_X1 U159 ( .A1(C[8]), .A2(n145), .B1(A[8]), .B2(n139), .ZN(n299) );
  AOI222_X1 U160 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n157), .ZN(n298) );
  NAND2_X1 U161 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  AOI22_X1 U162 ( .A1(C[12]), .A2(n150), .B1(A[12]), .B2(n144), .ZN(n181) );
  AOI222_X1 U163 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n153), .ZN(n180) );
  NAND2_X1 U164 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  AOI22_X1 U165 ( .A1(C[16]), .A2(n149), .B1(A[16]), .B2(n143), .ZN(n189) );
  AOI222_X1 U166 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n153), .ZN(n188) );
  NAND2_X1 U167 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  AOI22_X1 U168 ( .A1(C[20]), .A2(n149), .B1(A[20]), .B2(n143), .ZN(n199) );
  AOI222_X1 U169 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n154), .ZN(n198) );
  NAND2_X1 U170 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U171 ( .A1(C[1]), .A2(n149), .B1(A[1]), .B2(n143), .ZN(n197) );
  AOI222_X1 U172 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n153), .ZN(n196) );
  NAND2_X1 U173 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U174 ( .A1(C[5]), .A2(n145), .B1(A[5]), .B2(n139), .ZN(n285) );
  AOI222_X1 U175 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n157), .ZN(n284) );
  NAND2_X1 U176 ( .A1(n306), .A2(n305), .ZN(Y[9]) );
  AOI22_X1 U177 ( .A1(C[9]), .A2(n147), .B1(A[9]), .B2(n141), .ZN(n306) );
  AOI222_X1 U178 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n157), .ZN(n305) );
  NAND2_X1 U179 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U180 ( .A1(C[13]), .A2(n150), .B1(A[13]), .B2(n144), .ZN(n183) );
  AOI222_X1 U181 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n153), .ZN(n182) );
  NAND2_X1 U182 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI22_X1 U183 ( .A1(C[17]), .A2(n149), .B1(A[17]), .B2(n143), .ZN(n191) );
  AOI222_X1 U184 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n153), .ZN(n190) );
  NAND2_X1 U185 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI22_X1 U186 ( .A1(C[21]), .A2(n149), .B1(A[21]), .B2(n143), .ZN(n201) );
  AOI222_X1 U187 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n154), .ZN(n200) );
  NAND2_X1 U188 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U189 ( .A1(C[2]), .A2(n148), .B1(A[2]), .B2(n142), .ZN(n219) );
  AOI222_X1 U190 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n154), .ZN(n218) );
  NAND2_X1 U191 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U192 ( .A1(C[6]), .A2(n145), .B1(A[6]), .B2(n139), .ZN(n295) );
  AOI222_X1 U193 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n157), .ZN(n294) );
  NAND2_X1 U194 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U195 ( .A1(C[10]), .A2(n150), .B1(A[10]), .B2(n144), .ZN(n177) );
  AOI222_X1 U196 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n153), .ZN(n176) );
  NAND2_X1 U197 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U198 ( .A1(C[14]), .A2(n149), .B1(A[14]), .B2(n143), .ZN(n185) );
  AOI222_X1 U199 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n153), .ZN(n184) );
  NAND2_X1 U200 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI22_X1 U201 ( .A1(C[18]), .A2(n149), .B1(A[18]), .B2(n143), .ZN(n193) );
  AOI222_X1 U202 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n153), .ZN(n192) );
  NAND2_X1 U203 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U204 ( .A1(C[3]), .A2(n147), .B1(A[3]), .B2(n141), .ZN(n241) );
  AOI222_X1 U205 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n155), .ZN(n240) );
  NAND2_X1 U206 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U207 ( .A1(C[7]), .A2(n145), .B1(A[7]), .B2(n139), .ZN(n297) );
  AOI222_X1 U208 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n157), .ZN(n296) );
  NAND2_X1 U209 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U210 ( .A1(C[11]), .A2(n150), .B1(A[11]), .B2(n144), .ZN(n179) );
  AOI222_X1 U211 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n153), .ZN(n178) );
  NAND2_X1 U212 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U213 ( .A1(C[15]), .A2(n149), .B1(A[15]), .B2(n143), .ZN(n187) );
  AOI222_X1 U214 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n153), .ZN(n186) );
  NAND2_X1 U215 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI22_X1 U216 ( .A1(C[19]), .A2(n149), .B1(A[19]), .B2(n143), .ZN(n195) );
  AOI222_X1 U217 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n153), .ZN(n194) );
  AOI22_X1 U218 ( .A1(C[50]), .A2(n146), .B1(A[50]), .B2(n140), .ZN(n265) );
  AOI22_X1 U219 ( .A1(C[49]), .A2(n146), .B1(A[49]), .B2(n140), .ZN(n261) );
  AOI22_X1 U220 ( .A1(C[22]), .A2(n149), .B1(A[22]), .B2(n143), .ZN(n203) );
  AOI22_X1 U221 ( .A1(C[23]), .A2(n149), .B1(A[23]), .B2(n143), .ZN(n205) );
  NAND2_X1 U222 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  NAND2_X1 U223 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI222_X1 U224 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n154), .ZN(n212) );
  AOI222_X1 U225 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n154), .ZN(n210) );
  AOI22_X1 U226 ( .A1(C[45]), .A2(n147), .B1(A[45]), .B2(n141), .ZN(n253) );
  AOI22_X1 U227 ( .A1(C[53]), .A2(n146), .B1(A[53]), .B2(n140), .ZN(n271) );
  AOI222_X1 U228 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n154), .ZN(n208) );
  AOI222_X1 U229 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n154), .ZN(n206) );
  CLKBUF_X1 U230 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U231 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U232 ( .A(n158), .Z(n164) );
endmodule


module G_85 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_315 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_314 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_313 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_312 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_311 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_310 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_309 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_308 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_307 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_306 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_305 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_304 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_303 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_302 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_301 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_300 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_299 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_298 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_297 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_296 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_295 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_294 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_293 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_292 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_291 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_290 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_289 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_288 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_287 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_286 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_285 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_84 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_284 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_283 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_282 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_281 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_280 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_279 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_278 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_277 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_276 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_275 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_274 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_273 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_272 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_271 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3, n5;

  AND2_X1 U1 ( .A1(P_IK), .A2(G_K_1), .ZN(n3) );
  NOR2_X1 U2 ( .A1(n3), .A2(G_IK), .ZN(n5) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U4 ( .A(n5), .ZN(Gx) );
endmodule


module PG_270 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_83 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_269 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_268 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_267 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_266 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  OR2_X2 U2 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U3 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
endmodule


module PG_265 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_264 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  OR2_X1 U2 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_263 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_82 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_81 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_262 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_261 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_260 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3;

  OR2_X1 U1 ( .A1(G_IK), .A2(n3), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n3) );
endmodule


module PG_259 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_258 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_257 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_80 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_79 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_78 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_77 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_256 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_255 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_254 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_253 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_76 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_75 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_74 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_73 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_72 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_71 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_70 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
endmodule


module G_69 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module carry_generator_N64_NPB4_5 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U101 ( .A(B[37]), .B(A[37]), .Z(\PG_Network[0][0][37] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U108 ( .A(B[30]), .B(A[30]), .Z(\PG_Network[0][0][30] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U110 ( .A(B[29]), .B(A[29]), .Z(\PG_Network[0][0][29] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U114 ( .A(B[25]), .B(A[25]), .Z(\PG_Network[0][0][25] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U116 ( .A(B[23]), .B(A[23]), .Z(\PG_Network[0][0][23] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U121 ( .A(B[19]), .B(A[19]), .Z(\PG_Network[0][0][19] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U125 ( .A(B[15]), .B(A[15]), .Z(\PG_Network[0][0][15] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_85 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n29), .Gx(\PG_Network[1][1][1] ) );
  PG_315 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_314 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_313 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_312 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_311 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_310 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_309 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_308 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_307 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_306 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_305 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_304 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_303 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_302 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_301 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_300 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_299 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_298 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_297 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_296 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_295 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_294 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_293 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_292 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_291 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_290 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_289 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_288 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_287 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_286 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_285 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_84 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_284 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_283 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_282 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_281 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_280 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_279 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_278 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_277 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_276 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_275 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_274 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_273 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_272 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_271 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_270 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_83 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_269 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_268 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_267 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_266 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_265 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_264 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_263 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_82 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), 
        .G_K_1(Co[1]), .Gx(Co[3]) );
  G_81 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), 
        .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_262 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_261 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_260 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][47] ), .Px(
        \PG_Network[4][0][47] ) );
  PG_259 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][43] ), .Px(
        \PG_Network[4][0][43] ) );
  PG_258 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(n28), .P_K_1(n19), .Gx(
        \PG_Network[4][1][63] ), .Px(\PG_Network[4][0][63] ) );
  PG_257 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(n28), .P_K_1(n19), .Gx(
        \PG_Network[4][1][59] ), .Px(\PG_Network[4][0][59] ) );
  G_80 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), 
        .G_K_1(Co[3]), .Gx(Co[7]) );
  G_79 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), 
        .G_K_1(Co[3]), .Gx(Co[6]) );
  G_78 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), 
        .G_K_1(Co[3]), .Gx(Co[5]) );
  G_77 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), 
        .G_K_1(Co[3]), .Gx(Co[4]) );
  PG_256 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(n26), .P_K_1(n8), .Gx(
        \PG_Network[5][1][63] ), .Px(\PG_Network[5][0][63] ) );
  PG_255 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(n26), .P_K_1(n8), .Gx(
        \PG_Network[5][1][59] ), .Px(\PG_Network[5][0][59] ) );
  PG_254 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(n26), .P_K_1(n8), .Gx(
        \PG_Network[5][1][55] ), .Px(\PG_Network[5][0][55] ) );
  PG_253 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(n7), 
        .Gx(\PG_Network[5][1][51] ), .Px(\PG_Network[5][0][51] ) );
  G_76 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), 
        .G_K_1(n12), .Gx(Co[15]) );
  G_75 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), 
        .G_K_1(n12), .Gx(Co[14]) );
  G_74 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), 
        .G_K_1(n12), .Gx(Co[13]) );
  G_73 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), 
        .G_K_1(n5), .Gx(Co[12]) );
  G_72 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), 
        .G_K_1(n12), .Gx(Co[11]) );
  G_71 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), 
        .G_K_1(Co[7]), .Gx(Co[10]) );
  G_70 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), 
        .G_K_1(Co[7]), .Gx(Co[9]) );
  G_69 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), 
        .G_K_1(Co[7]), .Gx(Co[8]) );
  INV_X1 U1 ( .A(A[44]), .ZN(n13) );
  CLKBUF_X1 U2 ( .A(Co[7]), .Z(n5) );
  INV_X1 U3 ( .A(A[38]), .ZN(n18) );
  INV_X1 U4 ( .A(A[59]), .ZN(n11) );
  INV_X1 U5 ( .A(A[35]), .ZN(n16) );
  INV_X1 U6 ( .A(A[27]), .ZN(n17) );
  INV_X1 U7 ( .A(A[31]), .ZN(n23) );
  INV_X1 U8 ( .A(A[39]), .ZN(n22) );
  INV_X1 U9 ( .A(A[46]), .ZN(n9) );
  INV_X1 U10 ( .A(A[41]), .ZN(n6) );
  INV_X1 U11 ( .A(A[43]), .ZN(n21) );
  INV_X1 U12 ( .A(A[55]), .ZN(n27) );
  INV_X1 U13 ( .A(A[47]), .ZN(n24) );
  INV_X1 U14 ( .A(A[51]), .ZN(n25) );
  INV_X1 U15 ( .A(A[36]), .ZN(n10) );
  INV_X1 U16 ( .A(A[48]), .ZN(n14) );
  INV_X1 U17 ( .A(A[49]), .ZN(n15) );
  INV_X1 U18 ( .A(A[45]), .ZN(n20) );
  XNOR2_X1 U19 ( .A(B[41]), .B(n6), .ZN(\PG_Network[0][0][41] ) );
  CLKBUF_X1 U20 ( .A(\PG_Network[4][0][47] ), .Z(n7) );
  CLKBUF_X1 U21 ( .A(n7), .Z(n8) );
  XNOR2_X1 U22 ( .A(B[46]), .B(n9), .ZN(\PG_Network[0][0][46] ) );
  XNOR2_X1 U23 ( .A(B[36]), .B(n10), .ZN(\PG_Network[0][0][36] ) );
  XNOR2_X1 U24 ( .A(B[59]), .B(n11), .ZN(\PG_Network[0][0][59] ) );
  CLKBUF_X1 U25 ( .A(Co[7]), .Z(n12) );
  XNOR2_X1 U26 ( .A(B[44]), .B(n13), .ZN(\PG_Network[0][0][44] ) );
  XNOR2_X1 U27 ( .A(B[48]), .B(n14), .ZN(\PG_Network[0][0][48] ) );
  XNOR2_X1 U28 ( .A(B[49]), .B(n15), .ZN(\PG_Network[0][0][49] ) );
  XNOR2_X1 U29 ( .A(B[35]), .B(n16), .ZN(\PG_Network[0][0][35] ) );
  XNOR2_X1 U30 ( .A(B[27]), .B(n17), .ZN(\PG_Network[0][0][27] ) );
  XNOR2_X1 U31 ( .A(B[38]), .B(n18), .ZN(\PG_Network[0][0][38] ) );
  CLKBUF_X1 U32 ( .A(\PG_Network[3][0][55] ), .Z(n19) );
  XNOR2_X1 U33 ( .A(B[45]), .B(n20), .ZN(\PG_Network[0][0][45] ) );
  XNOR2_X1 U34 ( .A(B[43]), .B(n21), .ZN(\PG_Network[0][0][43] ) );
  XNOR2_X1 U35 ( .A(B[39]), .B(n22), .ZN(\PG_Network[0][0][39] ) );
  XNOR2_X1 U36 ( .A(B[31]), .B(n23), .ZN(\PG_Network[0][0][31] ) );
  XNOR2_X1 U37 ( .A(B[47]), .B(n24), .ZN(\PG_Network[0][0][47] ) );
  XNOR2_X1 U38 ( .A(B[51]), .B(n25), .ZN(\PG_Network[0][0][51] ) );
  CLKBUF_X1 U39 ( .A(\PG_Network[4][1][47] ), .Z(n26) );
  XNOR2_X1 U40 ( .A(B[55]), .B(n27), .ZN(\PG_Network[0][0][55] ) );
  CLKBUF_X1 U41 ( .A(\PG_Network[3][1][55] ), .Z(n28) );
  AND2_X1 U42 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U43 ( .A1(B[27]), .A2(A[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U44 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U45 ( .A1(B[31]), .A2(A[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U46 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U47 ( .A1(A[59]), .A2(B[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U48 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U49 ( .A1(B[43]), .A2(A[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U50 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U51 ( .A1(B[46]), .A2(A[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U52 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U53 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U54 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U55 ( .A1(B[41]), .A2(A[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U56 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U57 ( .A1(B[49]), .A2(A[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U58 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U59 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U60 ( .A1(B[45]), .A2(A[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U61 ( .A1(A[25]), .A2(B[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U62 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U63 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U64 ( .A1(A[35]), .A2(B[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U65 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U66 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U67 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U77 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U81 ( .A1(A[37]), .A2(B[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U85 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AND2_X1 U88 ( .A1(A[23]), .A2(B[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U89 ( .A1(B[29]), .A2(A[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U90 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U91 ( .A1(A[53]), .A2(B[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U92 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U93 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U94 ( .A1(A[11]), .A2(B[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U96 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U99 ( .A1(A[15]), .A2(B[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U100 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U102 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U103 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U107 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U112 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U131 ( .A1(A[19]), .A2(B[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U132 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U133 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U134 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U135 ( .A(n32), .ZN(n29) );
  AND2_X1 U136 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U137 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U138 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U139 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U140 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U141 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U142 ( .A1(A[7]), .A2(B[7]), .ZN(\PG_Network[0][1][7] ) );
  AND2_X1 U143 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U144 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AND2_X1 U145 ( .A1(A[21]), .A2(B[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U146 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AOI21_X1 U147 ( .B1(A[0]), .B2(B[0]), .A(n30), .ZN(n32) );
  INV_X1 U148 ( .A(n31), .ZN(n30) );
  OAI21_X1 U149 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n31) );
  AND2_X1 U150 ( .A1(B[55]), .A2(A[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U151 ( .A1(B[51]), .A2(A[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U152 ( .A1(B[47]), .A2(A[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U153 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U154 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
endmodule


module FA_640 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_639 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_638 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_637 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_160 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_640 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_639 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_638 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_637 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_636 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_635 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_634 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_633 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_159 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_636 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_635 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_634 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_633 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_80 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U2 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_80 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_160 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_159 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_80 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_632 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_631 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_630 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_629 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_158 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_632 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_631 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_630 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_629 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_628 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_627 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_626 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_625 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_157 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_628 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_627 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_626 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_625 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_79 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_79 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_158 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_157 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_79 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_624 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_623 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_622 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_621 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_156 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_624 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_623 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_622 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_621 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_620 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_619 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_618 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_617 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_155 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_620 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_619 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_618 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_617 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_78 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_78 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_156 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_155 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_78 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_616 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_615 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_614 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_613 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_154 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_616 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_615 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_614 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_613 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_612 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_611 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_610 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_609 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_153 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_612 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_611 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_610 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_609 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_77 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_77 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_154 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_153 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_77 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_608 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_607 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_606 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_605 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_152 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_608 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_607 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_606 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_605 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_604 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_603 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_602 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_601 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_151 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_604 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_603 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_602 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_601 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_76 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_76 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_152 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_151 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_76 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_600 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_599 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_598 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_597 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_150 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_600 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_599 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_598 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_597 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_596 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_595 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_594 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_593 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_149 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_596 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_595 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_594 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_593 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_75 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_75 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_150 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_149 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_75 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_592 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_591 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_590 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_589 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_148 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_592 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_591 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_590 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_589 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_588 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_587 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_586 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_585 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_147 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_588 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_587 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_586 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_585 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_74 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(sel), .ZN(n13) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n13), .ZN(n17) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_74 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_148 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_147 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_74 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_584 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(n6), .B(B), .ZN(n8) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_583 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_582 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_581 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_146 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_584 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_583 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_582 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_581 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_580 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_579 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_578 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_577 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_145 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_580 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_579 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_578 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_577 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_73 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U4 ( .A(sel), .ZN(n13) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n13), .ZN(n17) );
endmodule


module carry_select_block_NPB4_73 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_146 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_145 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_73 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_576 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_575 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_574 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_573 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_144 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_576 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_575 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_574 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_573 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_572 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_571 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_570 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_569 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_143 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_572 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_571 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_570 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_569 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_72 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U4 ( .A(sel), .ZN(n13) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_72 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_144 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_143 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_72 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_568 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n8), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  AOI22_X1 U6 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_567 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_566 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_565 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_142 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_568 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_567 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_566 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_565 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_564 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_563 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_562 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_561 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_141 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_564 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_563 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_562 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_561 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_71 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19;

  INV_X2 U1 ( .A(n18), .ZN(Y[2]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n5) );
  INV_X1 U3 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U4 ( .A(sel), .ZN(n10) );
  INV_X1 U5 ( .A(sel), .ZN(n11) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[2]), .B1(B[2]), .B2(n11), .ZN(n18) );
  INV_X1 U7 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U8 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n11), .ZN(n17) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n10), .ZN(n16) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n5), .B1(n11), .B2(B[3]), .ZN(n19) );
endmodule


module carry_select_block_NPB4_71 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_142 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_141 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_71 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_560 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7, n8, n9;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n6) );
  CLKBUF_X1 U2 ( .A(n9), .Z(n4) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Co) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n9) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(n7) );
  NAND2_X1 U7 ( .A1(n9), .A2(Ci), .ZN(n8) );
endmodule


module FA_559 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_558 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_557 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  OR2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_140 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_560 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_559 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_558 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_557 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_556 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_555 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_554 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_553 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_139 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_556 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_555 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_554 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_553 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_70 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n16), .ZN(Y[0]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n5) );
  INV_X1 U3 ( .A(sel), .ZN(n10) );
  INV_X1 U4 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n10), .ZN(n16) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n15), .ZN(n17) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n15), .ZN(n19) );
endmodule


module carry_select_block_NPB4_70 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_140 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_139 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_70 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_552 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68176, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  assign Co = net68176;

  INV_X1 U1 ( .A(n6), .ZN(n5) );
  INV_X1 U2 ( .A(Ci), .ZN(n11) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  OR2_X1 U4 ( .A1(B), .A2(n5), .ZN(n8) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(n7), .A2(n8), .ZN(n10) );
  INV_X1 U7 ( .A(A), .ZN(n6) );
  XNOR2_X1 U8 ( .A(n4), .B(A), .ZN(n9) );
  NAND2_X1 U9 ( .A1(A), .A2(n4), .ZN(n12) );
  XNOR2_X1 U10 ( .A(Ci), .B(n9), .ZN(S) );
  OAI21_X1 U11 ( .B1(n10), .B2(n11), .A(n12), .ZN(net68176) );
endmodule


module FA_551 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68175, n4, n5, n6, n7;
  assign Co = net68175;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(n5), .B(B), .ZN(n7) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n7), .ZN(n6) );
  INV_X1 U6 ( .A(n6), .ZN(net68175) );
endmodule


module FA_550 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_549 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(n4), .ZN(n7) );
endmodule


module RCA_N4_138 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_552 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_551 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_550 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_549 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_548 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_547 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(n4), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_546 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_545 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(n4), .ZN(n7) );
endmodule


module RCA_N4_137 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_548 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_547 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_546 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_545 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_69 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X2 U1 ( .A(n16), .ZN(Y[0]) );
  INV_X2 U2 ( .A(n17), .ZN(Y[1]) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n10) );
  INV_X1 U4 ( .A(sel), .ZN(n5) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[2]), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n15), .ZN(n17) );
  INV_X1 U8 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n5), .ZN(n16) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n15), .ZN(n19) );
endmodule


module carry_select_block_NPB4_69 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_138 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_137 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_69 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_544 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68168, n4, n5, n6, n7;
  assign Co = net68168;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  XNOR2_X1 U1 ( .A(B), .B(n7), .ZN(n4) );
  INV_X1 U2 ( .A(A), .ZN(n7) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n5) );
  INV_X1 U5 ( .A(n5), .ZN(net68168) );
  XNOR2_X1 U6 ( .A(B), .B(n7), .ZN(n6) );
endmodule


module FA_543 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68167, net88607, n4, n5, n6;
  assign Co = net68167;

  XOR2_X1 U3 ( .A(Ci), .B(net88607), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n6) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n4) );
  INV_X1 U4 ( .A(n4), .ZN(net68167) );
  XNOR2_X1 U5 ( .A(n6), .B(B), .ZN(n5) );
  CLKBUF_X1 U6 ( .A(n5), .Z(net88607) );
endmodule


module FA_542 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_541 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n8, n10, n11;

  INV_X1 U1 ( .A(n5), .ZN(n4) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n10) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n5), .A2(n10), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n8), .A2(n7), .ZN(S) );
  INV_X1 U6 ( .A(Ci), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(n6) );
  INV_X1 U8 ( .A(n11), .ZN(Co) );
  AOI22_X1 U9 ( .A1(B), .A2(A), .B1(n10), .B2(n4), .ZN(n11) );
endmodule


module RCA_N4_136 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_544 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_543 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_542 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_541 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_540 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_539 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_538 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_537 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_135 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_540 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_539 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_538 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_537 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_68 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n12, n17, n18, n19, n20;

  CLKBUF_X1 U1 ( .A(n10), .Z(n12) );
  CLKBUF_X1 U2 ( .A(n11), .Z(n5) );
  BUF_X1 U3 ( .A(sel), .Z(n11) );
  INV_X1 U4 ( .A(sel), .ZN(n10) );
  INV_X1 U5 ( .A(n17), .ZN(Y[0]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n11), .B1(n12), .B2(B[2]), .ZN(n19) );
  INV_X1 U8 ( .A(n18), .ZN(Y[1]) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[0]), .B1(n10), .B2(B[0]), .ZN(n17) );
  INV_X1 U10 ( .A(n20), .ZN(Y[3]) );
  AOI22_X1 U11 ( .A1(n11), .A2(A[1]), .B1(n10), .B2(B[1]), .ZN(n18) );
  AOI22_X1 U12 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n12), .ZN(n20) );
endmodule


module carry_select_block_NPB4_68 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_136 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_135 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_68 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_536 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68160, n4, n5, n6, n7;
  assign Co = net68160;

  INV_X1 U1 ( .A(Ci), .ZN(n6) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n4) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n7) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n5) );
  XNOR2_X1 U5 ( .A(Ci), .B(n4), .ZN(S) );
  OAI21_X1 U6 ( .B1(n5), .B2(n6), .A(n7), .ZN(net68160) );
endmodule


module FA_535 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n5), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n5) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n7), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_534 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_533 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_134 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_536 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_535 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_534 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_533 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_532 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_531 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_530 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_529 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_133 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_532 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_531 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_530 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_529 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_67 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19, n20;

  CLKBUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(n17), .ZN(Y[0]) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n10) );
  INV_X1 U4 ( .A(n18), .ZN(Y[1]) );
  INV_X1 U5 ( .A(sel), .ZN(n11) );
  INV_X1 U6 ( .A(n19), .ZN(Y[2]) );
  INV_X1 U7 ( .A(n20), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(n5), .A2(A[2]), .B1(n11), .B2(B[2]), .ZN(n19) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[1]), .B1(n16), .B2(B[1]), .ZN(n18) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n16), .B2(B[0]), .ZN(n17) );
  INV_X1 U11 ( .A(sel), .ZN(n16) );
  AOI22_X1 U12 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n11), .ZN(n20) );
endmodule


module carry_select_block_NPB4_67 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_134 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_133 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_67 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_528 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_527 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_526 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_525 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_132 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_528 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_527 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_526 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_525 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_524 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_523 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_522 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_521 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_131 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_524 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_523 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_522 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_521 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_66 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n10), .ZN(n5) );
  INV_X1 U2 ( .A(n16), .ZN(Y[0]) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n10) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(n10), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U11 ( .A(sel), .ZN(n15) );
endmodule


module carry_select_block_NPB4_66 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_132 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_131 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_66 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_520 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_519 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_518 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_517 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_130 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_520 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_519 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_518 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_517 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_516 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_515 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_514 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_513 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_129 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_516 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_515 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_514 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_513 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_65 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n15), .ZN(Y[0]) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n5) );
  INV_X1 U3 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U4 ( .A(sel), .ZN(n14) );
  INV_X1 U5 ( .A(n17), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n14), .ZN(n17) );
  INV_X1 U7 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U9 ( .A1(n5), .A2(A[3]), .B1(B[3]), .B2(n14), .ZN(n18) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n14), .ZN(n15) );
endmodule


module carry_select_block_NPB4_65 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_130 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_129 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_65 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_5 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_80 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_79 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_78 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_77 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_76 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_75 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_74 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_73 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_72 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_71 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_70 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), 
        .S(S[43:40]) );
  carry_select_block_NPB4_69 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), 
        .S(S[47:44]) );
  carry_select_block_NPB4_68 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), 
        .S(S[51:48]) );
  carry_select_block_NPB4_67 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), 
        .S(S[55:52]) );
  carry_select_block_NPB4_66 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), 
        .S(S[59:56]) );
  carry_select_block_NPB4_65 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), 
        .S(S[63:60]) );
endmodule


module P4_ADDER_N64_5 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_5 CGEN ( .A(A), .B({B[63:57], n6, B[55:54], n8, n10, 
        B[51:49], n15, B[47:37], n19, B[35:25], n1, B[23:0]}), .Cin(Cin), .Co(
        CoutCgen) );
  sum_generator_N64_NPB4_5 SGEN ( .A(A), .B({B[63:56], n14, B[54:52], n5, 
        B[50:48], n11, n9, n16, B[44], n13, n7, B[41:40], n2, B[38:36], n12, 
        B[34:32], n3, B[30:28], n18, B[26:0]}), .Ci({CoutCgen, Cin}), .S(S), 
        .Co(Cout) );
  BUF_X1 U1 ( .A(B[45]), .Z(n16) );
  CLKBUF_X1 U2 ( .A(B[24]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(B[39]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(B[31]), .Z(n3) );
  BUF_X1 U5 ( .A(B[36]), .Z(n19) );
  INV_X1 U6 ( .A(B[51]), .ZN(n4) );
  INV_X1 U7 ( .A(n4), .ZN(n5) );
  BUF_X1 U8 ( .A(B[55]), .Z(n14) );
  BUF_X1 U9 ( .A(B[53]), .Z(n8) );
  CLKBUF_X1 U10 ( .A(B[56]), .Z(n6) );
  CLKBUF_X1 U11 ( .A(B[42]), .Z(n7) );
  CLKBUF_X1 U12 ( .A(B[46]), .Z(n9) );
  CLKBUF_X1 U13 ( .A(B[52]), .Z(n10) );
  CLKBUF_X1 U14 ( .A(B[47]), .Z(n11) );
  CLKBUF_X1 U15 ( .A(B[35]), .Z(n12) );
  CLKBUF_X1 U16 ( .A(B[43]), .Z(n13) );
  CLKBUF_X1 U17 ( .A(B[48]), .Z(n15) );
  INV_X1 U18 ( .A(B[27]), .ZN(n17) );
  INV_X1 U19 ( .A(n17), .ZN(n18) );
endmodule


module Booth_Encoder_4 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_4 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306;

  NAND2_X1 U1 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  NAND2_X1 U2 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  NAND2_X1 U3 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  NAND2_X1 U4 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  NOR3_X1 U5 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U6 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  AOI222_X1 U7 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n155), .ZN(n230) );
  BUF_X1 U8 ( .A(n158), .Z(n161) );
  BUF_X1 U9 ( .A(n158), .Z(n160) );
  BUF_X1 U10 ( .A(n158), .Z(n163) );
  BUF_X1 U11 ( .A(n158), .Z(n162) );
  BUF_X1 U12 ( .A(n158), .Z(n159) );
  BUF_X1 U13 ( .A(n151), .Z(n153) );
  BUF_X1 U14 ( .A(n165), .Z(n167) );
  BUF_X1 U15 ( .A(n303), .Z(n158) );
  NOR4_X1 U16 ( .A1(n150), .A2(n144), .A3(n153), .A4(n167), .ZN(n303) );
  BUF_X1 U17 ( .A(n151), .Z(n155) );
  BUF_X1 U18 ( .A(n165), .Z(n169) );
  BUF_X1 U19 ( .A(n151), .Z(n154) );
  BUF_X1 U20 ( .A(n165), .Z(n168) );
  BUF_X1 U21 ( .A(n152), .Z(n156) );
  BUF_X1 U22 ( .A(n166), .Z(n170) );
  BUF_X1 U23 ( .A(n152), .Z(n157) );
  BUF_X1 U24 ( .A(n166), .Z(n171) );
  BUF_X1 U25 ( .A(n304), .Z(n165) );
  BUF_X1 U26 ( .A(n302), .Z(n151) );
  BUF_X1 U27 ( .A(n301), .Z(n147) );
  BUF_X1 U28 ( .A(n301), .Z(n149) );
  BUF_X1 U29 ( .A(n301), .Z(n148) );
  BUF_X1 U30 ( .A(n301), .Z(n146) );
  BUF_X1 U31 ( .A(n304), .Z(n166) );
  BUF_X1 U32 ( .A(n302), .Z(n152) );
  BUF_X1 U33 ( .A(n301), .Z(n145) );
  BUF_X1 U34 ( .A(n300), .Z(n141) );
  BUF_X1 U35 ( .A(n300), .Z(n139) );
  BUF_X1 U36 ( .A(n300), .Z(n143) );
  BUF_X1 U37 ( .A(n300), .Z(n142) );
  BUF_X1 U38 ( .A(n300), .Z(n140) );
  INV_X1 U39 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U40 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n304) );
  AND3_X1 U41 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U42 ( .A(sel[2]), .ZN(n173) );
  AOI22_X1 U43 ( .A1(C[44]), .A2(n147), .B1(A[44]), .B2(n141), .ZN(n251) );
  AOI222_X1 U44 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n156), .ZN(n250) );
  NAND2_X1 U45 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI22_X1 U46 ( .A1(C[50]), .A2(n146), .B1(A[50]), .B2(n140), .ZN(n265) );
  AOI222_X1 U47 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n156), .ZN(n264) );
  AOI222_X1 U48 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n154), .ZN(n208) );
  NAND2_X1 U49 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI22_X1 U50 ( .A1(C[26]), .A2(n148), .B1(A[26]), .B2(n142), .ZN(n211) );
  NAND2_X1 U51 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI22_X1 U52 ( .A1(C[29]), .A2(n148), .B1(A[29]), .B2(n142), .ZN(n217) );
  NAND2_X1 U53 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI22_X1 U54 ( .A1(C[27]), .A2(n148), .B1(A[27]), .B2(n142), .ZN(n213) );
  NAND2_X1 U55 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U56 ( .A1(C[30]), .A2(n148), .B1(A[30]), .B2(n142), .ZN(n221) );
  AOI222_X1 U57 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n154), .ZN(n220) );
  NAND2_X1 U58 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI22_X1 U59 ( .A1(C[31]), .A2(n148), .B1(A[31]), .B2(n142), .ZN(n223) );
  AOI222_X1 U60 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n154), .ZN(n222) );
  NAND2_X1 U61 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI222_X1 U62 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n155), .ZN(n248) );
  AOI22_X1 U63 ( .A1(C[43]), .A2(n147), .B1(A[43]), .B2(n141), .ZN(n249) );
  AOI22_X1 U64 ( .A1(C[48]), .A2(n146), .B1(A[48]), .B2(n140), .ZN(n259) );
  NAND2_X1 U65 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  AOI22_X1 U66 ( .A1(C[28]), .A2(n148), .B1(A[28]), .B2(n142), .ZN(n215) );
  NAND2_X1 U67 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI22_X1 U68 ( .A1(C[46]), .A2(n146), .B1(A[46]), .B2(n140), .ZN(n255) );
  AOI222_X1 U69 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n156), .ZN(n254) );
  NAND2_X1 U70 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI22_X1 U71 ( .A1(C[54]), .A2(n146), .B1(A[54]), .B2(n140), .ZN(n273) );
  AOI222_X1 U72 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n156), .ZN(n272) );
  NAND2_X1 U73 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  AOI22_X1 U74 ( .A1(C[57]), .A2(n145), .B1(A[57]), .B2(n139), .ZN(n279) );
  AOI222_X1 U75 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n157), .ZN(n278) );
  NAND2_X1 U76 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI222_X1 U77 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n156), .ZN(n260) );
  AOI22_X1 U78 ( .A1(C[49]), .A2(n146), .B1(A[49]), .B2(n140), .ZN(n261) );
  NAND2_X1 U79 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  AOI22_X1 U80 ( .A1(C[53]), .A2(n146), .B1(A[53]), .B2(n140), .ZN(n271) );
  AOI222_X1 U81 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n156), .ZN(n270) );
  NAND2_X1 U82 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI222_X1 U83 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n156), .ZN(n252) );
  AOI22_X1 U84 ( .A1(C[45]), .A2(n147), .B1(A[45]), .B2(n141), .ZN(n253) );
  NAND2_X1 U85 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  NAND2_X1 U86 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  NAND2_X1 U87 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  NAND2_X1 U88 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  NAND2_X1 U89 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  AOI222_X1 U90 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n157), .ZN(n276) );
  AOI22_X1 U91 ( .A1(C[56]), .A2(n146), .B1(A[56]), .B2(n140), .ZN(n277) );
  AOI222_X1 U92 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n154), .ZN(n206) );
  AOI22_X1 U93 ( .A1(C[40]), .A2(n147), .B1(A[40]), .B2(n141), .ZN(n243) );
  AOI222_X1 U94 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n155), .ZN(n242) );
  NAND2_X1 U95 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  AOI22_X1 U96 ( .A1(C[32]), .A2(n148), .B1(A[32]), .B2(n142), .ZN(n225) );
  AOI222_X1 U97 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n155), .ZN(n224) );
  NAND2_X1 U98 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI22_X1 U99 ( .A1(C[34]), .A2(n148), .B1(A[34]), .B2(n142), .ZN(n229) );
  AOI222_X1 U100 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n155), .ZN(n228) );
  NAND2_X1 U101 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI222_X1 U102 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n155), .ZN(n236) );
  AOI22_X1 U103 ( .A1(C[38]), .A2(n147), .B1(A[38]), .B2(n141), .ZN(n237) );
  NAND2_X1 U104 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U105 ( .A1(C[61]), .A2(n145), .B1(A[61]), .B2(n139), .ZN(n289) );
  AOI222_X1 U106 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n157), .ZN(n288) );
  NAND2_X1 U107 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI22_X1 U108 ( .A1(C[58]), .A2(n145), .B1(A[58]), .B2(n139), .ZN(n281) );
  AOI222_X1 U109 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n157), .ZN(n280) );
  NAND2_X1 U110 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U111 ( .A1(C[59]), .A2(n145), .B1(A[59]), .B2(n139), .ZN(n283) );
  AOI222_X1 U112 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n157), .ZN(n282) );
  NAND2_X1 U113 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI22_X1 U114 ( .A1(C[35]), .A2(n148), .B1(A[35]), .B2(n142), .ZN(n231) );
  NAND2_X1 U115 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI22_X1 U116 ( .A1(C[33]), .A2(n148), .B1(A[33]), .B2(n142), .ZN(n227) );
  AOI222_X1 U117 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n155), .ZN(n226) );
  NAND2_X1 U118 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI222_X1 U119 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n155), .ZN(n234) );
  AOI22_X1 U120 ( .A1(C[37]), .A2(n147), .B1(A[37]), .B2(n141), .ZN(n235) );
  NAND2_X1 U121 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U122 ( .A1(C[63]), .A2(n145), .B1(A[63]), .B2(n139), .ZN(n293) );
  AOI222_X1 U123 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n157), .ZN(n292) );
  AOI22_X1 U124 ( .A1(C[36]), .A2(n147), .B1(A[36]), .B2(n141), .ZN(n233) );
  AOI222_X1 U125 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n155), .ZN(n232) );
  NAND2_X1 U126 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI222_X1 U127 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n155), .ZN(n246) );
  AOI22_X1 U128 ( .A1(C[42]), .A2(n147), .B1(A[42]), .B2(n141), .ZN(n247) );
  NAND2_X1 U129 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U130 ( .A1(C[60]), .A2(n145), .B1(A[60]), .B2(n139), .ZN(n287) );
  AOI222_X1 U131 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n157), .ZN(n286) );
  NAND2_X1 U132 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI222_X1 U133 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n155), .ZN(n244) );
  AOI22_X1 U134 ( .A1(C[41]), .A2(n147), .B1(A[41]), .B2(n141), .ZN(n245) );
  NAND2_X1 U135 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U136 ( .A1(C[62]), .A2(n145), .B1(A[62]), .B2(n139), .ZN(n291) );
  AOI222_X1 U137 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n157), .ZN(n290) );
  NAND2_X1 U138 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI222_X1 U139 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n155), .ZN(n238) );
  AOI22_X1 U140 ( .A1(C[39]), .A2(n147), .B1(A[39]), .B2(n141), .ZN(n239) );
  NAND2_X1 U141 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U142 ( .A1(C[0]), .A2(n145), .B1(A[0]), .B2(n139), .ZN(n175) );
  AOI222_X1 U143 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n153), .ZN(n174) );
  NAND2_X1 U144 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U145 ( .A1(C[4]), .A2(n146), .B1(A[4]), .B2(n140), .ZN(n263) );
  AOI222_X1 U146 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n156), .ZN(n262) );
  NAND2_X1 U147 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI22_X1 U148 ( .A1(C[8]), .A2(n145), .B1(A[8]), .B2(n139), .ZN(n299) );
  AOI222_X1 U149 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n157), .ZN(n298) );
  NAND2_X1 U150 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  AOI22_X1 U151 ( .A1(C[12]), .A2(n150), .B1(A[12]), .B2(n144), .ZN(n181) );
  AOI222_X1 U152 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n153), .ZN(n180) );
  NAND2_X1 U153 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  AOI22_X1 U154 ( .A1(C[16]), .A2(n149), .B1(A[16]), .B2(n143), .ZN(n189) );
  AOI222_X1 U155 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n153), .ZN(n188) );
  NAND2_X1 U156 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  AOI22_X1 U157 ( .A1(C[20]), .A2(n149), .B1(A[20]), .B2(n143), .ZN(n199) );
  AOI222_X1 U158 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n154), .ZN(n198) );
  NAND2_X1 U159 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U160 ( .A1(C[1]), .A2(n149), .B1(A[1]), .B2(n143), .ZN(n197) );
  AOI222_X1 U161 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n153), .ZN(n196) );
  NAND2_X1 U162 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U163 ( .A1(C[5]), .A2(n145), .B1(A[5]), .B2(n139), .ZN(n285) );
  AOI222_X1 U164 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n157), .ZN(n284) );
  NAND2_X1 U165 ( .A1(n306), .A2(n305), .ZN(Y[9]) );
  AOI22_X1 U166 ( .A1(C[9]), .A2(n147), .B1(A[9]), .B2(n141), .ZN(n306) );
  AOI222_X1 U167 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n157), .ZN(n305) );
  NAND2_X1 U168 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U169 ( .A1(C[13]), .A2(n150), .B1(A[13]), .B2(n144), .ZN(n183) );
  AOI222_X1 U170 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n153), .ZN(n182) );
  NAND2_X1 U171 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI22_X1 U172 ( .A1(C[17]), .A2(n149), .B1(A[17]), .B2(n143), .ZN(n191) );
  AOI222_X1 U173 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n153), .ZN(n190) );
  NAND2_X1 U174 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI22_X1 U175 ( .A1(C[21]), .A2(n149), .B1(A[21]), .B2(n143), .ZN(n201) );
  AOI222_X1 U176 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n154), .ZN(n200) );
  NAND2_X1 U177 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U178 ( .A1(C[2]), .A2(n148), .B1(A[2]), .B2(n142), .ZN(n219) );
  AOI222_X1 U179 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n154), .ZN(n218) );
  NAND2_X1 U180 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U181 ( .A1(C[6]), .A2(n145), .B1(A[6]), .B2(n139), .ZN(n295) );
  AOI222_X1 U182 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n157), .ZN(n294) );
  NAND2_X1 U183 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U184 ( .A1(C[10]), .A2(n150), .B1(A[10]), .B2(n144), .ZN(n177) );
  AOI222_X1 U185 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n153), .ZN(n176) );
  NAND2_X1 U186 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U187 ( .A1(C[14]), .A2(n149), .B1(A[14]), .B2(n143), .ZN(n185) );
  AOI222_X1 U188 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n153), .ZN(n184) );
  NAND2_X1 U189 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI22_X1 U190 ( .A1(C[18]), .A2(n149), .B1(A[18]), .B2(n143), .ZN(n193) );
  AOI222_X1 U191 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n153), .ZN(n192) );
  NAND2_X1 U192 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI22_X1 U193 ( .A1(C[22]), .A2(n149), .B1(A[22]), .B2(n143), .ZN(n203) );
  AOI222_X1 U194 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n154), .ZN(n202) );
  NAND2_X1 U195 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U196 ( .A1(C[3]), .A2(n147), .B1(A[3]), .B2(n141), .ZN(n241) );
  AOI222_X1 U197 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n155), .ZN(n240) );
  NAND2_X1 U198 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U199 ( .A1(C[7]), .A2(n145), .B1(A[7]), .B2(n139), .ZN(n297) );
  AOI222_X1 U200 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n157), .ZN(n296) );
  NAND2_X1 U201 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U202 ( .A1(C[11]), .A2(n150), .B1(A[11]), .B2(n144), .ZN(n179) );
  AOI222_X1 U203 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n153), .ZN(n178) );
  NAND2_X1 U204 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U205 ( .A1(C[15]), .A2(n149), .B1(A[15]), .B2(n143), .ZN(n187) );
  AOI222_X1 U206 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n153), .ZN(n186) );
  NAND2_X1 U207 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI22_X1 U208 ( .A1(C[19]), .A2(n149), .B1(A[19]), .B2(n143), .ZN(n195) );
  AOI222_X1 U209 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n153), .ZN(n194) );
  NAND2_X1 U210 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI22_X1 U211 ( .A1(C[23]), .A2(n149), .B1(A[23]), .B2(n143), .ZN(n205) );
  AOI222_X1 U212 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n154), .ZN(n204) );
  AOI22_X1 U213 ( .A1(C[52]), .A2(n146), .B1(A[52]), .B2(n140), .ZN(n269) );
  AOI22_X1 U214 ( .A1(C[51]), .A2(n146), .B1(A[51]), .B2(n140), .ZN(n267) );
  AOI222_X1 U215 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n156), .ZN(n266) );
  AOI22_X1 U216 ( .A1(C[24]), .A2(n149), .B1(A[24]), .B2(n143), .ZN(n207) );
  AOI22_X1 U217 ( .A1(C[25]), .A2(n148), .B1(A[25]), .B2(n142), .ZN(n209) );
  NAND2_X1 U218 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  NAND2_X1 U219 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI222_X1 U220 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n154), .ZN(n216) );
  AOI222_X1 U221 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n154), .ZN(n214) );
  AOI22_X1 U222 ( .A1(C[47]), .A2(n146), .B1(A[47]), .B2(n140), .ZN(n257) );
  AOI222_X1 U223 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n156), .ZN(n268) );
  AOI222_X1 U224 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n156), .ZN(n256) );
  AOI222_X1 U225 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n156), .ZN(n258) );
  AOI22_X1 U226 ( .A1(C[55]), .A2(n146), .B1(A[55]), .B2(n140), .ZN(n275) );
  AOI222_X1 U227 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n156), .ZN(n274) );
  AOI222_X1 U228 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n154), .ZN(n210) );
  AOI222_X1 U229 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n154), .ZN(n212) );
  CLKBUF_X1 U230 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U231 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U232 ( .A(n158), .Z(n164) );
endmodule


module G_68 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_252 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_251 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_250 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_249 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_248 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_247 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_246 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_245 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_244 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_243 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_242 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_241 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_240 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3, n5;

  CLKBUF_X1 U1 ( .A(P_IK), .Z(n3) );
  INV_X1 U2 ( .A(n5), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n5) );
  AND2_X1 U4 ( .A1(n3), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_239 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_238 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_237 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_236 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_235 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3, n5;

  CLKBUF_X1 U1 ( .A(P_IK), .Z(n3) );
  INV_X1 U2 ( .A(n5), .ZN(Gx) );
  AND2_X1 U3 ( .A1(n3), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U4 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n5) );
endmodule


module PG_234 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_233 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_232 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_231 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_230 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_229 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_228 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_227 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_226 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_225 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_224 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_223 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_222 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_67 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_221 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_220 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_219 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_218 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_217 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_216 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_215 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_214 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_213 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3, n5;

  AND2_X1 U1 ( .A1(P_IK), .A2(G_K_1), .ZN(n3) );
  NOR2_X1 U2 ( .A1(n3), .A2(G_IK), .ZN(n5) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U4 ( .A(n5), .ZN(Gx) );
endmodule


module PG_212 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_211 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_210 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_209 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_208 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_207 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_66 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_206 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_205 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_204 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_203 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_202 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_201 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AND2_X1 U3 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
endmodule


module PG_200 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_65 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_64 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_199 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_198 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_197 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n3) );
  OR2_X2 U3 ( .A1(G_IK), .A2(n3), .ZN(Gx) );
endmodule


module PG_196 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_195 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_194 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_63 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_62 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_61 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_60 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_193 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_192 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_191 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_190 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module G_59 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_58 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_57 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_56 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_55 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_54 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_53 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_52 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module carry_generator_N64_NPB4_4 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   n29, \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n11, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U91 ( .A(B[46]), .B(A[46]), .Z(\PG_Network[0][0][46] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U100 ( .A(B[38]), .B(A[38]), .Z(\PG_Network[0][0][38] ) );
  XOR2_X1 U101 ( .A(B[37]), .B(A[37]), .Z(\PG_Network[0][0][37] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U108 ( .A(B[30]), .B(A[30]), .Z(\PG_Network[0][0][30] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U110 ( .A(B[29]), .B(A[29]), .Z(\PG_Network[0][0][29] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U114 ( .A(B[25]), .B(A[25]), .Z(\PG_Network[0][0][25] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U116 ( .A(B[23]), .B(A[23]), .Z(\PG_Network[0][0][23] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U121 ( .A(B[19]), .B(A[19]), .Z(\PG_Network[0][0][19] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U125 ( .A(B[15]), .B(A[15]), .Z(\PG_Network[0][0][15] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_68 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n25), .Gx(\PG_Network[1][1][1] ) );
  PG_252 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_251 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_250 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_249 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_248 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_247 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_246 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_245 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_244 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_243 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_242 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_241 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_240 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_239 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_238 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_237 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_236 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_235 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_234 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_233 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_232 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_231 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_230 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_229 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_228 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_227 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_226 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_225 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_224 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_223 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_222 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_67 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_221 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_220 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_219 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_218 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_217 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_216 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_215 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_214 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_213 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_212 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_211 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_210 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_209 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_208 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_207 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_66 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_206 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_205 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_204 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_203 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_202 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_201 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_200 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(n5), .P_K_1(\PG_Network[2][0][59] ), 
        .Gx(\PG_Network[3][1][63] ), .Px(\PG_Network[3][0][63] ) );
  G_65 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), 
        .G_K_1(Co[1]), .Gx(Co[3]) );
  G_64 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), 
        .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_199 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_198 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_197 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][47] ), .Px(
        \PG_Network[4][0][47] ) );
  PG_196 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][43] ), .Px(
        \PG_Network[4][0][43] ) );
  PG_195 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(n16), .P_K_1(n18), .Gx(
        \PG_Network[4][1][63] ), .Px(\PG_Network[4][0][63] ) );
  PG_194 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(n16), .P_K_1(n18), .Gx(
        \PG_Network[4][1][59] ), .Px(\PG_Network[4][0][59] ) );
  G_63 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), 
        .G_K_1(Co[3]), .Gx(n29) );
  G_62 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), 
        .G_K_1(Co[3]), .Gx(Co[6]) );
  G_61 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), 
        .G_K_1(Co[3]), .Gx(Co[5]) );
  G_60 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), 
        .G_K_1(Co[3]), .Gx(Co[4]) );
  PG_193 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(n19), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][63] ), .Px(\PG_Network[5][0][63] ) );
  PG_192 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(n19), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][59] ), .Px(\PG_Network[5][0][59] ) );
  PG_191 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(n11), .P_K_1(\PG_Network[4][0][47] ), 
        .Gx(\PG_Network[5][1][55] ), .Px(\PG_Network[5][0][55] ) );
  PG_190 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][51] ), .Px(
        \PG_Network[5][0][51] ) );
  G_59 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), 
        .G_K_1(n20), .Gx(Co[15]) );
  G_58 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), 
        .G_K_1(n20), .Gx(Co[14]) );
  G_57 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), 
        .G_K_1(n20), .Gx(Co[13]) );
  G_56 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), 
        .G_K_1(n20), .Gx(Co[12]) );
  G_55 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), 
        .G_K_1(n20), .Gx(Co[11]) );
  G_54 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), 
        .G_K_1(n10), .Gx(Co[10]) );
  G_53 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), 
        .G_K_1(n29), .Gx(Co[9]) );
  G_52 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), 
        .G_K_1(n29), .Gx(Co[8]) );
  CLKBUF_X1 U1 ( .A(\PG_Network[2][1][59] ), .Z(n5) );
  INV_X1 U2 ( .A(A[27]), .ZN(n12) );
  INV_X1 U3 ( .A(A[31]), .ZN(n14) );
  INV_X1 U4 ( .A(A[59]), .ZN(n15) );
  INV_X1 U5 ( .A(A[35]), .ZN(n7) );
  INV_X1 U6 ( .A(A[43]), .ZN(n8) );
  INV_X1 U7 ( .A(A[54]), .ZN(n6) );
  INV_X1 U8 ( .A(A[45]), .ZN(n21) );
  INV_X1 U9 ( .A(A[55]), .ZN(n24) );
  INV_X1 U10 ( .A(A[47]), .ZN(n23) );
  INV_X1 U11 ( .A(A[51]), .ZN(n22) );
  INV_X1 U12 ( .A(A[39]), .ZN(n17) );
  INV_X1 U13 ( .A(A[49]), .ZN(n9) );
  XNOR2_X1 U14 ( .A(B[54]), .B(n6), .ZN(\PG_Network[0][0][54] ) );
  XNOR2_X1 U15 ( .A(B[35]), .B(n7), .ZN(\PG_Network[0][0][35] ) );
  CLKBUF_X1 U16 ( .A(\PG_Network[4][1][47] ), .Z(n11) );
  XNOR2_X1 U17 ( .A(B[43]), .B(n8), .ZN(\PG_Network[0][0][43] ) );
  XNOR2_X1 U18 ( .A(B[49]), .B(n9), .ZN(\PG_Network[0][0][49] ) );
  CLKBUF_X1 U19 ( .A(n29), .Z(n10) );
  XNOR2_X1 U20 ( .A(B[27]), .B(n12), .ZN(\PG_Network[0][0][27] ) );
  BUF_X2 U21 ( .A(n29), .Z(Co[7]) );
  XNOR2_X1 U22 ( .A(B[31]), .B(n14), .ZN(\PG_Network[0][0][31] ) );
  XNOR2_X1 U23 ( .A(B[59]), .B(n15), .ZN(\PG_Network[0][0][59] ) );
  CLKBUF_X1 U24 ( .A(\PG_Network[3][1][55] ), .Z(n16) );
  XNOR2_X1 U25 ( .A(B[39]), .B(n17), .ZN(\PG_Network[0][0][39] ) );
  CLKBUF_X1 U26 ( .A(\PG_Network[3][0][55] ), .Z(n18) );
  CLKBUF_X1 U27 ( .A(n11), .Z(n19) );
  CLKBUF_X1 U28 ( .A(n10), .Z(n20) );
  XNOR2_X1 U29 ( .A(B[45]), .B(n21), .ZN(\PG_Network[0][0][45] ) );
  XNOR2_X1 U30 ( .A(B[51]), .B(n22), .ZN(\PG_Network[0][0][51] ) );
  XNOR2_X1 U31 ( .A(B[47]), .B(n23), .ZN(\PG_Network[0][0][47] ) );
  XNOR2_X1 U32 ( .A(B[55]), .B(n24), .ZN(\PG_Network[0][0][55] ) );
  AND2_X1 U33 ( .A1(A[46]), .A2(B[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U34 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U35 ( .A1(B[45]), .A2(A[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U36 ( .A1(B[54]), .A2(A[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U37 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U38 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U39 ( .A1(A[37]), .A2(B[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U40 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U41 ( .A1(B[41]), .A2(A[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U42 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U43 ( .A1(B[43]), .A2(A[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U44 ( .A1(B[49]), .A2(A[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U45 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U46 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U47 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U48 ( .A1(A[27]), .A2(B[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U49 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U50 ( .A1(A[25]), .A2(B[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U51 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U52 ( .A1(A[35]), .A2(B[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U53 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U54 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U55 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U56 ( .A1(A[29]), .A2(B[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U57 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U58 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U59 ( .A1(A[59]), .A2(B[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U60 ( .A1(B[53]), .A2(A[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U61 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U62 ( .A1(B[31]), .A2(A[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U63 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U64 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U65 ( .A1(A[11]), .A2(B[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U66 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U67 ( .A1(A[15]), .A2(B[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U77 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U81 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U82 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U85 ( .A1(A[19]), .A2(B[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U88 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U90 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U92 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U94 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U99 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U103 ( .A(n28), .ZN(n25) );
  AND2_X1 U107 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U112 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U131 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U132 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U133 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U134 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U135 ( .A1(A[7]), .A2(B[7]), .ZN(\PG_Network[0][1][7] ) );
  AND2_X1 U136 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U137 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AND2_X1 U138 ( .A1(A[21]), .A2(B[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U139 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U140 ( .A1(A[23]), .A2(B[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U141 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AOI21_X1 U142 ( .B1(A[0]), .B2(B[0]), .A(n26), .ZN(n28) );
  INV_X1 U143 ( .A(n27), .ZN(n26) );
  OAI21_X1 U144 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n27) );
  AND2_X1 U145 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U146 ( .A1(B[51]), .A2(A[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U147 ( .A1(B[47]), .A2(A[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U148 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U149 ( .A1(B[55]), .A2(A[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U150 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
endmodule


module FA_512 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_511 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_510 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_509 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_128 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_512 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_511 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_510 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_509 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_508 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_507 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_506 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_505 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_127 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_508 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_507 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_506 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_505 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_64 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U2 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U4 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U7 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_64 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_128 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_127 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_64 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_504 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_503 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_502 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_501 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_126 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_504 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_503 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_502 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_501 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_500 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_499 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_498 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_497 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_125 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_500 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_499 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_498 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_497 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_63 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_63 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_126 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_125 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_63 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_496 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_495 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_494 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_493 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_124 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_496 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_495 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_494 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_493 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_492 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_491 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_490 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_489 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_123 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_492 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_491 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_490 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_489 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_62 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_62 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_124 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_123 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_62 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_488 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_487 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_486 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_485 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_122 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_488 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_487 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_486 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_485 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_484 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_483 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_482 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_481 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_121 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_484 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_483 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_482 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_481 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_61 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_61 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_122 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_121 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_61 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_480 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_479 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_478 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_477 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_120 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_480 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_479 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_478 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_477 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_476 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_475 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_474 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_473 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_119 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_476 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_475 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_474 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_473 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_60 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_60 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_120 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_119 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_60 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_472 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_471 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_470 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_469 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_118 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_472 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_471 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_470 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_469 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_468 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_467 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_466 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_465 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_117 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_468 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_467 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_466 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_465 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_59 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_59 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_118 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_117 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_59 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_464 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_463 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_462 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_461 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_116 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_464 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_463 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_462 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_461 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_460 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_459 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_458 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_457 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_115 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_460 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_459 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_458 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_457 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_58 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U2 ( .A(sel), .ZN(n13) );
  INV_X1 U3 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U4 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_58 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_116 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_115 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_58 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_456 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_455 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_454 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_453 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_114 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_456 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_455 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_454 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_453 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_452 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_451 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_450 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_449 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_113 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_452 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_451 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_450 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_449 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_57 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X2 U1 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n17), .ZN(Y[2]) );
  CLKBUF_X1 U4 ( .A(sel), .Z(n5) );
  INV_X1 U5 ( .A(sel), .ZN(n14) );
  INV_X1 U6 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n14), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n14), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n14), .ZN(n15) );
endmodule


module carry_select_block_NPB4_57 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_114 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_113 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_57 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_448 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n5), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_447 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_446 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_445 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_112 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_448 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_447 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_446 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_445 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_444 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_443 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_442 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_441 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_111 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_444 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_443 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_442 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_441 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_56 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U3 ( .A(sel), .ZN(n5) );
  INV_X2 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n17) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n16) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n5), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n5), .ZN(n14) );
endmodule


module carry_select_block_NPB4_56 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_112 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_111 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_56 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_440 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_439 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_438 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_437 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_110 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_440 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_439 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_438 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_437 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_436 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_435 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_434 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_433 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_109 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_436 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_435 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_434 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_433 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_55 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n18), .ZN(Y[2]) );
  CLKBUF_X1 U4 ( .A(sel), .Z(n5) );
  INV_X1 U5 ( .A(sel), .ZN(n10) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n10), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n15), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
  INV_X1 U10 ( .A(sel), .ZN(n15) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n10), .ZN(n19) );
endmodule


module carry_select_block_NPB4_55 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_110 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_109 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_55 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_432 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(n5), .B(B), .ZN(n7) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_431 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_430 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_429 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_108 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_432 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_431 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_430 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_429 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_428 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_427 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_426 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_425 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_107 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_428 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_427 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_426 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_425 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_54 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17;

  INV_X2 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U3 ( .A(sel), .ZN(n5) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n16) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n5), .ZN(n17) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n5), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n5), .ZN(n14) );
endmodule


module carry_select_block_NPB4_54 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_108 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_107 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_54 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_424 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  XNOR2_X1 U1 ( .A(B), .B(n5), .ZN(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_423 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68047, n4, n5;
  assign Co = net68047;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(net68047) );
endmodule


module FA_422 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_421 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  OR2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n7) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n7), .A2(n6), .ZN(S) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(n4), .ZN(n10) );
endmodule


module RCA_N4_106 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_424 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_423 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_422 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_421 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_420 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_419 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_418 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_417 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_105 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_420 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_419 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_418 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_417 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_53 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X2 U1 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U3 ( .A(sel), .ZN(n5) );
  INV_X1 U4 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[2]), .B1(B[2]), .B2(n14), .ZN(n17) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[1]), .B1(n5), .B2(B[1]), .ZN(n16) );
  INV_X1 U8 ( .A(sel), .ZN(n14) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n14), .ZN(n18) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n5), .B2(B[0]), .ZN(n15) );
endmodule


module carry_select_block_NPB4_53 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_106 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_105 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_53 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_416 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(n4), .ZN(n8) );
  CLKBUF_X1 U4 ( .A(B), .Z(n5) );
  XOR2_X1 U5 ( .A(n5), .B(A), .Z(n6) );
  AOI22_X1 U6 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_415 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_414 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_413 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_104 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_416 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_415 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_414 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_413 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_412 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_411 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_410 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_409 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_103 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_412 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_411 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_410 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_409 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_52 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U2 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U3 ( .A(sel), .ZN(n5) );
  INV_X1 U4 ( .A(n15), .ZN(Y[0]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[2]), .B1(n5), .B2(B[2]), .ZN(n17) );
  INV_X1 U6 ( .A(n16), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[1]), .B1(n5), .B2(B[1]), .ZN(n16) );
  INV_X1 U8 ( .A(sel), .ZN(n14) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n5), .ZN(n18) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n14), .B2(B[0]), .ZN(n15) );
endmodule


module carry_select_block_NPB4_52 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_104 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_103 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_52 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_408 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net68032, n4, n5, n6, n7;
  assign Co = net68032;

  XNOR2_X1 U1 ( .A(Ci), .B(A), .ZN(n7) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  OAI21_X1 U3 ( .B1(n4), .B2(n5), .A(n6), .ZN(net68032) );
  NAND2_X1 U4 ( .A1(Ci), .A2(B), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n7), .ZN(S) );
  NOR2_X1 U6 ( .A1(B), .A2(Ci), .ZN(n4) );
endmodule


module FA_407 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  AOI22_X1 U2 ( .A1(n4), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_406 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_405 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(n4), .ZN(n7) );
endmodule


module RCA_N4_102 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_408 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_407 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_406 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_405 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_404 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_403 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  XOR2_X1 U2 ( .A(A), .B(n4), .Z(n5) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(Ci), .B2(n7), .ZN(n8) );
endmodule


module FA_402 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_401 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_101 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_404 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_403 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_402 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_401 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_51 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X2 U1 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U2 ( .A(sel), .ZN(n5) );
  INV_X1 U3 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[2]), .B1(n5), .B2(B[2]), .ZN(n17) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[1]), .B1(n14), .B2(B[1]), .ZN(n16) );
  INV_X1 U7 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U8 ( .A(sel), .ZN(n14) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[3]), .B1(n5), .B2(B[3]), .ZN(n18) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n14), .B2(B[0]), .ZN(n15) );
endmodule


module carry_select_block_NPB4_51 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_102 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_101 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_51 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_400 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n7), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(n4), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n5), .B2(Ci), .ZN(n8) );
endmodule


module FA_399 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_398 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_397 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  OR2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_100 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_400 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_399 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_398 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_397 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_396 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_395 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_394 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_393 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_99 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_396 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_395 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_394 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_393 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_50 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n12, n13, n18, n19, n20, n21, n22;

  BUF_X1 U1 ( .A(n12), .Z(n13) );
  BUF_X1 U2 ( .A(sel), .Z(n12) );
  INV_X1 U3 ( .A(n13), .ZN(n5) );
  CLKBUF_X1 U4 ( .A(sel), .Z(n10) );
  INV_X2 U5 ( .A(n19), .ZN(Y[0]) );
  INV_X1 U6 ( .A(n12), .ZN(n11) );
  INV_X1 U7 ( .A(n21), .ZN(Y[2]) );
  INV_X1 U8 ( .A(n20), .ZN(Y[1]) );
  INV_X1 U9 ( .A(n22), .ZN(Y[3]) );
  AOI22_X1 U10 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(n5), .ZN(n21) );
  AOI22_X1 U11 ( .A1(n10), .A2(A[1]), .B1(B[1]), .B2(n11), .ZN(n20) );
  INV_X1 U12 ( .A(sel), .ZN(n18) );
  AOI22_X1 U13 ( .A1(A[3]), .A2(n13), .B1(B[3]), .B2(n5), .ZN(n22) );
  AOI22_X1 U14 ( .A1(sel), .A2(A[0]), .B1(n18), .B2(B[0]), .ZN(n19) );
endmodule


module carry_select_block_NPB4_50 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_100 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_99 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_50 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_392 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_391 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_390 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_389 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_98 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_392 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_391 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_390 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_389 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_388 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_387 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_386 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_385 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_97 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_388 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_387 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_386 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_385 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_49 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(n16), .ZN(Y[0]) );
  BUF_X1 U2 ( .A(n15), .Z(n5) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n10) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U6 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U7 ( .A(sel), .ZN(n15) );
  AOI22_X1 U8 ( .A1(n10), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U10 ( .A1(A[1]), .A2(n10), .B1(B[1]), .B2(n5), .ZN(n17) );
  AOI22_X1 U11 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n15), .ZN(n16) );
endmodule


module carry_select_block_NPB4_49 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_98 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_97 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_49 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_4 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_64 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_63 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_62 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_61 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_60 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_59 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_58 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_57 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_56 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_55 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_54 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), 
        .S(S[43:40]) );
  carry_select_block_NPB4_53 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), 
        .S(S[47:44]) );
  carry_select_block_NPB4_52 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), 
        .S(S[51:48]) );
  carry_select_block_NPB4_51 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), 
        .S(S[55:52]) );
  carry_select_block_NPB4_50 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), 
        .S(S[59:56]) );
  carry_select_block_NPB4_49 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), 
        .S(S[63:60]) );
endmodule


module P4_ADDER_N64_4 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_4 CGEN ( .A(A), .B({B[63:61], n4, B[59:57], n13, 
        B[55:49], n5, B[47:41], n3, B[39:29], n12, B[27:0]}), .Cin(Cin), .Co(
        CoutCgen) );
  sum_generator_N64_NPB4_4 SGEN ( .A(A), .B({B[63:56], n11, B[54:52], n9, 
        B[50:48], n2, B[46:44], n6, B[42:40], n10, B[38], n8, B[36:32], n1, 
        B[30:28], n7, B[26:0]}), .Ci({CoutCgen, Cin}), .S(S), .Co(Cout) );
  BUF_X1 U1 ( .A(B[31]), .Z(n1) );
  BUF_X2 U2 ( .A(B[37]), .Z(n8) );
  CLKBUF_X1 U3 ( .A(B[47]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(B[40]), .Z(n3) );
  CLKBUF_X1 U5 ( .A(B[60]), .Z(n4) );
  CLKBUF_X1 U6 ( .A(B[48]), .Z(n5) );
  CLKBUF_X1 U7 ( .A(B[43]), .Z(n6) );
  BUF_X1 U8 ( .A(B[28]), .Z(n12) );
  CLKBUF_X1 U9 ( .A(B[27]), .Z(n7) );
  CLKBUF_X1 U10 ( .A(B[51]), .Z(n9) );
  CLKBUF_X1 U11 ( .A(B[39]), .Z(n10) );
  CLKBUF_X1 U12 ( .A(B[55]), .Z(n11) );
  CLKBUF_X1 U13 ( .A(B[56]), .Z(n13) );
endmodule


module Booth_Encoder_3 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_3 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306;

  NAND2_X1 U1 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  NAND2_X1 U2 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  NAND2_X1 U3 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  AOI222_X1 U4 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n155), .ZN(n234) );
  NOR3_X1 U5 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U6 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  BUF_X1 U7 ( .A(n158), .Z(n161) );
  BUF_X1 U8 ( .A(n158), .Z(n162) );
  BUF_X1 U9 ( .A(n158), .Z(n160) );
  BUF_X1 U10 ( .A(n158), .Z(n163) );
  BUF_X1 U11 ( .A(n158), .Z(n159) );
  BUF_X1 U12 ( .A(n151), .Z(n153) );
  BUF_X1 U13 ( .A(n151), .Z(n155) );
  BUF_X1 U14 ( .A(n165), .Z(n167) );
  BUF_X1 U15 ( .A(n165), .Z(n169) );
  BUF_X1 U16 ( .A(n151), .Z(n154) );
  BUF_X1 U17 ( .A(n165), .Z(n168) );
  BUF_X1 U18 ( .A(n303), .Z(n158) );
  NOR4_X1 U19 ( .A1(n150), .A2(n144), .A3(n153), .A4(n167), .ZN(n303) );
  BUF_X1 U20 ( .A(n152), .Z(n157) );
  BUF_X1 U21 ( .A(n166), .Z(n171) );
  BUF_X1 U22 ( .A(n152), .Z(n156) );
  BUF_X1 U23 ( .A(n166), .Z(n170) );
  BUF_X1 U24 ( .A(n301), .Z(n148) );
  BUF_X1 U25 ( .A(n304), .Z(n165) );
  BUF_X1 U26 ( .A(n302), .Z(n151) );
  BUF_X1 U27 ( .A(n301), .Z(n147) );
  BUF_X1 U28 ( .A(n301), .Z(n145) );
  BUF_X1 U29 ( .A(n301), .Z(n146) );
  BUF_X1 U30 ( .A(n304), .Z(n166) );
  BUF_X1 U31 ( .A(n302), .Z(n152) );
  BUF_X1 U32 ( .A(n301), .Z(n149) );
  BUF_X1 U33 ( .A(n300), .Z(n141) );
  BUF_X1 U34 ( .A(n300), .Z(n143) );
  BUF_X1 U35 ( .A(n300), .Z(n139) );
  BUF_X1 U36 ( .A(n300), .Z(n142) );
  BUF_X1 U37 ( .A(n300), .Z(n140) );
  INV_X1 U38 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U39 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n304) );
  AND3_X1 U40 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U41 ( .A(sel[2]), .ZN(n173) );
  NAND2_X1 U42 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  NAND2_X1 U43 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  NAND2_X1 U44 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  NAND2_X1 U45 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U46 ( .A1(C[60]), .A2(n145), .B1(A[60]), .B2(n139), .ZN(n287) );
  AOI222_X1 U47 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n157), .ZN(n286) );
  NAND2_X1 U48 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  AOI22_X1 U49 ( .A1(C[56]), .A2(n146), .B1(A[56]), .B2(n140), .ZN(n277) );
  AOI222_X1 U50 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n157), .ZN(n276) );
  AOI222_X1 U51 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n154), .ZN(n212) );
  AOI222_X1 U52 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n154), .ZN(n210) );
  NAND2_X1 U53 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  AOI22_X1 U54 ( .A1(C[28]), .A2(n148), .B1(A[28]), .B2(n142), .ZN(n215) );
  NAND2_X1 U55 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI22_X1 U56 ( .A1(C[29]), .A2(n148), .B1(A[29]), .B2(n142), .ZN(n217) );
  NAND2_X1 U57 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U58 ( .A1(C[30]), .A2(n148), .B1(A[30]), .B2(n142), .ZN(n221) );
  NAND2_X1 U59 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI22_X1 U60 ( .A1(C[31]), .A2(n148), .B1(A[31]), .B2(n142), .ZN(n223) );
  NAND2_X1 U61 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI22_X1 U62 ( .A1(C[34]), .A2(n148), .B1(A[34]), .B2(n142), .ZN(n229) );
  AOI222_X1 U63 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n155), .ZN(n228) );
  NAND2_X1 U64 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI22_X1 U65 ( .A1(C[38]), .A2(n147), .B1(A[38]), .B2(n141), .ZN(n237) );
  AOI222_X1 U66 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n155), .ZN(n236) );
  NAND2_X1 U67 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI22_X1 U68 ( .A1(C[42]), .A2(n147), .B1(A[42]), .B2(n141), .ZN(n247) );
  AOI222_X1 U69 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n155), .ZN(n246) );
  NAND2_X1 U70 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI22_X1 U71 ( .A1(C[46]), .A2(n146), .B1(A[46]), .B2(n140), .ZN(n255) );
  AOI222_X1 U72 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n156), .ZN(n254) );
  NAND2_X1 U73 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U74 ( .A1(C[63]), .A2(n145), .B1(A[63]), .B2(n139), .ZN(n293) );
  AOI222_X1 U75 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n157), .ZN(n292) );
  NAND2_X1 U76 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  AOI22_X1 U77 ( .A1(C[32]), .A2(n148), .B1(A[32]), .B2(n142), .ZN(n225) );
  AOI222_X1 U78 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n155), .ZN(n224) );
  AOI22_X1 U79 ( .A1(C[48]), .A2(n146), .B1(A[48]), .B2(n140), .ZN(n259) );
  AOI222_X1 U80 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n156), .ZN(n258) );
  NAND2_X1 U81 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI22_X1 U82 ( .A1(C[33]), .A2(n148), .B1(A[33]), .B2(n142), .ZN(n227) );
  AOI222_X1 U83 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n155), .ZN(n226) );
  NAND2_X1 U84 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI22_X1 U85 ( .A1(C[37]), .A2(n147), .B1(A[37]), .B2(n141), .ZN(n235) );
  NAND2_X1 U86 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI22_X1 U87 ( .A1(C[35]), .A2(n148), .B1(A[35]), .B2(n142), .ZN(n231) );
  AOI222_X1 U88 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n155), .ZN(n230) );
  NAND2_X1 U89 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI222_X1 U90 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n155), .ZN(n238) );
  AOI22_X1 U91 ( .A1(C[39]), .A2(n147), .B1(A[39]), .B2(n141), .ZN(n239) );
  NAND2_X1 U92 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI22_X1 U93 ( .A1(C[50]), .A2(n146), .B1(A[50]), .B2(n140), .ZN(n265) );
  NAND2_X1 U94 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  NAND2_X1 U95 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U96 ( .A1(C[61]), .A2(n145), .B1(A[61]), .B2(n139), .ZN(n289) );
  AOI222_X1 U97 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n157), .ZN(n288) );
  NAND2_X1 U98 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  AOI22_X1 U99 ( .A1(C[36]), .A2(n147), .B1(A[36]), .B2(n141), .ZN(n233) );
  AOI222_X1 U100 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n155), .ZN(n232) );
  AOI222_X1 U101 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n155), .ZN(n242) );
  AOI22_X1 U102 ( .A1(C[40]), .A2(n147), .B1(A[40]), .B2(n141), .ZN(n243) );
  NAND2_X1 U103 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U104 ( .A1(C[62]), .A2(n145), .B1(A[62]), .B2(n139), .ZN(n291) );
  AOI222_X1 U105 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n157), .ZN(n290) );
  NAND2_X1 U106 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI222_X1 U107 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n157), .ZN(n280) );
  AOI22_X1 U108 ( .A1(C[58]), .A2(n145), .B1(A[58]), .B2(n139), .ZN(n281) );
  NAND2_X1 U109 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI222_X1 U110 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n155), .ZN(n244) );
  AOI22_X1 U111 ( .A1(C[41]), .A2(n147), .B1(A[41]), .B2(n141), .ZN(n245) );
  NAND2_X1 U112 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI222_X1 U113 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n156), .ZN(n252) );
  AOI22_X1 U114 ( .A1(C[45]), .A2(n147), .B1(A[45]), .B2(n141), .ZN(n253) );
  AOI222_X1 U115 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n156), .ZN(n250) );
  AOI22_X1 U116 ( .A1(C[44]), .A2(n147), .B1(A[44]), .B2(n141), .ZN(n251) );
  NAND2_X1 U117 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI222_X1 U118 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n156), .ZN(n256) );
  AOI22_X1 U119 ( .A1(C[47]), .A2(n146), .B1(A[47]), .B2(n140), .ZN(n257) );
  NAND2_X1 U120 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  AOI222_X1 U121 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n156), .ZN(n266) );
  AOI22_X1 U122 ( .A1(C[51]), .A2(n146), .B1(A[51]), .B2(n140), .ZN(n267) );
  NAND2_X1 U123 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  AOI22_X1 U124 ( .A1(C[52]), .A2(n146), .B1(A[52]), .B2(n140), .ZN(n269) );
  AOI222_X1 U125 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n156), .ZN(n268) );
  NAND2_X1 U126 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U127 ( .A1(C[59]), .A2(n145), .B1(A[59]), .B2(n139), .ZN(n283) );
  AOI222_X1 U128 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n157), .ZN(n282) );
  NAND2_X1 U129 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI222_X1 U130 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n155), .ZN(n248) );
  AOI22_X1 U131 ( .A1(C[43]), .A2(n147), .B1(A[43]), .B2(n141), .ZN(n249) );
  NAND2_X1 U132 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI22_X1 U133 ( .A1(C[55]), .A2(n146), .B1(A[55]), .B2(n140), .ZN(n275) );
  AOI222_X1 U134 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n156), .ZN(n274) );
  NAND2_X1 U135 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U136 ( .A1(C[0]), .A2(n145), .B1(A[0]), .B2(n139), .ZN(n175) );
  AOI222_X1 U137 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n153), .ZN(n174) );
  NAND2_X1 U138 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U139 ( .A1(C[4]), .A2(n146), .B1(A[4]), .B2(n140), .ZN(n263) );
  AOI222_X1 U140 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n156), .ZN(n262) );
  NAND2_X1 U141 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI22_X1 U142 ( .A1(C[8]), .A2(n145), .B1(A[8]), .B2(n139), .ZN(n299) );
  AOI222_X1 U143 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n157), .ZN(n298) );
  NAND2_X1 U144 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  AOI22_X1 U145 ( .A1(C[12]), .A2(n150), .B1(A[12]), .B2(n144), .ZN(n181) );
  AOI222_X1 U146 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n153), .ZN(n180) );
  NAND2_X1 U147 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  AOI22_X1 U148 ( .A1(C[16]), .A2(n149), .B1(A[16]), .B2(n143), .ZN(n189) );
  AOI222_X1 U149 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n153), .ZN(n188) );
  NAND2_X1 U150 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  AOI22_X1 U151 ( .A1(C[20]), .A2(n149), .B1(A[20]), .B2(n143), .ZN(n199) );
  AOI222_X1 U152 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n154), .ZN(n198) );
  NAND2_X1 U153 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  AOI22_X1 U154 ( .A1(C[24]), .A2(n149), .B1(A[24]), .B2(n143), .ZN(n207) );
  AOI222_X1 U155 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n154), .ZN(n206) );
  NAND2_X1 U156 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U157 ( .A1(C[1]), .A2(n149), .B1(A[1]), .B2(n143), .ZN(n197) );
  AOI222_X1 U158 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n153), .ZN(n196) );
  NAND2_X1 U159 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U160 ( .A1(C[5]), .A2(n145), .B1(A[5]), .B2(n139), .ZN(n285) );
  AOI222_X1 U161 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n157), .ZN(n284) );
  NAND2_X1 U162 ( .A1(n306), .A2(n305), .ZN(Y[9]) );
  AOI22_X1 U163 ( .A1(C[9]), .A2(n147), .B1(A[9]), .B2(n141), .ZN(n306) );
  AOI222_X1 U164 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n157), .ZN(n305) );
  NAND2_X1 U165 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U166 ( .A1(C[13]), .A2(n150), .B1(A[13]), .B2(n144), .ZN(n183) );
  AOI222_X1 U167 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n153), .ZN(n182) );
  NAND2_X1 U168 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI22_X1 U169 ( .A1(C[17]), .A2(n149), .B1(A[17]), .B2(n143), .ZN(n191) );
  AOI222_X1 U170 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n153), .ZN(n190) );
  NAND2_X1 U171 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI22_X1 U172 ( .A1(C[21]), .A2(n149), .B1(A[21]), .B2(n143), .ZN(n201) );
  AOI222_X1 U173 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n154), .ZN(n200) );
  NAND2_X1 U174 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI22_X1 U175 ( .A1(C[25]), .A2(n148), .B1(A[25]), .B2(n142), .ZN(n209) );
  AOI222_X1 U176 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n154), .ZN(n208) );
  NAND2_X1 U177 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U178 ( .A1(C[2]), .A2(n148), .B1(A[2]), .B2(n142), .ZN(n219) );
  AOI222_X1 U179 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n154), .ZN(n218) );
  NAND2_X1 U180 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U181 ( .A1(C[6]), .A2(n145), .B1(A[6]), .B2(n139), .ZN(n295) );
  AOI222_X1 U182 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n157), .ZN(n294) );
  NAND2_X1 U183 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U184 ( .A1(C[10]), .A2(n150), .B1(A[10]), .B2(n144), .ZN(n177) );
  AOI222_X1 U185 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n153), .ZN(n176) );
  NAND2_X1 U186 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U187 ( .A1(C[14]), .A2(n149), .B1(A[14]), .B2(n143), .ZN(n185) );
  AOI222_X1 U188 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n153), .ZN(n184) );
  NAND2_X1 U189 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI22_X1 U190 ( .A1(C[18]), .A2(n149), .B1(A[18]), .B2(n143), .ZN(n193) );
  AOI222_X1 U191 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n153), .ZN(n192) );
  NAND2_X1 U192 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI22_X1 U193 ( .A1(C[22]), .A2(n149), .B1(A[22]), .B2(n143), .ZN(n203) );
  AOI222_X1 U194 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n154), .ZN(n202) );
  NAND2_X1 U195 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U196 ( .A1(C[3]), .A2(n147), .B1(A[3]), .B2(n141), .ZN(n241) );
  AOI222_X1 U197 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n155), .ZN(n240) );
  NAND2_X1 U198 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U199 ( .A1(C[7]), .A2(n145), .B1(A[7]), .B2(n139), .ZN(n297) );
  AOI222_X1 U200 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n157), .ZN(n296) );
  NAND2_X1 U201 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U202 ( .A1(C[11]), .A2(n150), .B1(A[11]), .B2(n144), .ZN(n179) );
  AOI222_X1 U203 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n153), .ZN(n178) );
  NAND2_X1 U204 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U205 ( .A1(C[15]), .A2(n149), .B1(A[15]), .B2(n143), .ZN(n187) );
  AOI222_X1 U206 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n153), .ZN(n186) );
  NAND2_X1 U207 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI22_X1 U208 ( .A1(C[19]), .A2(n149), .B1(A[19]), .B2(n143), .ZN(n195) );
  AOI222_X1 U209 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n153), .ZN(n194) );
  NAND2_X1 U210 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI22_X1 U211 ( .A1(C[23]), .A2(n149), .B1(A[23]), .B2(n143), .ZN(n205) );
  AOI222_X1 U212 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n154), .ZN(n204) );
  AOI22_X1 U213 ( .A1(C[54]), .A2(n146), .B1(A[54]), .B2(n140), .ZN(n273) );
  AOI22_X1 U214 ( .A1(C[53]), .A2(n146), .B1(A[53]), .B2(n140), .ZN(n271) );
  AOI222_X1 U215 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n156), .ZN(n270) );
  AOI22_X1 U216 ( .A1(C[26]), .A2(n148), .B1(A[26]), .B2(n142), .ZN(n211) );
  AOI22_X1 U217 ( .A1(C[27]), .A2(n148), .B1(A[27]), .B2(n142), .ZN(n213) );
  NAND2_X1 U218 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  NAND2_X1 U219 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI222_X1 U220 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n154), .ZN(n222) );
  AOI222_X1 U221 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n154), .ZN(n220) );
  AOI22_X1 U222 ( .A1(C[49]), .A2(n146), .B1(A[49]), .B2(n140), .ZN(n261) );
  AOI222_X1 U223 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n156), .ZN(n272) );
  AOI222_X1 U224 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n156), .ZN(n260) );
  AOI222_X1 U225 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n156), .ZN(n264) );
  AOI22_X1 U226 ( .A1(C[57]), .A2(n145), .B1(A[57]), .B2(n139), .ZN(n279) );
  AOI222_X1 U227 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n157), .ZN(n278) );
  AOI222_X1 U228 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n154), .ZN(n214) );
  AOI222_X1 U229 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n154), .ZN(n216) );
  CLKBUF_X1 U230 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U231 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U232 ( .A(n158), .Z(n164) );
endmodule


module G_51 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_189 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_188 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_187 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_186 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_185 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_184 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_183 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_182 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_181 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_180 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_179 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_178 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_177 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_176 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_175 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_174 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_173 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_172 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_171 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_170 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_169 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n3, n5;

  CLKBUF_X1 U1 ( .A(P_IK), .Z(n3) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n5) );
  AND2_X1 U3 ( .A1(n3), .A2(P_K_1), .ZN(Px) );
  INV_X1 U4 ( .A(n5), .ZN(Gx) );
endmodule


module PG_168 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_167 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_166 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_165 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_164 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_163 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_162 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_161 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_160 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_159 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_50 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_158 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_157 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_156 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_155 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_154 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_153 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_152 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_151 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_150 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_149 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_148 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_147 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_146 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_145 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_144 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_49 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_143 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_142 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_141 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_140 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_139 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_138 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_137 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_48 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_47 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_136 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_135 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_134 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_133 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_132 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_131 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module G_46 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_45 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_44 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_43 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_130 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_129 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_128 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_127 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module G_42 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_41 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_40 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_39 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_38 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_37 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_36 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n3, n5;

  AND2_X1 U1 ( .A1(P_IK), .A2(G_K_1), .ZN(n3) );
  NOR2_X1 U2 ( .A1(n3), .A2(G_IK), .ZN(n5) );
  INV_X1 U3 ( .A(n5), .ZN(Gx) );
endmodule


module G_35 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
endmodule


module carry_generator_N64_NPB4_3 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   n27, \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U83 ( .A(B[53]), .B(A[53]), .Z(\PG_Network[0][0][53] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U100 ( .A(B[38]), .B(A[38]), .Z(\PG_Network[0][0][38] ) );
  XOR2_X1 U101 ( .A(B[37]), .B(A[37]), .Z(\PG_Network[0][0][37] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U103 ( .A(B[35]), .B(A[35]), .Z(\PG_Network[0][0][35] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U108 ( .A(B[30]), .B(A[30]), .Z(\PG_Network[0][0][30] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U110 ( .A(B[29]), .B(A[29]), .Z(\PG_Network[0][0][29] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U112 ( .A(B[27]), .B(A[27]), .Z(\PG_Network[0][0][27] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U114 ( .A(B[25]), .B(A[25]), .Z(\PG_Network[0][0][25] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U116 ( .A(B[23]), .B(A[23]), .Z(\PG_Network[0][0][23] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U121 ( .A(B[19]), .B(A[19]), .Z(\PG_Network[0][0][19] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U125 ( .A(B[15]), .B(A[15]), .Z(\PG_Network[0][0][15] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_51 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n23), .Gx(\PG_Network[1][1][1] ) );
  PG_189 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_188 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_187 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_186 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_185 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_184 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_183 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_182 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_181 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_180 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_179 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_178 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_177 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_176 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_175 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_174 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_173 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_172 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_171 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_170 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_169 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_168 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_167 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_166 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_165 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_164 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_163 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_162 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_161 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_160 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_159 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_50 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_158 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_157 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_156 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_155 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_154 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_153 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_152 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_151 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_150 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_149 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_148 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_147 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_146 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_145 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_144 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_49 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_143 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_142 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_141 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_140 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_139 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_138 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_137 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_48 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), 
        .G_K_1(Co[1]), .Gx(Co[3]) );
  G_47 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), 
        .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_136 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_135 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_134 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][47] ), .Px(
        \PG_Network[4][0][47] ) );
  PG_133 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(
        \PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][43] ), .Px(
        \PG_Network[4][0][43] ) );
  PG_132 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(n11), .P_K_1(n13), .Gx(
        \PG_Network[4][1][63] ), .Px(\PG_Network[4][0][63] ) );
  PG_131 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(n11), .P_K_1(n13), .Gx(
        \PG_Network[4][1][59] ), .Px(\PG_Network[4][0][59] ) );
  G_46 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), 
        .G_K_1(Co[3]), .Gx(n27) );
  G_45 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), 
        .G_K_1(Co[3]), .Gx(Co[6]) );
  G_44 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), 
        .G_K_1(Co[3]), .Gx(Co[5]) );
  G_43 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), 
        .G_K_1(Co[3]), .Gx(Co[4]) );
  PG_130 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(n17), .P_K_1(n7), .Gx(
        \PG_Network[5][1][63] ), .Px(\PG_Network[5][0][63] ) );
  PG_129 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(n17), .P_K_1(n7), .Gx(
        \PG_Network[5][1][59] ), .Px(\PG_Network[5][0][59] ) );
  PG_128 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(n9), .P_K_1(n7), .Gx(
        \PG_Network[5][1][55] ), .Px(\PG_Network[5][0][55] ) );
  PG_127 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][51] ), .Px(
        \PG_Network[5][0][51] ) );
  G_42 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), 
        .G_K_1(n10), .Gx(Co[15]) );
  G_41 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), 
        .G_K_1(n10), .Gx(Co[14]) );
  G_40 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), 
        .G_K_1(n10), .Gx(Co[13]) );
  G_39 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), 
        .G_K_1(n10), .Gx(Co[12]) );
  G_38 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), 
        .G_K_1(n10), .Gx(Co[11]) );
  G_37 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), 
        .G_K_1(Co[7]), .Gx(Co[10]) );
  G_36 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), 
        .G_K_1(n27), .Gx(Co[9]) );
  G_35 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), 
        .G_K_1(n27), .Gx(Co[8]) );
  INV_X1 U1 ( .A(A[31]), .ZN(n12) );
  INV_X1 U2 ( .A(A[46]), .ZN(n6) );
  INV_X1 U3 ( .A(A[45]), .ZN(n16) );
  INV_X1 U4 ( .A(A[49]), .ZN(n14) );
  INV_X1 U5 ( .A(A[47]), .ZN(n19) );
  INV_X1 U6 ( .A(A[51]), .ZN(n18) );
  INV_X1 U7 ( .A(A[43]), .ZN(n15) );
  INV_X1 U8 ( .A(A[55]), .ZN(n21) );
  INV_X1 U9 ( .A(A[39]), .ZN(n20) );
  INV_X1 U10 ( .A(A[59]), .ZN(n22) );
  INV_X1 U11 ( .A(A[48]), .ZN(n5) );
  XNOR2_X1 U12 ( .A(n5), .B(B[48]), .ZN(\PG_Network[0][0][48] ) );
  XNOR2_X1 U13 ( .A(B[46]), .B(n6), .ZN(\PG_Network[0][0][46] ) );
  CLKBUF_X1 U14 ( .A(\PG_Network[4][0][47] ), .Z(n7) );
  BUF_X2 U15 ( .A(n27), .Z(Co[7]) );
  CLKBUF_X1 U16 ( .A(\PG_Network[4][1][47] ), .Z(n9) );
  CLKBUF_X1 U17 ( .A(n27), .Z(n10) );
  CLKBUF_X1 U18 ( .A(\PG_Network[3][1][55] ), .Z(n11) );
  XNOR2_X1 U19 ( .A(B[31]), .B(n12), .ZN(\PG_Network[0][0][31] ) );
  CLKBUF_X1 U20 ( .A(\PG_Network[3][0][55] ), .Z(n13) );
  XNOR2_X1 U21 ( .A(B[49]), .B(n14), .ZN(\PG_Network[0][0][49] ) );
  XNOR2_X1 U22 ( .A(B[43]), .B(n15), .ZN(\PG_Network[0][0][43] ) );
  XNOR2_X1 U23 ( .A(B[45]), .B(n16), .ZN(\PG_Network[0][0][45] ) );
  CLKBUF_X1 U24 ( .A(n9), .Z(n17) );
  XNOR2_X1 U25 ( .A(B[51]), .B(n18), .ZN(\PG_Network[0][0][51] ) );
  XNOR2_X1 U26 ( .A(B[47]), .B(n19), .ZN(\PG_Network[0][0][47] ) );
  XNOR2_X1 U27 ( .A(B[39]), .B(n20), .ZN(\PG_Network[0][0][39] ) );
  XNOR2_X1 U28 ( .A(B[55]), .B(n21), .ZN(\PG_Network[0][0][55] ) );
  XNOR2_X1 U29 ( .A(B[59]), .B(n22), .ZN(\PG_Network[0][0][59] ) );
  AND2_X1 U30 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U31 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U32 ( .A1(A[41]), .A2(B[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U33 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U34 ( .A1(A[35]), .A2(B[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U35 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U36 ( .A1(A[31]), .A2(B[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U37 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U38 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U39 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U40 ( .A1(B[49]), .A2(A[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U41 ( .A1(B[48]), .A2(A[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U42 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U43 ( .A1(B[51]), .A2(A[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U44 ( .A1(A[46]), .A2(B[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U45 ( .A1(B[47]), .A2(A[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U46 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U47 ( .A1(A[27]), .A2(B[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U48 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U49 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U50 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U51 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U52 ( .A1(A[45]), .A2(B[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U53 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U54 ( .A1(A[29]), .A2(B[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U55 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U56 ( .A1(A[37]), .A2(B[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U57 ( .A1(B[53]), .A2(A[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U58 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U59 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U60 ( .A1(A[19]), .A2(B[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U61 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U62 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U63 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U64 ( .A1(A[11]), .A2(B[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U65 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U66 ( .A1(A[15]), .A2(B[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U67 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U77 ( .A1(A[25]), .A2(B[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U81 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U85 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U88 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U89 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U90 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U91 ( .A(n26), .ZN(n23) );
  AND2_X1 U92 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U94 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U99 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U107 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U131 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U132 ( .A1(A[7]), .A2(B[7]), .ZN(\PG_Network[0][1][7] ) );
  AND2_X1 U133 ( .A1(A[21]), .A2(B[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U134 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U135 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U136 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AND2_X1 U137 ( .A1(A[23]), .A2(B[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U138 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AOI21_X1 U139 ( .B1(A[0]), .B2(B[0]), .A(n24), .ZN(n26) );
  INV_X1 U140 ( .A(n25), .ZN(n24) );
  OAI21_X1 U141 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n25) );
  AND2_X1 U142 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
  AND2_X1 U143 ( .A1(A[52]), .A2(B[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U144 ( .A1(B[43]), .A2(A[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U145 ( .A1(B[44]), .A2(A[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U146 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U147 ( .A1(B[55]), .A2(A[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U148 ( .A1(B[59]), .A2(A[59]), .ZN(\PG_Network[0][1][59] ) );
endmodule


module FA_384 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_383 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_382 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_381 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_96 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_384 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_383 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_382 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_381 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_380 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_379 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_378 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_377 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_95 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_380 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_379 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_378 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_377 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_48 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U2 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U4 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U5 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U7 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_48 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_96 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_95 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_48 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_376 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_375 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_374 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_373 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_94 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_376 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_375 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_374 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_373 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_372 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_371 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_370 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_369 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_93 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_372 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_371 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_370 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_369 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_47 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_47 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_94 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_93 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_47 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_368 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_367 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_366 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_365 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_92 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_368 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_367 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_366 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_365 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_364 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_363 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_362 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_361 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_91 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_364 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_363 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_362 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_361 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_46 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_46 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_92 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_91 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_46 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_360 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_359 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_358 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_357 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_90 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_360 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_359 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_358 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_357 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_356 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_355 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_354 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_353 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_89 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_356 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_355 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_354 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_353 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_45 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_45 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_90 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_89 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_45 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_352 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_351 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_350 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_349 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_88 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_352 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_351 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_350 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_349 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_348 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_347 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_346 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_345 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_87 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_348 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_347 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_346 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_345 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_44 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_44 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_88 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_87 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_44 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_344 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_343 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_342 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_341 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_86 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_344 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_343 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_342 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_341 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_340 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_339 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_338 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_337 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_85 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_340 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_339 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_338 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_337 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_43 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_43 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_86 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_85 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_43 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_336 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_335 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_334 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_333 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_84 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_336 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_335 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_334 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_333 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_332 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_331 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_330 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_329 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_83 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_332 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_331 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_330 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_329 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_42 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_42 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_84 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_83 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_42 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_328 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_327 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_326 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_325 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_82 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_328 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_327 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_326 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_325 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_324 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_323 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_322 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_321 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_81 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_324 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_323 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_322 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_321 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_41 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U3 ( .A(sel), .ZN(n13) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_41 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_82 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_81 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_41 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_320 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_319 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_318 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_317 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_80 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_320 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_319 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_318 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_317 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_316 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_315 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_314 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_313 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_79 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_316 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_315 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_314 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_313 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_40 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U5 ( .A(sel), .ZN(n13) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_40 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_80 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_79 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_40 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_312 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_311 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_310 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_309 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_78 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_312 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_311 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_310 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_309 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_308 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_307 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_306 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_305 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_77 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_308 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_307 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_306 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_305 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_39 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n13), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(sel), .ZN(n13) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n13), .ZN(n17) );
endmodule


module carry_select_block_NPB4_39 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_78 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_77 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_39 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_304 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_303 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_302 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_301 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  OR2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_76 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_304 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_303 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_302 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_301 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_300 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_299 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_298 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_297 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_75 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_300 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_299 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_298 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_297 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_38 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  BUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U6 ( .A(sel), .ZN(n14) );
  AOI22_X1 U7 ( .A1(n5), .A2(A[2]), .B1(B[2]), .B2(n14), .ZN(n17) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n14), .ZN(n15) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n14), .ZN(n18) );
endmodule


module carry_select_block_NPB4_38 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_76 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_75 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_38 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_296 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n5) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  XOR2_X1 U5 ( .A(n4), .B(A), .Z(n6) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n9) );
endmodule


module FA_295 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_294 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_293 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_74 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_296 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_295 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_294 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_293 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_292 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_291 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_290 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_289 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_73 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_292 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_291 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_290 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_289 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_37 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U4 ( .A(sel), .ZN(n5) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n16) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n5), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n5), .ZN(n14) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n5), .ZN(n17) );
endmodule


module carry_select_block_NPB4_37 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_74 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_73 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_37 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_288 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_287 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_286 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_285 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  OR2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n6) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n8) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_72 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_288 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_287 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_286 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_285 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_284 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_283 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_282 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_281 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_71 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_284 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_283 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_282 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_281 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_36 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19, n20;

  CLKBUF_X1 U1 ( .A(sel), .Z(n5) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n10) );
  INV_X1 U3 ( .A(sel), .ZN(n11) );
  INV_X1 U4 ( .A(n20), .ZN(Y[3]) );
  INV_X1 U5 ( .A(n19), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n18), .ZN(Y[1]) );
  INV_X1 U7 ( .A(n17), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n11), .ZN(n19) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(sel), .B1(n16), .B2(B[1]), .ZN(n18) );
  AOI22_X1 U10 ( .A1(n10), .A2(A[3]), .B1(B[3]), .B2(n11), .ZN(n20) );
  AOI22_X1 U11 ( .A1(A[0]), .A2(sel), .B1(n16), .B2(B[0]), .ZN(n17) );
  INV_X1 U12 ( .A(sel), .ZN(n16) );
endmodule


module carry_select_block_NPB4_36 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_72 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_71 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_36 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_280 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net67904, n4, n5, n6, n7;
  assign Co = net67904;

  INV_X1 U1 ( .A(Ci), .ZN(n6) );
  CLKBUF_X1 U2 ( .A(n5), .Z(n4) );
  XNOR2_X1 U3 ( .A(n4), .B(Ci), .ZN(S) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n7) );
  OAI21_X1 U5 ( .B1(n5), .B2(n6), .A(n7), .ZN(net67904) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n5) );
endmodule


module FA_279 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_278 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_277 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  OR2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n6) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n8) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_70 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_280 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_279 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_278 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_277 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_276 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_275 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_274 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_273 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_69 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_276 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_275 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_274 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_273 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_35 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n11, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(n11), .Z(n5) );
  INV_X2 U2 ( .A(n17), .ZN(Y[1]) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n10) );
  INV_X1 U4 ( .A(sel), .ZN(n11) );
  INV_X1 U5 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U6 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U7 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[1]), .B1(n11), .B2(B[1]), .ZN(n17) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n11), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_35 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_70 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_69 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_35 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_272 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net67896, n4, n5, n6, n7;
  assign Co = net67896;

  INV_X1 U1 ( .A(Ci), .ZN(n6) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n4) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n7) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n5) );
  XNOR2_X1 U5 ( .A(Ci), .B(n4), .ZN(S) );
  OAI21_X1 U6 ( .B1(n5), .B2(n6), .A(n7), .ZN(net67896) );
endmodule


module FA_271 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n5), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n5) );
  CLKBUF_X1 U5 ( .A(n8), .Z(n6) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(Ci), .B2(n8), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_270 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_269 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n5) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n4), .B2(Ci), .ZN(n8) );
endmodule


module RCA_N4_68 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_272 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_271 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_270 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_269 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_268 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_267 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_266 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_265 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n4) );
  XNOR2_X1 U2 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U3 ( .A(n6), .B(B), .ZN(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n8) );
endmodule


module RCA_N4_67 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_268 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_267 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_266 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_265 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_34 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(sel), .ZN(n5) );
  INV_X1 U2 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[2]), .B1(B[2]), .B2(n5), .ZN(n17) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[1]), .B1(n5), .B2(B[1]), .ZN(n16) );
  INV_X1 U8 ( .A(sel), .ZN(n14) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n5), .ZN(n18) );
  AOI22_X1 U10 ( .A1(sel), .A2(A[0]), .B1(n14), .B2(B[0]), .ZN(n15) );
endmodule


module carry_select_block_NPB4_34 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_68 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_67 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_34 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_264 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_263 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_262 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_261 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module RCA_N4_66 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_264 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_263 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_262 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_261 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_260 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_259 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_258 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_257 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module RCA_N4_65 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_260 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_259 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_258 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_257 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_33 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X1 U1 ( .A(sel), .ZN(n5) );
  INV_X1 U2 ( .A(n19), .ZN(Y[3]) );
  INV_X1 U3 ( .A(n18), .ZN(Y[2]) );
  CLKBUF_X1 U4 ( .A(sel), .Z(n10) );
  INV_X1 U5 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U6 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n15), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(n10), .B1(B[1]), .B2(n15), .ZN(n17) );
  INV_X1 U9 ( .A(sel), .ZN(n15) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n15), .ZN(n19) );
  AOI22_X1 U11 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n5), .ZN(n16) );
endmodule


module carry_select_block_NPB4_33 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_66 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_65 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_33 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_3 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_48 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_47 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_46 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_45 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_44 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_43 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_42 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_41 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_40 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_39 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_38 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), 
        .S(S[43:40]) );
  carry_select_block_NPB4_37 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), 
        .S(S[47:44]) );
  carry_select_block_NPB4_36 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), 
        .S(S[51:48]) );
  carry_select_block_NPB4_35 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), 
        .S(S[55:52]) );
  carry_select_block_NPB4_34 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), 
        .S(S[59:56]) );
  carry_select_block_NPB4_33 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), 
        .S(S[63:60]) );
endmodule


module P4_ADDER_N64_3 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_3 CGEN ( .A(A), .B({B[63:61], n8, B[59:58], n10, 
        n16, B[55:49], n17, B[47:0]}), .Cin(Cin), .Co(CoutCgen) );
  sum_generator_N64_NPB4_3 SGEN ( .A(A), .B({B[63:60], n2, B[58:54], n9, B[52], 
        n12, B[50:48], n11, n1, n7, B[44], n13, B[42], n3, B[40], n6, B[38:36], 
        n4, B[34:32], n15, B[30:0]}), .Ci({CoutCgen, Cin}), .S(S), .Co(Cout)
         );
  BUF_X1 U1 ( .A(B[41]), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B[48]), .Z(n17) );
  CLKBUF_X1 U3 ( .A(B[46]), .Z(n1) );
  BUF_X1 U4 ( .A(B[45]), .Z(n7) );
  BUF_X1 U5 ( .A(B[59]), .Z(n2) );
  BUF_X2 U6 ( .A(B[53]), .Z(n9) );
  CLKBUF_X1 U7 ( .A(B[35]), .Z(n4) );
  INV_X1 U8 ( .A(B[39]), .ZN(n5) );
  INV_X1 U9 ( .A(n5), .ZN(n6) );
  CLKBUF_X1 U10 ( .A(B[60]), .Z(n8) );
  CLKBUF_X1 U11 ( .A(B[57]), .Z(n10) );
  CLKBUF_X1 U12 ( .A(B[47]), .Z(n11) );
  CLKBUF_X1 U13 ( .A(B[51]), .Z(n12) );
  CLKBUF_X1 U14 ( .A(B[43]), .Z(n13) );
  INV_X1 U15 ( .A(B[31]), .ZN(n14) );
  INV_X1 U16 ( .A(n14), .ZN(n15) );
  CLKBUF_X1 U17 ( .A(B[56]), .Z(n16) );
endmodule


module Booth_Encoder_2 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_2 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306;

  NAND2_X1 U1 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  NAND2_X1 U2 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  NOR3_X1 U3 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U4 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  NAND2_X1 U5 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  NAND2_X1 U6 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI222_X1 U7 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n155), .ZN(n238) );
  BUF_X1 U8 ( .A(n158), .Z(n160) );
  BUF_X1 U9 ( .A(n158), .Z(n161) );
  BUF_X1 U10 ( .A(n158), .Z(n162) );
  BUF_X1 U11 ( .A(n158), .Z(n163) );
  BUF_X1 U12 ( .A(n158), .Z(n159) );
  BUF_X1 U13 ( .A(n151), .Z(n153) );
  BUF_X1 U14 ( .A(n165), .Z(n167) );
  BUF_X1 U15 ( .A(n151), .Z(n155) );
  BUF_X1 U16 ( .A(n165), .Z(n169) );
  BUF_X1 U17 ( .A(n152), .Z(n157) );
  BUF_X1 U18 ( .A(n151), .Z(n154) );
  BUF_X1 U19 ( .A(n166), .Z(n171) );
  BUF_X1 U20 ( .A(n165), .Z(n168) );
  BUF_X1 U21 ( .A(n152), .Z(n156) );
  BUF_X1 U22 ( .A(n166), .Z(n170) );
  BUF_X1 U23 ( .A(n303), .Z(n158) );
  NOR4_X1 U24 ( .A1(n150), .A2(n144), .A3(n153), .A4(n167), .ZN(n303) );
  BUF_X1 U25 ( .A(n301), .Z(n147) );
  BUF_X1 U26 ( .A(n301), .Z(n145) );
  BUF_X1 U27 ( .A(n301), .Z(n148) );
  BUF_X1 U28 ( .A(n301), .Z(n146) );
  BUF_X1 U29 ( .A(n304), .Z(n165) );
  BUF_X1 U30 ( .A(n302), .Z(n151) );
  BUF_X1 U31 ( .A(n304), .Z(n166) );
  BUF_X1 U32 ( .A(n302), .Z(n152) );
  BUF_X1 U33 ( .A(n301), .Z(n149) );
  BUF_X1 U34 ( .A(n300), .Z(n141) );
  BUF_X1 U35 ( .A(n300), .Z(n143) );
  BUF_X1 U36 ( .A(n300), .Z(n139) );
  BUF_X1 U37 ( .A(n300), .Z(n142) );
  BUF_X1 U38 ( .A(n300), .Z(n140) );
  INV_X1 U39 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U40 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n304) );
  AND3_X1 U41 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U42 ( .A(sel[2]), .ZN(n173) );
  NAND2_X1 U43 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI22_X1 U44 ( .A1(C[54]), .A2(n146), .B1(A[54]), .B2(n140), .ZN(n273) );
  AOI222_X1 U45 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n156), .ZN(n272) );
  NAND2_X1 U46 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  AOI22_X1 U47 ( .A1(C[58]), .A2(n145), .B1(A[58]), .B2(n139), .ZN(n281) );
  AOI222_X1 U48 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n157), .ZN(n280) );
  NAND2_X1 U49 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  AOI22_X1 U50 ( .A1(C[57]), .A2(n145), .B1(A[57]), .B2(n139), .ZN(n279) );
  AOI222_X1 U51 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n157), .ZN(n278) );
  NAND2_X1 U52 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  AOI222_X1 U53 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n156), .ZN(n270) );
  AOI22_X1 U54 ( .A1(C[53]), .A2(n146), .B1(A[53]), .B2(n140), .ZN(n271) );
  NAND2_X1 U55 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  NAND2_X1 U56 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  NAND2_X1 U57 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI22_X1 U58 ( .A1(C[52]), .A2(n146), .B1(A[52]), .B2(n140), .ZN(n269) );
  NAND2_X1 U59 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U60 ( .A1(C[63]), .A2(n145), .B1(A[63]), .B2(n139), .ZN(n293) );
  AOI222_X1 U61 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n157), .ZN(n292) );
  AOI222_X1 U62 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n154), .ZN(n214) );
  AOI222_X1 U63 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n154), .ZN(n216) );
  NAND2_X1 U64 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  AOI22_X1 U65 ( .A1(C[30]), .A2(n148), .B1(A[30]), .B2(n142), .ZN(n221) );
  NAND2_X1 U66 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI22_X1 U67 ( .A1(C[33]), .A2(n148), .B1(A[33]), .B2(n142), .ZN(n227) );
  NAND2_X1 U68 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI22_X1 U69 ( .A1(C[31]), .A2(n148), .B1(A[31]), .B2(n142), .ZN(n223) );
  NAND2_X1 U70 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  NAND2_X1 U71 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI22_X1 U72 ( .A1(C[34]), .A2(n148), .B1(A[34]), .B2(n142), .ZN(n229) );
  AOI222_X1 U73 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n155), .ZN(n228) );
  NAND2_X1 U74 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI22_X1 U75 ( .A1(C[38]), .A2(n147), .B1(A[38]), .B2(n141), .ZN(n237) );
  AOI222_X1 U76 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n155), .ZN(n236) );
  NAND2_X1 U77 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI222_X1 U78 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n155), .ZN(n246) );
  AOI22_X1 U79 ( .A1(C[42]), .A2(n147), .B1(A[42]), .B2(n141), .ZN(n247) );
  NAND2_X1 U80 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI22_X1 U81 ( .A1(C[50]), .A2(n146), .B1(A[50]), .B2(n140), .ZN(n265) );
  AOI222_X1 U82 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n156), .ZN(n264) );
  AOI22_X1 U83 ( .A1(C[35]), .A2(n148), .B1(A[35]), .B2(n142), .ZN(n231) );
  AOI222_X1 U84 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n155), .ZN(n230) );
  NAND2_X1 U85 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI22_X1 U86 ( .A1(C[39]), .A2(n147), .B1(A[39]), .B2(n141), .ZN(n239) );
  NAND2_X1 U87 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI222_X1 U88 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n155), .ZN(n248) );
  AOI22_X1 U89 ( .A1(C[43]), .A2(n147), .B1(A[43]), .B2(n141), .ZN(n249) );
  NAND2_X1 U90 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  AOI22_X1 U91 ( .A1(C[32]), .A2(n148), .B1(A[32]), .B2(n142), .ZN(n225) );
  AOI222_X1 U92 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n155), .ZN(n224) );
  NAND2_X1 U93 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  AOI22_X1 U94 ( .A1(C[36]), .A2(n147), .B1(A[36]), .B2(n141), .ZN(n233) );
  AOI222_X1 U95 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n155), .ZN(n232) );
  NAND2_X1 U96 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI22_X1 U97 ( .A1(C[37]), .A2(n147), .B1(A[37]), .B2(n141), .ZN(n235) );
  AOI222_X1 U98 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n155), .ZN(n234) );
  NAND2_X1 U99 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  AOI22_X1 U100 ( .A1(C[40]), .A2(n147), .B1(A[40]), .B2(n141), .ZN(n243) );
  AOI222_X1 U101 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n155), .ZN(n242) );
  NAND2_X1 U102 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI222_X1 U103 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n155), .ZN(n244) );
  AOI22_X1 U104 ( .A1(C[41]), .A2(n147), .B1(A[41]), .B2(n141), .ZN(n245) );
  NAND2_X1 U105 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  AOI22_X1 U106 ( .A1(C[44]), .A2(n147), .B1(A[44]), .B2(n141), .ZN(n251) );
  AOI222_X1 U107 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n156), .ZN(n250) );
  NAND2_X1 U108 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  AOI22_X1 U109 ( .A1(C[61]), .A2(n145), .B1(A[61]), .B2(n139), .ZN(n289) );
  AOI222_X1 U110 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n157), .ZN(n288) );
  NAND2_X1 U111 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI22_X1 U112 ( .A1(C[62]), .A2(n145), .B1(A[62]), .B2(n139), .ZN(n291) );
  AOI222_X1 U113 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n157), .ZN(n290) );
  AOI22_X1 U114 ( .A1(C[48]), .A2(n146), .B1(A[48]), .B2(n140), .ZN(n259) );
  AOI222_X1 U115 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n156), .ZN(n258) );
  NAND2_X1 U116 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI222_X1 U117 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n156), .ZN(n260) );
  AOI22_X1 U118 ( .A1(C[49]), .A2(n146), .B1(A[49]), .B2(n140), .ZN(n261) );
  NAND2_X1 U119 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI222_X1 U120 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n156), .ZN(n254) );
  AOI22_X1 U121 ( .A1(C[46]), .A2(n146), .B1(A[46]), .B2(n140), .ZN(n255) );
  AOI222_X1 U122 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n157), .ZN(n286) );
  AOI22_X1 U123 ( .A1(C[60]), .A2(n145), .B1(A[60]), .B2(n139), .ZN(n287) );
  NAND2_X1 U124 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI222_X1 U125 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n156), .ZN(n256) );
  AOI22_X1 U126 ( .A1(C[47]), .A2(n146), .B1(A[47]), .B2(n140), .ZN(n257) );
  NAND2_X1 U127 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI222_X1 U128 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n156), .ZN(n252) );
  AOI22_X1 U129 ( .A1(C[45]), .A2(n147), .B1(A[45]), .B2(n141), .ZN(n253) );
  NAND2_X1 U130 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U131 ( .A1(C[0]), .A2(n145), .B1(A[0]), .B2(n139), .ZN(n175) );
  AOI222_X1 U132 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n153), .ZN(n174) );
  NAND2_X1 U133 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U134 ( .A1(C[1]), .A2(n149), .B1(A[1]), .B2(n143), .ZN(n197) );
  AOI222_X1 U135 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n153), .ZN(n196) );
  NAND2_X1 U136 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U137 ( .A1(C[4]), .A2(n146), .B1(A[4]), .B2(n140), .ZN(n263) );
  AOI222_X1 U138 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n156), .ZN(n262) );
  NAND2_X1 U139 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U140 ( .A1(C[5]), .A2(n145), .B1(A[5]), .B2(n139), .ZN(n285) );
  AOI222_X1 U141 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n157), .ZN(n284) );
  NAND2_X1 U142 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI22_X1 U143 ( .A1(C[8]), .A2(n145), .B1(A[8]), .B2(n139), .ZN(n299) );
  AOI222_X1 U144 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n157), .ZN(n298) );
  NAND2_X1 U145 ( .A1(n306), .A2(n305), .ZN(Y[9]) );
  AOI22_X1 U146 ( .A1(C[9]), .A2(n147), .B1(A[9]), .B2(n141), .ZN(n306) );
  AOI222_X1 U147 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n157), .ZN(n305) );
  NAND2_X1 U148 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  AOI22_X1 U149 ( .A1(C[12]), .A2(n150), .B1(A[12]), .B2(n144), .ZN(n181) );
  AOI222_X1 U150 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n153), .ZN(n180) );
  NAND2_X1 U151 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U152 ( .A1(C[13]), .A2(n150), .B1(A[13]), .B2(n144), .ZN(n183) );
  AOI222_X1 U153 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n153), .ZN(n182) );
  NAND2_X1 U154 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  AOI22_X1 U155 ( .A1(C[16]), .A2(n149), .B1(A[16]), .B2(n143), .ZN(n189) );
  AOI222_X1 U156 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n153), .ZN(n188) );
  NAND2_X1 U157 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI22_X1 U158 ( .A1(C[17]), .A2(n149), .B1(A[17]), .B2(n143), .ZN(n191) );
  AOI222_X1 U159 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n153), .ZN(n190) );
  NAND2_X1 U160 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  AOI22_X1 U161 ( .A1(C[20]), .A2(n149), .B1(A[20]), .B2(n143), .ZN(n199) );
  AOI222_X1 U162 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n154), .ZN(n198) );
  NAND2_X1 U163 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI22_X1 U164 ( .A1(C[21]), .A2(n149), .B1(A[21]), .B2(n143), .ZN(n201) );
  AOI222_X1 U165 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n154), .ZN(n200) );
  NAND2_X1 U166 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  AOI22_X1 U167 ( .A1(C[24]), .A2(n149), .B1(A[24]), .B2(n143), .ZN(n207) );
  AOI222_X1 U168 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n154), .ZN(n206) );
  NAND2_X1 U169 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI22_X1 U170 ( .A1(C[25]), .A2(n148), .B1(A[25]), .B2(n142), .ZN(n209) );
  AOI222_X1 U171 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n154), .ZN(n208) );
  NAND2_X1 U172 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U173 ( .A1(C[2]), .A2(n148), .B1(A[2]), .B2(n142), .ZN(n219) );
  AOI222_X1 U174 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n154), .ZN(n218) );
  NAND2_X1 U175 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U176 ( .A1(C[6]), .A2(n145), .B1(A[6]), .B2(n139), .ZN(n295) );
  AOI222_X1 U177 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n157), .ZN(n294) );
  NAND2_X1 U178 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U179 ( .A1(C[10]), .A2(n150), .B1(A[10]), .B2(n144), .ZN(n177) );
  AOI222_X1 U180 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n153), .ZN(n176) );
  NAND2_X1 U181 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U182 ( .A1(C[14]), .A2(n149), .B1(A[14]), .B2(n143), .ZN(n185) );
  AOI222_X1 U183 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n153), .ZN(n184) );
  NAND2_X1 U184 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI22_X1 U185 ( .A1(C[18]), .A2(n149), .B1(A[18]), .B2(n143), .ZN(n193) );
  AOI222_X1 U186 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n153), .ZN(n192) );
  NAND2_X1 U187 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI22_X1 U188 ( .A1(C[22]), .A2(n149), .B1(A[22]), .B2(n143), .ZN(n203) );
  AOI222_X1 U189 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n154), .ZN(n202) );
  NAND2_X1 U190 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI22_X1 U191 ( .A1(C[26]), .A2(n148), .B1(A[26]), .B2(n142), .ZN(n211) );
  AOI222_X1 U192 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n154), .ZN(n210) );
  NAND2_X1 U193 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U194 ( .A1(C[3]), .A2(n147), .B1(A[3]), .B2(n141), .ZN(n241) );
  AOI222_X1 U195 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n155), .ZN(n240) );
  NAND2_X1 U196 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U197 ( .A1(C[7]), .A2(n145), .B1(A[7]), .B2(n139), .ZN(n297) );
  AOI222_X1 U198 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n157), .ZN(n296) );
  NAND2_X1 U199 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U200 ( .A1(C[11]), .A2(n150), .B1(A[11]), .B2(n144), .ZN(n179) );
  AOI222_X1 U201 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n153), .ZN(n178) );
  NAND2_X1 U202 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U203 ( .A1(C[15]), .A2(n149), .B1(A[15]), .B2(n143), .ZN(n187) );
  AOI222_X1 U204 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n153), .ZN(n186) );
  NAND2_X1 U205 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI22_X1 U206 ( .A1(C[19]), .A2(n149), .B1(A[19]), .B2(n143), .ZN(n195) );
  AOI222_X1 U207 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n153), .ZN(n194) );
  NAND2_X1 U208 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI22_X1 U209 ( .A1(C[23]), .A2(n149), .B1(A[23]), .B2(n143), .ZN(n205) );
  AOI222_X1 U210 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n154), .ZN(n204) );
  NAND2_X1 U211 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI22_X1 U212 ( .A1(C[27]), .A2(n148), .B1(A[27]), .B2(n142), .ZN(n213) );
  AOI222_X1 U213 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n154), .ZN(n212) );
  AOI22_X1 U214 ( .A1(C[56]), .A2(n146), .B1(A[56]), .B2(n140), .ZN(n277) );
  AOI22_X1 U215 ( .A1(C[55]), .A2(n146), .B1(A[55]), .B2(n140), .ZN(n275) );
  AOI222_X1 U216 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n156), .ZN(n274) );
  AOI22_X1 U217 ( .A1(C[28]), .A2(n148), .B1(A[28]), .B2(n142), .ZN(n215) );
  AOI22_X1 U218 ( .A1(C[29]), .A2(n148), .B1(A[29]), .B2(n142), .ZN(n217) );
  AOI222_X1 U219 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n154), .ZN(n220) );
  NAND2_X1 U220 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  NAND2_X1 U221 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI222_X1 U222 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n155), .ZN(n226) );
  AOI22_X1 U223 ( .A1(C[51]), .A2(n146), .B1(A[51]), .B2(n140), .ZN(n267) );
  AOI222_X1 U224 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n157), .ZN(n276) );
  AOI222_X1 U225 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n156), .ZN(n266) );
  AOI222_X1 U226 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n156), .ZN(n268) );
  AOI22_X1 U227 ( .A1(C[59]), .A2(n145), .B1(A[59]), .B2(n139), .ZN(n283) );
  AOI222_X1 U228 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n157), .ZN(n282) );
  AOI222_X1 U229 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n154), .ZN(n222) );
  CLKBUF_X1 U230 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U231 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U232 ( .A(n158), .Z(n164) );
endmodule


module G_34 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_126 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_125 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_124 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_123 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_122 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_121 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_120 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_119 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_118 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_117 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_116 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_115 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_114 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_113 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_112 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_111 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_110 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_109 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_108 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_107 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_106 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_105 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_104 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_103 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_102 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_101 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_100 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_99 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_98 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_97 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_96 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_33 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_95 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_94 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_93 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_92 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_91 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_90 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_89 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_88 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_87 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_86 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_85 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_84 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_83 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_82 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_81 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_32 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_80 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_79 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_78 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_77 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_76 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_75 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_74 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_31 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_30 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_73 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_72 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_71 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  OR2_X2 U2 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U3 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module PG_70 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_69 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_68 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_29 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_28 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_27 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_26 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_67 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_66 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_65 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_64 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module G_25 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_24 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_23 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_22 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_21 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_20 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_19 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_18 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module carry_generator_N64_NPB4_2 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   n26, \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n11, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U79 ( .A(B[57]), .B(A[57]), .Z(\PG_Network[0][0][57] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U88 ( .A(B[49]), .B(A[49]), .Z(\PG_Network[0][0][49] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U91 ( .A(B[46]), .B(A[46]), .Z(\PG_Network[0][0][46] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U100 ( .A(B[38]), .B(A[38]), .Z(\PG_Network[0][0][38] ) );
  XOR2_X1 U101 ( .A(B[37]), .B(A[37]), .Z(\PG_Network[0][0][37] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U108 ( .A(B[30]), .B(A[30]), .Z(\PG_Network[0][0][30] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U110 ( .A(B[29]), .B(A[29]), .Z(\PG_Network[0][0][29] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U112 ( .A(B[27]), .B(A[27]), .Z(\PG_Network[0][0][27] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U114 ( .A(B[25]), .B(A[25]), .Z(\PG_Network[0][0][25] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U116 ( .A(B[23]), .B(A[23]), .Z(\PG_Network[0][0][23] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U121 ( .A(B[19]), .B(A[19]), .Z(\PG_Network[0][0][19] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U125 ( .A(B[15]), .B(A[15]), .Z(\PG_Network[0][0][15] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_34 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n22), .Gx(\PG_Network[1][1][1] ) );
  PG_126 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_125 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_124 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_123 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_122 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_121 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_120 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_119 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_118 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_117 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_116 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_115 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_114 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_113 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_112 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_111 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_110 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_109 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_108 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_107 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_106 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_105 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_104 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_103 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_102 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_101 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_100 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_99 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_98 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_97 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_96 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_33 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_95 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), 
        .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_94 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_93 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_92 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_91 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_90 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_89 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_88 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_87 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_86 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_85 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_84 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_83 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_82 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_81 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_32 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_80 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_79 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_78 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_77 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_76 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_75 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_74 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(\PG_Network[2][1][59] ), .P_K_1(
        \PG_Network[2][0][59] ), .Gx(\PG_Network[3][1][63] ), .Px(
        \PG_Network[3][0][63] ) );
  G_31 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), 
        .G_K_1(Co[1]), .Gx(Co[3]) );
  G_30 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), 
        .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_73 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_72 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(
        \PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][27] ), .Px(
        \PG_Network[4][0][27] ) );
  PG_71 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(
        \PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(
        \PG_Network[3][0][39] ), .Gx(\PG_Network[4][1][47] ), .Px(
        \PG_Network[4][0][47] ) );
  PG_70 PGJ_3_2_1 ( .G_IK(n9), .P_IK(\PG_Network[2][0][43] ), .G_K_1(
        \PG_Network[3][1][39] ), .P_K_1(\PG_Network[3][0][39] ), .Gx(
        \PG_Network[4][1][43] ), .Px(\PG_Network[4][0][43] ) );
  PG_69 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(
        \PG_Network[3][0][63] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][63] ), .Px(
        \PG_Network[4][0][63] ) );
  PG_68 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(
        \PG_Network[2][0][59] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(
        \PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][59] ), .Px(
        \PG_Network[4][0][59] ) );
  G_29 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), 
        .G_K_1(Co[3]), .Gx(n26) );
  G_28 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), 
        .G_K_1(Co[3]), .Gx(Co[6]) );
  G_27 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), 
        .G_K_1(Co[3]), .Gx(Co[5]) );
  G_26 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), 
        .G_K_1(Co[3]), .Gx(Co[4]) );
  PG_67 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(
        \PG_Network[4][0][63] ), .G_K_1(n17), .P_K_1(n12), .Gx(
        \PG_Network[5][1][63] ), .Px(\PG_Network[5][0][63] ) );
  PG_66 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(
        \PG_Network[4][0][59] ), .G_K_1(n17), .P_K_1(n12), .Gx(
        \PG_Network[5][1][59] ), .Px(\PG_Network[5][0][59] ) );
  PG_65 PGJ_4_1_2 ( .G_IK(\PG_Network[3][1][55] ), .P_IK(
        \PG_Network[3][0][55] ), .G_K_1(n17), .P_K_1(n12), .Gx(
        \PG_Network[5][1][55] ), .Px(\PG_Network[5][0][55] ) );
  PG_64 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(
        \PG_Network[2][0][51] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(
        \PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][51] ), .Px(
        \PG_Network[5][0][51] ) );
  G_25 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), 
        .G_K_1(Co[7]), .Gx(Co[15]) );
  G_24 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), 
        .G_K_1(Co[7]), .Gx(Co[14]) );
  G_23 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), 
        .G_K_1(Co[7]), .Gx(Co[13]) );
  G_22 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), 
        .G_K_1(Co[7]), .Gx(Co[12]) );
  G_21 GJ_5_0_4 ( .G_IK(\PG_Network[4][1][47] ), .P_IK(\PG_Network[4][0][47] ), 
        .G_K_1(n26), .Gx(Co[11]) );
  G_20 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), 
        .G_K_1(n26), .Gx(Co[10]) );
  G_19 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), 
        .G_K_1(n26), .Gx(Co[9]) );
  G_18 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), 
        .G_K_1(n26), .Gx(Co[8]) );
  BUF_X2 U1 ( .A(n26), .Z(Co[7]) );
  NAND2_X1 U2 ( .A1(B[35]), .A2(n6), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n5), .A2(A[35]), .ZN(n8) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(\PG_Network[0][0][35] ) );
  INV_X1 U5 ( .A(B[35]), .ZN(n5) );
  INV_X1 U6 ( .A(A[35]), .ZN(n6) );
  CLKBUF_X1 U7 ( .A(\PG_Network[2][1][43] ), .Z(n9) );
  INV_X1 U8 ( .A(A[31]), .ZN(n15) );
  INV_X1 U9 ( .A(A[43]), .ZN(n14) );
  INV_X1 U10 ( .A(A[45]), .ZN(n11) );
  INV_X1 U11 ( .A(A[53]), .ZN(n10) );
  INV_X1 U12 ( .A(A[59]), .ZN(n21) );
  INV_X1 U13 ( .A(A[55]), .ZN(n18) );
  INV_X1 U14 ( .A(A[39]), .ZN(n16) );
  INV_X1 U15 ( .A(A[47]), .ZN(n20) );
  INV_X1 U16 ( .A(A[51]), .ZN(n19) );
  XNOR2_X1 U17 ( .A(B[53]), .B(n10), .ZN(\PG_Network[0][0][53] ) );
  XNOR2_X1 U18 ( .A(B[45]), .B(n11), .ZN(\PG_Network[0][0][45] ) );
  CLKBUF_X1 U19 ( .A(\PG_Network[4][1][47] ), .Z(n17) );
  CLKBUF_X1 U20 ( .A(\PG_Network[4][0][47] ), .Z(n12) );
  XNOR2_X1 U21 ( .A(B[43]), .B(n14), .ZN(\PG_Network[0][0][43] ) );
  XNOR2_X1 U22 ( .A(B[31]), .B(n15), .ZN(\PG_Network[0][0][31] ) );
  XNOR2_X1 U23 ( .A(B[39]), .B(n16), .ZN(\PG_Network[0][0][39] ) );
  XNOR2_X1 U24 ( .A(B[55]), .B(n18), .ZN(\PG_Network[0][0][55] ) );
  XNOR2_X1 U25 ( .A(B[51]), .B(n19), .ZN(\PG_Network[0][0][51] ) );
  XNOR2_X1 U26 ( .A(B[47]), .B(n20), .ZN(\PG_Network[0][0][47] ) );
  XNOR2_X1 U27 ( .A(B[59]), .B(n21), .ZN(\PG_Network[0][0][59] ) );
  AND2_X1 U28 ( .A1(B[50]), .A2(A[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U29 ( .A1(B[51]), .A2(A[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U30 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U31 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U32 ( .A1(A[46]), .A2(B[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U33 ( .A1(A[57]), .A2(B[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U34 ( .A1(A[37]), .A2(B[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U35 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U36 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U37 ( .A1(B[31]), .A2(A[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U38 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U39 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U40 ( .A1(B[35]), .A2(A[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U41 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U42 ( .A1(A[41]), .A2(B[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U43 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U44 ( .A1(B[49]), .A2(A[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U45 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U46 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U47 ( .A1(A[43]), .A2(B[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U48 ( .A1(B[39]), .A2(A[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U49 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U50 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U51 ( .A1(A[29]), .A2(B[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U52 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U53 ( .A1(B[52]), .A2(A[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U54 ( .A1(B[53]), .A2(A[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U55 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U56 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U57 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U58 ( .A1(A[19]), .A2(B[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U59 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U60 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U61 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U62 ( .A1(A[11]), .A2(B[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U63 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U64 ( .A1(A[15]), .A2(B[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U65 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U66 ( .A1(A[25]), .A2(B[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U67 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U77 ( .A1(A[27]), .A2(B[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U81 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U83 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U85 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U90 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U92 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U94 ( .A(n25), .ZN(n22) );
  AND2_X1 U99 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U103 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U107 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U131 ( .A1(A[7]), .A2(B[7]), .ZN(\PG_Network[0][1][7] ) );
  AND2_X1 U132 ( .A1(A[21]), .A2(B[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U133 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U134 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U135 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AND2_X1 U136 ( .A1(A[23]), .A2(B[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U137 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AOI21_X1 U138 ( .B1(A[0]), .B2(B[0]), .A(n23), .ZN(n25) );
  INV_X1 U139 ( .A(n24), .ZN(n23) );
  OAI21_X1 U140 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n24) );
  AND2_X1 U141 ( .A1(B[55]), .A2(A[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U142 ( .A1(B[47]), .A2(A[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U143 ( .A1(A[45]), .A2(B[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U144 ( .A1(B[59]), .A2(A[59]), .ZN(\PG_Network[0][1][59] ) );
  AND2_X1 U145 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U146 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U147 ( .A1(A[56]), .A2(B[56]), .ZN(\PG_Network[0][1][56] ) );
endmodule


module FA_256 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_64 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_256 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_255 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_254 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_253 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_252 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_251 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_250 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_249 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_63 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_252 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_251 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_250 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_249 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_32 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U2 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U4 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U5 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U7 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_32 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_64 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_63 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_32 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_62 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_248 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_247 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_246 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_245 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_244 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_243 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_242 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_241 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_61 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_244 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_243 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_242 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_241 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_31 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_31 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_62 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_61 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_31 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_60 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_240 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_239 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_238 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_237 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_236 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_235 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_234 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_233 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_59 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_236 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_235 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_234 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_233 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_30 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_30 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_60 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_59 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_30 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_58 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_232 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_231 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_230 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_229 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_228 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_227 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_226 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_225 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_57 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_228 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_227 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_226 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_225 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_29 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_29 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_58 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_57 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_29 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_56 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_224 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_223 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_222 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_221 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_220 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_219 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_218 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_217 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_55 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_220 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_219 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_218 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_217 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_28 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_28 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_56 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_55 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_28 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_216 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_215 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_214 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_213 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_54 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_216 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_215 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_214 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_213 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_212 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_211 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_210 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_209 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_53 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_212 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_211 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_210 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_209 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_27 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_27 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_54 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_53 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_27 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_208 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_207 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_206 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_205 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_52 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_208 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_207 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_206 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_205 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_204 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_203 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_202 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_201 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_51 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_204 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_203 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_202 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_201 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_26 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_26 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_52 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_51 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_26 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_200 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_50 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_200 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_199 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_198 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_197 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_196 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_195 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_194 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_193 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_49 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_196 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_195 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_194 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_193 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_25 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_25 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_50 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_49 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_25 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_192 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_191 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_190 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_189 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_48 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_192 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_191 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_190 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_189 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_188 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_187 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_186 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_185 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_47 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_188 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_187 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_186 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_185 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_24 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_24 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_48 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_47 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_24 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_184 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_183 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_182 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_181 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_46 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_184 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_183 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_182 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_181 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_180 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_179 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_178 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_177 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_45 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_180 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_179 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_178 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_177 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_23 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X2 U1 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(sel), .ZN(n13) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_23 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_46 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_45 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_23 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_176 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n5) );
  INV_X1 U5 ( .A(n8), .ZN(Co) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
endmodule


module FA_175 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_174 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_173 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_44 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_176 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_175 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_174 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_173 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_172 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_171 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_170 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_169 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_43 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_172 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_171 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_170 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_169 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_22 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_22 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_44 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_43 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_22 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_168 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_167 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_166 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_165 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_42 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_168 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_167 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_166 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_165 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_164 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_163 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_162 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_161 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_41 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_164 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_163 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_162 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_161 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_21 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U2 ( .A(sel), .ZN(n13) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U5 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U6 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U7 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n13), .ZN(n17) );
endmodule


module carry_select_block_NPB4_21 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_42 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_41 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_21 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_160 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n4), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_159 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_158 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_157 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_40 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_160 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_159 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_158 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_157 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_156 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_155 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_154 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_153 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_39 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_156 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_155 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_154 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_153 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_20 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(sel), .ZN(n5) );
  INV_X1 U2 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U3 ( .A(sel), .ZN(n14) );
  INV_X1 U4 ( .A(n17), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n5), .ZN(n17) );
  INV_X1 U6 ( .A(n16), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  INV_X1 U8 ( .A(n15), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n14), .ZN(n15) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n14), .ZN(n18) );
endmodule


module carry_select_block_NPB4_20 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_40 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_39 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_20 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net67776, n4, n5, n6, n7;
  assign Co = net67776;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n7) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n5) );
  INV_X1 U5 ( .A(n5), .ZN(net67776) );
  XNOR2_X1 U6 ( .A(B), .B(n7), .ZN(n6) );
endmodule


module FA_151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net67775, n4, n5, n6;
  assign Co = net67775;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n5) );
  INV_X1 U5 ( .A(n5), .ZN(net67775) );
endmodule


module FA_150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  OR2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n7) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(n4), .ZN(n10) );
endmodule


module RCA_N4_38 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_152 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_151 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_150 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_149 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_148 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_147 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_146 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_145 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_37 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_148 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_147 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_146 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_145 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_19 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U2 ( .A(sel), .ZN(n5) );
  INV_X1 U3 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U5 ( .A(n15), .ZN(Y[0]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[2]), .B1(B[2]), .B2(n5), .ZN(n17) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[0]), .B1(B[0]), .B2(n5), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(sel), .B1(n14), .B2(B[3]), .ZN(n18) );
  AOI22_X1 U9 ( .A1(sel), .A2(A[1]), .B1(n14), .B2(B[1]), .ZN(n16) );
  INV_X1 U10 ( .A(sel), .ZN(n14) );
endmodule


module carry_select_block_NPB4_19 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_38 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_37 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_19 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n5) );
  INV_X1 U4 ( .A(A), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  AOI22_X1 U6 ( .A1(n4), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  INV_X1 U7 ( .A(n9), .ZN(Co) );
endmodule


module FA_143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n4) );
  OR2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n7) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(n4), .ZN(n10) );
endmodule


module RCA_N4_36 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_144 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_143 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_142 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_141 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_140 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_139 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  INV_X1 U1 ( .A(B), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(n5) );
  XOR2_X1 U5 ( .A(A), .B(n5), .Z(n6) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n5), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_138 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_137 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(n9), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_35 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_140 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_139 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_138 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_137 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_18 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(sel), .ZN(n5) );
  INV_X1 U2 ( .A(n16), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n17), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[0]), .B1(n14), .B2(B[0]), .ZN(n15) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[2]), .B1(n14), .B2(B[2]), .ZN(n17) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[1]), .B1(B[1]), .B2(n5), .ZN(n16) );
  INV_X1 U9 ( .A(sel), .ZN(n14) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n14), .ZN(n18) );
endmodule


module carry_select_block_NPB4_18 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_36 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_35 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_18 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  CLKBUF_X1 U1 ( .A(B), .Z(n4) );
  INV_X1 U2 ( .A(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(n5), .B(B), .ZN(n8) );
  XOR2_X1 U5 ( .A(A), .B(n4), .Z(n6) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n4), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
endmodule


module FA_135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n4), .B2(Ci), .ZN(n7) );
endmodule


module RCA_N4_34 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_136 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_135 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_134 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_133 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_132 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_131 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(n4), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_130 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(n4), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_129 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n7, n9, n10;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n4) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n5), .A2(n9), .ZN(n7) );
  NAND2_X1 U5 ( .A1(n6), .A2(n7), .ZN(S) );
  INV_X1 U6 ( .A(Ci), .ZN(n5) );
  INV_X1 U7 ( .A(n10), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
endmodule


module RCA_N4_33 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_132 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_131 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_130 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_129 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_17 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n10, n15, n16, n17, n18, n19;

  INV_X2 U1 ( .A(n16), .ZN(Y[0]) );
  INV_X1 U2 ( .A(sel), .ZN(n5) );
  INV_X1 U3 ( .A(n5), .ZN(n10) );
  INV_X1 U4 ( .A(n18), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[1]) );
  INV_X1 U6 ( .A(n19), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n10), .B1(B[2]), .B2(n5), .ZN(n18) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n5), .ZN(n17) );
  INV_X1 U9 ( .A(sel), .ZN(n15) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(n10), .B1(B[3]), .B2(n5), .ZN(n19) );
  AOI22_X1 U11 ( .A1(sel), .A2(A[0]), .B1(n15), .B2(B[0]), .ZN(n16) );
endmodule


module carry_select_block_NPB4_17 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_34 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_33 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_17 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_2 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_32 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_31 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_30 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_29 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_28 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_27 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_26 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_25 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_24 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_23 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_22 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), 
        .S(S[43:40]) );
  carry_select_block_NPB4_21 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), 
        .S(S[47:44]) );
  carry_select_block_NPB4_20 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), 
        .S(S[51:48]) );
  carry_select_block_NPB4_19 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), 
        .S(S[55:52]) );
  carry_select_block_NPB4_18 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), 
        .S(S[59:56]) );
  carry_select_block_NPB4_17 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), 
        .S(S[63:60]) );
endmodule


module P4_ADDER_N64_2 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_2 CGEN ( .A(A), .B({n1, B[62:61], n17, B[59:57], n3, 
        B[55:53], n16, B[51:49], n8, B[47:0]}), .Cin(Cin), .Co(CoutCgen) );
  sum_generator_N64_NPB4_2 SGEN ( .A(A), .B({B[63:60], n15, n13, B[57:56], n14, 
        n5, B[53:52], n6, n2, B[49:48], n7, B[46:44], n10, B[42:40], n11, 
        B[38:36], n4, B[34:0]}), .Ci({CoutCgen, Cin}), .S(S), .Co(Cout) );
  CLKBUF_X1 U1 ( .A(B[63]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(B[50]), .Z(n2) );
  CLKBUF_X1 U3 ( .A(B[56]), .Z(n3) );
  CLKBUF_X1 U4 ( .A(B[35]), .Z(n4) );
  BUF_X1 U5 ( .A(B[52]), .Z(n16) );
  BUF_X1 U6 ( .A(B[48]), .Z(n8) );
  BUF_X1 U7 ( .A(B[54]), .Z(n5) );
  CLKBUF_X1 U8 ( .A(B[51]), .Z(n6) );
  CLKBUF_X1 U9 ( .A(B[47]), .Z(n7) );
  INV_X1 U10 ( .A(B[43]), .ZN(n9) );
  INV_X1 U11 ( .A(n9), .ZN(n10) );
  CLKBUF_X1 U12 ( .A(B[39]), .Z(n11) );
  INV_X1 U13 ( .A(B[58]), .ZN(n12) );
  INV_X1 U14 ( .A(n12), .ZN(n13) );
  CLKBUF_X1 U15 ( .A(B[55]), .Z(n14) );
  CLKBUF_X1 U16 ( .A(B[59]), .Z(n15) );
  CLKBUF_X1 U17 ( .A(B[60]), .Z(n17) );
endmodule


module Booth_Encoder_1 ( i, o );
  input [2:0] i;
  output [2:0] o;
  wire   n4, n6, n7;

  OAI22_X1 U3 ( .A1(n4), .A2(n6), .B1(i[2]), .B2(n7), .ZN(o[1]) );
  INV_X1 U4 ( .A(i[2]), .ZN(n4) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(i[2]), .ZN(o[0]) );
  OAI21_X1 U6 ( .B1(i[1]), .B2(i[0]), .A(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(i[1]), .A2(i[0]), .ZN(n7) );
  AND3_X1 U8 ( .A1(i[2]), .A2(n7), .A3(n6), .ZN(o[2]) );
endmodule


module MUX_booth_N64_1 ( A, B, C, D, E, sel, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] sel;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306;

  NOR3_X1 U1 ( .A1(sel[0]), .A2(sel[2]), .A3(n172), .ZN(n301) );
  NOR3_X1 U2 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n300) );
  AOI222_X1 U3 ( .A1(D[41]), .A2(n169), .B1(E[41]), .B2(n161), .C1(B[41]), 
        .C2(n155), .ZN(n244) );
  BUF_X1 U4 ( .A(n158), .Z(n162) );
  BUF_X1 U5 ( .A(n158), .Z(n161) );
  BUF_X1 U6 ( .A(n158), .Z(n163) );
  BUF_X1 U7 ( .A(n158), .Z(n159) );
  BUF_X1 U8 ( .A(n158), .Z(n160) );
  BUF_X1 U9 ( .A(n151), .Z(n153) );
  BUF_X1 U10 ( .A(n165), .Z(n167) );
  BUF_X1 U11 ( .A(n303), .Z(n158) );
  NOR4_X1 U12 ( .A1(n150), .A2(n144), .A3(n153), .A4(n167), .ZN(n303) );
  BUF_X1 U13 ( .A(n151), .Z(n154) );
  BUF_X1 U14 ( .A(n165), .Z(n168) );
  BUF_X1 U15 ( .A(n152), .Z(n156) );
  BUF_X1 U16 ( .A(n166), .Z(n170) );
  BUF_X1 U17 ( .A(n151), .Z(n155) );
  BUF_X1 U18 ( .A(n152), .Z(n157) );
  BUF_X1 U19 ( .A(n165), .Z(n169) );
  BUF_X1 U20 ( .A(n166), .Z(n171) );
  BUF_X1 U21 ( .A(n304), .Z(n165) );
  BUF_X1 U22 ( .A(n302), .Z(n151) );
  BUF_X1 U23 ( .A(n301), .Z(n147) );
  BUF_X1 U24 ( .A(n301), .Z(n146) );
  BUF_X1 U25 ( .A(n301), .Z(n148) );
  BUF_X1 U26 ( .A(n301), .Z(n145) );
  BUF_X1 U27 ( .A(n304), .Z(n166) );
  BUF_X1 U28 ( .A(n302), .Z(n152) );
  BUF_X1 U29 ( .A(n301), .Z(n149) );
  BUF_X1 U30 ( .A(n300), .Z(n143) );
  BUF_X1 U31 ( .A(n300), .Z(n141) );
  BUF_X1 U32 ( .A(n300), .Z(n140) );
  BUF_X1 U33 ( .A(n300), .Z(n142) );
  BUF_X1 U34 ( .A(n300), .Z(n139) );
  INV_X1 U35 ( .A(sel[1]), .ZN(n172) );
  AND3_X1 U36 ( .A1(sel[0]), .A2(n173), .A3(sel[1]), .ZN(n304) );
  AND3_X1 U37 ( .A1(n172), .A2(n173), .A3(sel[0]), .ZN(n302) );
  INV_X1 U38 ( .A(sel[2]), .ZN(n173) );
  NAND2_X1 U39 ( .A1(n225), .A2(n224), .ZN(Y[32]) );
  AOI22_X1 U40 ( .A1(C[32]), .A2(n148), .B1(A[32]), .B2(n142), .ZN(n225) );
  NAND2_X1 U41 ( .A1(n271), .A2(n270), .ZN(Y[53]) );
  NAND2_X1 U42 ( .A1(n273), .A2(n272), .ZN(Y[54]) );
  AOI22_X1 U43 ( .A1(C[54]), .A2(n146), .B1(A[54]), .B2(n140), .ZN(n273) );
  NAND2_X1 U44 ( .A1(n279), .A2(n278), .ZN(Y[57]) );
  NAND2_X1 U45 ( .A1(n281), .A2(n280), .ZN(Y[58]) );
  NAND2_X1 U46 ( .A1(n277), .A2(n276), .ZN(Y[56]) );
  AOI22_X1 U47 ( .A1(C[56]), .A2(n146), .B1(A[56]), .B2(n140), .ZN(n277) );
  AOI222_X1 U48 ( .A1(D[56]), .A2(n171), .B1(E[56]), .B2(n163), .C1(B[56]), 
        .C2(n157), .ZN(n276) );
  NAND2_X1 U49 ( .A1(n287), .A2(n286), .ZN(Y[60]) );
  AOI22_X1 U50 ( .A1(C[60]), .A2(n145), .B1(A[60]), .B2(n139), .ZN(n287) );
  AOI222_X1 U51 ( .A1(D[60]), .A2(n171), .B1(E[60]), .B2(n163), .C1(B[60]), 
        .C2(n157), .ZN(n286) );
  NAND2_X1 U52 ( .A1(n293), .A2(n292), .ZN(Y[63]) );
  AOI22_X1 U53 ( .A1(C[63]), .A2(n145), .B1(A[63]), .B2(n139), .ZN(n293) );
  AOI222_X1 U54 ( .A1(D[63]), .A2(n171), .B1(E[63]), .B2(n163), .C1(B[63]), 
        .C2(n157), .ZN(n292) );
  AOI222_X1 U55 ( .A1(D[31]), .A2(n168), .B1(E[31]), .B2(n161), .C1(B[31]), 
        .C2(n154), .ZN(n222) );
  NAND2_X1 U56 ( .A1(n227), .A2(n226), .ZN(Y[33]) );
  AOI22_X1 U57 ( .A1(C[33]), .A2(n148), .B1(A[33]), .B2(n142), .ZN(n227) );
  NAND2_X1 U58 ( .A1(n231), .A2(n230), .ZN(Y[35]) );
  AOI22_X1 U59 ( .A1(C[35]), .A2(n148), .B1(A[35]), .B2(n142), .ZN(n231) );
  NAND2_X1 U60 ( .A1(n233), .A2(n232), .ZN(Y[36]) );
  AOI22_X1 U61 ( .A1(C[36]), .A2(n147), .B1(A[36]), .B2(n141), .ZN(n233) );
  AOI222_X1 U62 ( .A1(D[36]), .A2(n169), .B1(E[36]), .B2(n161), .C1(B[36]), 
        .C2(n155), .ZN(n232) );
  NAND2_X1 U63 ( .A1(n243), .A2(n242), .ZN(Y[40]) );
  AOI22_X1 U64 ( .A1(C[40]), .A2(n147), .B1(A[40]), .B2(n141), .ZN(n243) );
  AOI222_X1 U65 ( .A1(D[40]), .A2(n169), .B1(E[40]), .B2(n161), .C1(B[40]), 
        .C2(n155), .ZN(n242) );
  NAND2_X1 U66 ( .A1(n251), .A2(n250), .ZN(Y[44]) );
  AOI222_X1 U67 ( .A1(D[44]), .A2(n170), .B1(E[44]), .B2(n162), .C1(B[44]), 
        .C2(n156), .ZN(n250) );
  AOI22_X1 U68 ( .A1(C[44]), .A2(n147), .B1(A[44]), .B2(n141), .ZN(n251) );
  NAND2_X1 U69 ( .A1(n269), .A2(n268), .ZN(Y[52]) );
  AOI22_X1 U70 ( .A1(C[52]), .A2(n146), .B1(A[52]), .B2(n140), .ZN(n269) );
  AOI222_X1 U71 ( .A1(D[52]), .A2(n170), .B1(E[52]), .B2(n162), .C1(B[52]), 
        .C2(n156), .ZN(n268) );
  NAND2_X1 U72 ( .A1(n265), .A2(n264), .ZN(Y[50]) );
  AOI22_X1 U73 ( .A1(C[50]), .A2(n146), .B1(A[50]), .B2(n140), .ZN(n265) );
  AOI222_X1 U74 ( .A1(D[50]), .A2(n170), .B1(E[50]), .B2(n162), .C1(B[50]), 
        .C2(n156), .ZN(n264) );
  NAND2_X1 U75 ( .A1(n235), .A2(n234), .ZN(Y[37]) );
  AOI22_X1 U76 ( .A1(C[37]), .A2(n147), .B1(A[37]), .B2(n141), .ZN(n235) );
  AOI222_X1 U77 ( .A1(D[37]), .A2(n169), .B1(E[37]), .B2(n161), .C1(B[37]), 
        .C2(n155), .ZN(n234) );
  NAND2_X1 U78 ( .A1(n245), .A2(n244), .ZN(Y[41]) );
  AOI22_X1 U79 ( .A1(C[41]), .A2(n147), .B1(A[41]), .B2(n141), .ZN(n245) );
  NAND2_X1 U80 ( .A1(n253), .A2(n252), .ZN(Y[45]) );
  AOI222_X1 U81 ( .A1(D[45]), .A2(n170), .B1(E[45]), .B2(n162), .C1(B[45]), 
        .C2(n156), .ZN(n252) );
  AOI22_X1 U82 ( .A1(C[45]), .A2(n147), .B1(A[45]), .B2(n141), .ZN(n253) );
  NAND2_X1 U83 ( .A1(n261), .A2(n260), .ZN(Y[49]) );
  AOI222_X1 U84 ( .A1(D[49]), .A2(n170), .B1(E[49]), .B2(n162), .C1(B[49]), 
        .C2(n156), .ZN(n260) );
  AOI22_X1 U85 ( .A1(C[49]), .A2(n146), .B1(A[49]), .B2(n140), .ZN(n261) );
  NAND2_X1 U86 ( .A1(n255), .A2(n254), .ZN(Y[46]) );
  AOI22_X1 U87 ( .A1(C[46]), .A2(n146), .B1(A[46]), .B2(n140), .ZN(n255) );
  AOI222_X1 U88 ( .A1(D[46]), .A2(n170), .B1(E[46]), .B2(n162), .C1(B[46]), 
        .C2(n156), .ZN(n254) );
  NAND2_X1 U89 ( .A1(n257), .A2(n256), .ZN(Y[47]) );
  AOI222_X1 U90 ( .A1(D[47]), .A2(n170), .B1(E[47]), .B2(n162), .C1(B[47]), 
        .C2(n156), .ZN(n256) );
  AOI22_X1 U91 ( .A1(C[47]), .A2(n146), .B1(A[47]), .B2(n140), .ZN(n257) );
  NAND2_X1 U92 ( .A1(n275), .A2(n274), .ZN(Y[55]) );
  AOI222_X1 U93 ( .A1(D[55]), .A2(n170), .B1(E[55]), .B2(n163), .C1(B[55]), 
        .C2(n156), .ZN(n274) );
  AOI22_X1 U94 ( .A1(C[55]), .A2(n146), .B1(A[55]), .B2(n140), .ZN(n275) );
  NAND2_X1 U95 ( .A1(n239), .A2(n238), .ZN(Y[39]) );
  AOI22_X1 U96 ( .A1(C[39]), .A2(n147), .B1(A[39]), .B2(n141), .ZN(n239) );
  AOI222_X1 U97 ( .A1(D[39]), .A2(n169), .B1(E[39]), .B2(n161), .C1(B[39]), 
        .C2(n155), .ZN(n238) );
  NAND2_X1 U98 ( .A1(n249), .A2(n248), .ZN(Y[43]) );
  AOI222_X1 U99 ( .A1(D[43]), .A2(n169), .B1(E[43]), .B2(n162), .C1(B[43]), 
        .C2(n155), .ZN(n248) );
  AOI22_X1 U100 ( .A1(C[43]), .A2(n147), .B1(A[43]), .B2(n141), .ZN(n249) );
  NAND2_X1 U101 ( .A1(n229), .A2(n228), .ZN(Y[34]) );
  AOI22_X1 U102 ( .A1(C[34]), .A2(n148), .B1(A[34]), .B2(n142), .ZN(n229) );
  AOI222_X1 U103 ( .A1(D[34]), .A2(n169), .B1(E[34]), .B2(n161), .C1(B[34]), 
        .C2(n155), .ZN(n228) );
  NAND2_X1 U104 ( .A1(n237), .A2(n236), .ZN(Y[38]) );
  AOI22_X1 U105 ( .A1(C[38]), .A2(n147), .B1(A[38]), .B2(n141), .ZN(n237) );
  AOI222_X1 U106 ( .A1(D[38]), .A2(n169), .B1(E[38]), .B2(n161), .C1(B[38]), 
        .C2(n155), .ZN(n236) );
  NAND2_X1 U107 ( .A1(n247), .A2(n246), .ZN(Y[42]) );
  AOI22_X1 U108 ( .A1(C[42]), .A2(n147), .B1(A[42]), .B2(n141), .ZN(n247) );
  AOI222_X1 U109 ( .A1(D[42]), .A2(n169), .B1(E[42]), .B2(n162), .C1(B[42]), 
        .C2(n155), .ZN(n246) );
  NAND2_X1 U110 ( .A1(n291), .A2(n290), .ZN(Y[62]) );
  AOI222_X1 U111 ( .A1(D[62]), .A2(n171), .B1(E[62]), .B2(n163), .C1(B[62]), 
        .C2(n157), .ZN(n290) );
  AOI22_X1 U112 ( .A1(C[62]), .A2(n145), .B1(A[62]), .B2(n139), .ZN(n291) );
  NAND2_X1 U113 ( .A1(n289), .A2(n288), .ZN(Y[61]) );
  NAND2_X1 U114 ( .A1(n259), .A2(n258), .ZN(Y[48]) );
  AOI222_X1 U115 ( .A1(D[48]), .A2(n170), .B1(E[48]), .B2(n162), .C1(B[48]), 
        .C2(n156), .ZN(n258) );
  AOI22_X1 U116 ( .A1(C[48]), .A2(n146), .B1(A[48]), .B2(n140), .ZN(n259) );
  NAND2_X1 U117 ( .A1(n267), .A2(n266), .ZN(Y[51]) );
  AOI222_X1 U118 ( .A1(D[51]), .A2(n170), .B1(E[51]), .B2(n162), .C1(B[51]), 
        .C2(n156), .ZN(n266) );
  AOI22_X1 U119 ( .A1(C[51]), .A2(n146), .B1(A[51]), .B2(n140), .ZN(n267) );
  NAND2_X1 U120 ( .A1(n283), .A2(n282), .ZN(Y[59]) );
  AOI22_X1 U121 ( .A1(C[59]), .A2(n145), .B1(A[59]), .B2(n139), .ZN(n283) );
  AOI222_X1 U122 ( .A1(D[59]), .A2(n171), .B1(E[59]), .B2(n163), .C1(B[59]), 
        .C2(n157), .ZN(n282) );
  AOI222_X1 U123 ( .A1(D[30]), .A2(n168), .B1(E[30]), .B2(n160), .C1(B[30]), 
        .C2(n154), .ZN(n220) );
  NAND2_X1 U124 ( .A1(n175), .A2(n174), .ZN(Y[0]) );
  AOI22_X1 U125 ( .A1(C[0]), .A2(n145), .B1(A[0]), .B2(n139), .ZN(n175) );
  AOI222_X1 U126 ( .A1(D[0]), .A2(n167), .B1(E[0]), .B2(n159), .C1(B[0]), .C2(
        n153), .ZN(n174) );
  NAND2_X1 U127 ( .A1(n197), .A2(n196), .ZN(Y[1]) );
  AOI22_X1 U128 ( .A1(C[1]), .A2(n149), .B1(A[1]), .B2(n143), .ZN(n197) );
  AOI222_X1 U129 ( .A1(D[1]), .A2(n167), .B1(E[1]), .B2(n159), .C1(B[1]), .C2(
        n153), .ZN(n196) );
  NAND2_X1 U130 ( .A1(n219), .A2(n218), .ZN(Y[2]) );
  AOI22_X1 U131 ( .A1(C[2]), .A2(n148), .B1(A[2]), .B2(n142), .ZN(n219) );
  AOI222_X1 U132 ( .A1(D[2]), .A2(n168), .B1(E[2]), .B2(n160), .C1(B[2]), .C2(
        n154), .ZN(n218) );
  NAND2_X1 U133 ( .A1(n263), .A2(n262), .ZN(Y[4]) );
  AOI22_X1 U134 ( .A1(C[4]), .A2(n146), .B1(A[4]), .B2(n140), .ZN(n263) );
  AOI222_X1 U135 ( .A1(D[4]), .A2(n170), .B1(E[4]), .B2(n162), .C1(B[4]), .C2(
        n156), .ZN(n262) );
  NAND2_X1 U136 ( .A1(n285), .A2(n284), .ZN(Y[5]) );
  AOI22_X1 U137 ( .A1(C[5]), .A2(n145), .B1(A[5]), .B2(n139), .ZN(n285) );
  AOI222_X1 U138 ( .A1(D[5]), .A2(n171), .B1(E[5]), .B2(n163), .C1(B[5]), .C2(
        n157), .ZN(n284) );
  NAND2_X1 U139 ( .A1(n295), .A2(n294), .ZN(Y[6]) );
  AOI22_X1 U140 ( .A1(C[6]), .A2(n145), .B1(A[6]), .B2(n139), .ZN(n295) );
  AOI222_X1 U141 ( .A1(D[6]), .A2(n171), .B1(E[6]), .B2(n164), .C1(B[6]), .C2(
        n157), .ZN(n294) );
  NAND2_X1 U142 ( .A1(n299), .A2(n298), .ZN(Y[8]) );
  AOI22_X1 U143 ( .A1(C[8]), .A2(n145), .B1(A[8]), .B2(n139), .ZN(n299) );
  AOI222_X1 U144 ( .A1(D[8]), .A2(n171), .B1(E[8]), .B2(n164), .C1(B[8]), .C2(
        n157), .ZN(n298) );
  NAND2_X1 U145 ( .A1(n306), .A2(n305), .ZN(Y[9]) );
  AOI22_X1 U146 ( .A1(C[9]), .A2(n147), .B1(A[9]), .B2(n141), .ZN(n306) );
  AOI222_X1 U147 ( .A1(D[9]), .A2(n171), .B1(E[9]), .B2(n164), .C1(B[9]), .C2(
        n157), .ZN(n305) );
  NAND2_X1 U148 ( .A1(n177), .A2(n176), .ZN(Y[10]) );
  AOI22_X1 U149 ( .A1(C[10]), .A2(n150), .B1(A[10]), .B2(n144), .ZN(n177) );
  AOI222_X1 U150 ( .A1(D[10]), .A2(n167), .B1(E[10]), .B2(n159), .C1(B[10]), 
        .C2(n153), .ZN(n176) );
  NAND2_X1 U151 ( .A1(n181), .A2(n180), .ZN(Y[12]) );
  AOI22_X1 U152 ( .A1(C[12]), .A2(n150), .B1(A[12]), .B2(n144), .ZN(n181) );
  AOI222_X1 U153 ( .A1(D[12]), .A2(n167), .B1(E[12]), .B2(n159), .C1(B[12]), 
        .C2(n153), .ZN(n180) );
  NAND2_X1 U154 ( .A1(n183), .A2(n182), .ZN(Y[13]) );
  AOI22_X1 U155 ( .A1(C[13]), .A2(n150), .B1(A[13]), .B2(n144), .ZN(n183) );
  AOI222_X1 U156 ( .A1(D[13]), .A2(n167), .B1(E[13]), .B2(n159), .C1(B[13]), 
        .C2(n153), .ZN(n182) );
  NAND2_X1 U157 ( .A1(n185), .A2(n184), .ZN(Y[14]) );
  AOI22_X1 U158 ( .A1(C[14]), .A2(n149), .B1(A[14]), .B2(n143), .ZN(n185) );
  AOI222_X1 U159 ( .A1(D[14]), .A2(n167), .B1(E[14]), .B2(n159), .C1(B[14]), 
        .C2(n153), .ZN(n184) );
  NAND2_X1 U160 ( .A1(n189), .A2(n188), .ZN(Y[16]) );
  AOI22_X1 U161 ( .A1(C[16]), .A2(n149), .B1(A[16]), .B2(n143), .ZN(n189) );
  AOI222_X1 U162 ( .A1(D[16]), .A2(n167), .B1(E[16]), .B2(n159), .C1(B[16]), 
        .C2(n153), .ZN(n188) );
  NAND2_X1 U163 ( .A1(n191), .A2(n190), .ZN(Y[17]) );
  AOI22_X1 U164 ( .A1(C[17]), .A2(n149), .B1(A[17]), .B2(n143), .ZN(n191) );
  AOI222_X1 U165 ( .A1(D[17]), .A2(n167), .B1(E[17]), .B2(n159), .C1(B[17]), 
        .C2(n153), .ZN(n190) );
  NAND2_X1 U166 ( .A1(n193), .A2(n192), .ZN(Y[18]) );
  AOI22_X1 U167 ( .A1(C[18]), .A2(n149), .B1(A[18]), .B2(n143), .ZN(n193) );
  AOI222_X1 U168 ( .A1(D[18]), .A2(n167), .B1(E[18]), .B2(n159), .C1(B[18]), 
        .C2(n153), .ZN(n192) );
  NAND2_X1 U169 ( .A1(n199), .A2(n198), .ZN(Y[20]) );
  AOI22_X1 U170 ( .A1(C[20]), .A2(n149), .B1(A[20]), .B2(n143), .ZN(n199) );
  AOI222_X1 U171 ( .A1(D[20]), .A2(n168), .B1(E[20]), .B2(n160), .C1(B[20]), 
        .C2(n154), .ZN(n198) );
  NAND2_X1 U172 ( .A1(n201), .A2(n200), .ZN(Y[21]) );
  AOI22_X1 U173 ( .A1(C[21]), .A2(n149), .B1(A[21]), .B2(n143), .ZN(n201) );
  AOI222_X1 U174 ( .A1(D[21]), .A2(n168), .B1(E[21]), .B2(n160), .C1(B[21]), 
        .C2(n154), .ZN(n200) );
  NAND2_X1 U175 ( .A1(n203), .A2(n202), .ZN(Y[22]) );
  AOI22_X1 U176 ( .A1(C[22]), .A2(n149), .B1(A[22]), .B2(n143), .ZN(n203) );
  AOI222_X1 U177 ( .A1(D[22]), .A2(n168), .B1(E[22]), .B2(n160), .C1(B[22]), 
        .C2(n154), .ZN(n202) );
  NAND2_X1 U178 ( .A1(n207), .A2(n206), .ZN(Y[24]) );
  AOI22_X1 U179 ( .A1(C[24]), .A2(n149), .B1(A[24]), .B2(n143), .ZN(n207) );
  AOI222_X1 U180 ( .A1(D[24]), .A2(n168), .B1(E[24]), .B2(n160), .C1(B[24]), 
        .C2(n154), .ZN(n206) );
  NAND2_X1 U181 ( .A1(n209), .A2(n208), .ZN(Y[25]) );
  AOI22_X1 U182 ( .A1(C[25]), .A2(n148), .B1(A[25]), .B2(n142), .ZN(n209) );
  AOI222_X1 U183 ( .A1(D[25]), .A2(n168), .B1(E[25]), .B2(n160), .C1(B[25]), 
        .C2(n154), .ZN(n208) );
  NAND2_X1 U184 ( .A1(n211), .A2(n210), .ZN(Y[26]) );
  AOI22_X1 U185 ( .A1(C[26]), .A2(n148), .B1(A[26]), .B2(n142), .ZN(n211) );
  AOI222_X1 U186 ( .A1(D[26]), .A2(n168), .B1(E[26]), .B2(n160), .C1(B[26]), 
        .C2(n154), .ZN(n210) );
  NAND2_X1 U187 ( .A1(n215), .A2(n214), .ZN(Y[28]) );
  AOI22_X1 U188 ( .A1(C[28]), .A2(n148), .B1(A[28]), .B2(n142), .ZN(n215) );
  AOI222_X1 U189 ( .A1(D[28]), .A2(n168), .B1(E[28]), .B2(n160), .C1(B[28]), 
        .C2(n154), .ZN(n214) );
  NAND2_X1 U190 ( .A1(n217), .A2(n216), .ZN(Y[29]) );
  AOI22_X1 U191 ( .A1(C[29]), .A2(n148), .B1(A[29]), .B2(n142), .ZN(n217) );
  AOI222_X1 U192 ( .A1(D[29]), .A2(n168), .B1(E[29]), .B2(n160), .C1(B[29]), 
        .C2(n154), .ZN(n216) );
  NAND2_X1 U193 ( .A1(n241), .A2(n240), .ZN(Y[3]) );
  AOI22_X1 U194 ( .A1(C[3]), .A2(n147), .B1(A[3]), .B2(n141), .ZN(n241) );
  AOI222_X1 U195 ( .A1(D[3]), .A2(n169), .B1(E[3]), .B2(n161), .C1(B[3]), .C2(
        n155), .ZN(n240) );
  NAND2_X1 U196 ( .A1(n297), .A2(n296), .ZN(Y[7]) );
  AOI22_X1 U197 ( .A1(C[7]), .A2(n145), .B1(A[7]), .B2(n139), .ZN(n297) );
  AOI222_X1 U198 ( .A1(D[7]), .A2(n171), .B1(E[7]), .B2(n164), .C1(B[7]), .C2(
        n157), .ZN(n296) );
  NAND2_X1 U199 ( .A1(n179), .A2(n178), .ZN(Y[11]) );
  AOI22_X1 U200 ( .A1(C[11]), .A2(n150), .B1(A[11]), .B2(n144), .ZN(n179) );
  AOI222_X1 U201 ( .A1(D[11]), .A2(n167), .B1(E[11]), .B2(n159), .C1(B[11]), 
        .C2(n153), .ZN(n178) );
  NAND2_X1 U202 ( .A1(n187), .A2(n186), .ZN(Y[15]) );
  AOI22_X1 U203 ( .A1(C[15]), .A2(n149), .B1(A[15]), .B2(n143), .ZN(n187) );
  AOI222_X1 U204 ( .A1(D[15]), .A2(n167), .B1(E[15]), .B2(n159), .C1(B[15]), 
        .C2(n153), .ZN(n186) );
  NAND2_X1 U205 ( .A1(n195), .A2(n194), .ZN(Y[19]) );
  AOI22_X1 U206 ( .A1(C[19]), .A2(n149), .B1(A[19]), .B2(n143), .ZN(n195) );
  AOI222_X1 U207 ( .A1(D[19]), .A2(n167), .B1(E[19]), .B2(n159), .C1(B[19]), 
        .C2(n153), .ZN(n194) );
  NAND2_X1 U208 ( .A1(n205), .A2(n204), .ZN(Y[23]) );
  AOI22_X1 U209 ( .A1(C[23]), .A2(n149), .B1(A[23]), .B2(n143), .ZN(n205) );
  AOI222_X1 U210 ( .A1(D[23]), .A2(n168), .B1(E[23]), .B2(n160), .C1(B[23]), 
        .C2(n154), .ZN(n204) );
  NAND2_X1 U211 ( .A1(n213), .A2(n212), .ZN(Y[27]) );
  AOI22_X1 U212 ( .A1(C[27]), .A2(n148), .B1(A[27]), .B2(n142), .ZN(n213) );
  AOI222_X1 U213 ( .A1(D[27]), .A2(n168), .B1(E[27]), .B2(n160), .C1(B[27]), 
        .C2(n154), .ZN(n212) );
  AOI22_X1 U214 ( .A1(C[58]), .A2(n145), .B1(A[58]), .B2(n139), .ZN(n281) );
  AOI22_X1 U215 ( .A1(C[57]), .A2(n145), .B1(A[57]), .B2(n139), .ZN(n279) );
  AOI222_X1 U216 ( .A1(D[57]), .A2(n171), .B1(E[57]), .B2(n163), .C1(B[57]), 
        .C2(n157), .ZN(n278) );
  AOI22_X1 U217 ( .A1(C[30]), .A2(n148), .B1(A[30]), .B2(n142), .ZN(n221) );
  AOI22_X1 U218 ( .A1(C[31]), .A2(n148), .B1(A[31]), .B2(n142), .ZN(n223) );
  AOI222_X1 U219 ( .A1(D[32]), .A2(n169), .B1(E[32]), .B2(n161), .C1(B[32]), 
        .C2(n155), .ZN(n224) );
  NAND2_X1 U220 ( .A1(n221), .A2(n220), .ZN(Y[30]) );
  NAND2_X1 U221 ( .A1(n223), .A2(n222), .ZN(Y[31]) );
  AOI222_X1 U222 ( .A1(D[35]), .A2(n169), .B1(E[35]), .B2(n161), .C1(B[35]), 
        .C2(n155), .ZN(n230) );
  AOI22_X1 U223 ( .A1(C[53]), .A2(n146), .B1(A[53]), .B2(n140), .ZN(n271) );
  AOI222_X1 U224 ( .A1(D[58]), .A2(n171), .B1(E[58]), .B2(n163), .C1(B[58]), 
        .C2(n157), .ZN(n280) );
  AOI222_X1 U225 ( .A1(D[53]), .A2(n170), .B1(E[53]), .B2(n163), .C1(B[53]), 
        .C2(n156), .ZN(n270) );
  AOI222_X1 U226 ( .A1(D[54]), .A2(n170), .B1(E[54]), .B2(n163), .C1(B[54]), 
        .C2(n156), .ZN(n272) );
  AOI22_X1 U227 ( .A1(C[61]), .A2(n145), .B1(A[61]), .B2(n139), .ZN(n289) );
  AOI222_X1 U228 ( .A1(D[61]), .A2(n171), .B1(E[61]), .B2(n163), .C1(B[61]), 
        .C2(n157), .ZN(n288) );
  AOI222_X1 U229 ( .A1(D[33]), .A2(n169), .B1(E[33]), .B2(n161), .C1(B[33]), 
        .C2(n155), .ZN(n226) );
  CLKBUF_X1 U230 ( .A(n300), .Z(n144) );
  CLKBUF_X1 U231 ( .A(n301), .Z(n150) );
  CLKBUF_X1 U232 ( .A(n158), .Z(n164) );
endmodule


module G_17 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_63 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_62 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_61 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_60 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_59 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_58 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_57 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_56 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_55 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_54 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_53 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_52 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_51 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_50 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_49 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_48 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_47 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_46 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_45 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_44 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_43 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_42 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_41 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_40 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_39 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_38 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_37 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_36 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_35 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_34 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_33 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_16 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_32 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_31 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_30 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_29 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_28 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_27 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_26 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_25 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_24 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_23 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_22 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_21 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(G_K_1), .B2(P_IK), .A(G_IK), .ZN(n4) );
endmodule


module PG_20 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_19 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AND2_X1 U3 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
endmodule


module PG_18 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module G_15 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_17 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_16 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_15 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_14 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_13 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_12 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_11 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_14 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_13 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_10 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_9 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_8 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
endmodule


module PG_7 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_6 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AND2_X1 U1 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U2 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_5 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(G_K_1), .A2(P_IK), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module G_12 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_11 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_10 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_9 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_4 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  AOI21_X1 U3 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module PG_3 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  OR2_X1 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_IK), .A2(P_K_1), .ZN(Px) );
endmodule


module PG_2 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module PG_1 ( G_IK, P_IK, G_K_1, P_K_1, Gx, Px );
  input G_IK, P_IK, G_K_1, P_K_1;
  output Gx, Px;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
  AND2_X1 U2 ( .A1(P_K_1), .A2(P_IK), .ZN(Px) );
  INV_X1 U3 ( .A(n4), .ZN(Gx) );
endmodule


module G_8 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_7 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X2 U1 ( .A1(G_IK), .A2(n4), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_6 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_5 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G_IK), .ZN(Gx) );
  AND2_X1 U2 ( .A1(P_IK), .A2(G_K_1), .ZN(n4) );
endmodule


module G_4 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_3 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_2 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module G_1 ( G_IK, P_IK, G_K_1, Gx );
  input G_IK, P_IK, G_K_1;
  output Gx;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gx) );
  AOI21_X1 U2 ( .B1(P_IK), .B2(G_K_1), .A(G_IK), .ZN(n4) );
endmodule


module carry_generator_N64_NPB4_1 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   \PG_Network[5][1][63] , \PG_Network[5][1][59] ,
         \PG_Network[5][1][55] , \PG_Network[5][1][51] ,
         \PG_Network[5][0][63] , \PG_Network[5][0][59] ,
         \PG_Network[5][0][55] , \PG_Network[5][0][51] ,
         \PG_Network[4][1][63] , \PG_Network[4][1][59] ,
         \PG_Network[4][1][47] , \PG_Network[4][1][43] ,
         \PG_Network[4][1][31] , \PG_Network[4][1][27] ,
         \PG_Network[4][0][63] , \PG_Network[4][0][59] ,
         \PG_Network[4][0][47] , \PG_Network[4][0][43] ,
         \PG_Network[4][0][31] , \PG_Network[4][0][27] ,
         \PG_Network[3][1][63] , \PG_Network[3][1][55] ,
         \PG_Network[3][1][47] , \PG_Network[3][1][39] ,
         \PG_Network[3][1][31] , \PG_Network[3][1][23] ,
         \PG_Network[3][1][15] , \PG_Network[3][0][63] ,
         \PG_Network[3][0][55] , \PG_Network[3][0][47] ,
         \PG_Network[3][0][39] , \PG_Network[3][0][31] ,
         \PG_Network[3][0][23] , \PG_Network[3][0][15] ,
         \PG_Network[2][1][63] , \PG_Network[2][1][59] ,
         \PG_Network[2][1][55] , \PG_Network[2][1][51] ,
         \PG_Network[2][1][47] , \PG_Network[2][1][43] ,
         \PG_Network[2][1][39] , \PG_Network[2][1][35] ,
         \PG_Network[2][1][31] , \PG_Network[2][1][27] ,
         \PG_Network[2][1][23] , \PG_Network[2][1][19] ,
         \PG_Network[2][1][15] , \PG_Network[2][1][11] , \PG_Network[2][1][7] ,
         \PG_Network[2][0][63] , \PG_Network[2][0][59] ,
         \PG_Network[2][0][55] , \PG_Network[2][0][51] ,
         \PG_Network[2][0][47] , \PG_Network[2][0][43] ,
         \PG_Network[2][0][39] , \PG_Network[2][0][35] ,
         \PG_Network[2][0][31] , \PG_Network[2][0][27] ,
         \PG_Network[2][0][23] , \PG_Network[2][0][19] ,
         \PG_Network[2][0][15] , \PG_Network[2][0][11] , \PG_Network[2][0][7] ,
         \PG_Network[1][1][63] , \PG_Network[1][1][61] ,
         \PG_Network[1][1][59] , \PG_Network[1][1][57] ,
         \PG_Network[1][1][55] , \PG_Network[1][1][53] ,
         \PG_Network[1][1][51] , \PG_Network[1][1][49] ,
         \PG_Network[1][1][47] , \PG_Network[1][1][45] ,
         \PG_Network[1][1][43] , \PG_Network[1][1][41] ,
         \PG_Network[1][1][39] , \PG_Network[1][1][37] ,
         \PG_Network[1][1][35] , \PG_Network[1][1][33] ,
         \PG_Network[1][1][31] , \PG_Network[1][1][29] ,
         \PG_Network[1][1][27] , \PG_Network[1][1][25] ,
         \PG_Network[1][1][23] , \PG_Network[1][1][21] ,
         \PG_Network[1][1][19] , \PG_Network[1][1][17] ,
         \PG_Network[1][1][15] , \PG_Network[1][1][13] ,
         \PG_Network[1][1][11] , \PG_Network[1][1][9] , \PG_Network[1][1][7] ,
         \PG_Network[1][1][5] , \PG_Network[1][1][3] , \PG_Network[1][1][1] ,
         \PG_Network[1][0][63] , \PG_Network[1][0][61] ,
         \PG_Network[1][0][59] , \PG_Network[1][0][57] ,
         \PG_Network[1][0][55] , \PG_Network[1][0][53] ,
         \PG_Network[1][0][51] , \PG_Network[1][0][49] ,
         \PG_Network[1][0][47] , \PG_Network[1][0][45] ,
         \PG_Network[1][0][43] , \PG_Network[1][0][41] ,
         \PG_Network[1][0][39] , \PG_Network[1][0][37] ,
         \PG_Network[1][0][35] , \PG_Network[1][0][33] ,
         \PG_Network[1][0][31] , \PG_Network[1][0][29] ,
         \PG_Network[1][0][27] , \PG_Network[1][0][25] ,
         \PG_Network[1][0][23] , \PG_Network[1][0][21] ,
         \PG_Network[1][0][19] , \PG_Network[1][0][17] ,
         \PG_Network[1][0][15] , \PG_Network[1][0][13] ,
         \PG_Network[1][0][11] , \PG_Network[1][0][9] , \PG_Network[1][0][7] ,
         \PG_Network[1][0][5] , \PG_Network[1][0][3] , \PG_Network[0][1][63] ,
         \PG_Network[0][1][62] , \PG_Network[0][1][61] ,
         \PG_Network[0][1][60] , \PG_Network[0][1][59] ,
         \PG_Network[0][1][58] , \PG_Network[0][1][57] ,
         \PG_Network[0][1][56] , \PG_Network[0][1][55] ,
         \PG_Network[0][1][54] , \PG_Network[0][1][53] ,
         \PG_Network[0][1][52] , \PG_Network[0][1][51] ,
         \PG_Network[0][1][50] , \PG_Network[0][1][49] ,
         \PG_Network[0][1][48] , \PG_Network[0][1][47] ,
         \PG_Network[0][1][46] , \PG_Network[0][1][45] ,
         \PG_Network[0][1][44] , \PG_Network[0][1][43] ,
         \PG_Network[0][1][42] , \PG_Network[0][1][41] ,
         \PG_Network[0][1][40] , \PG_Network[0][1][39] ,
         \PG_Network[0][1][38] , \PG_Network[0][1][37] ,
         \PG_Network[0][1][36] , \PG_Network[0][1][35] ,
         \PG_Network[0][1][34] , \PG_Network[0][1][33] ,
         \PG_Network[0][1][32] , \PG_Network[0][1][31] ,
         \PG_Network[0][1][30] , \PG_Network[0][1][29] ,
         \PG_Network[0][1][28] , \PG_Network[0][1][27] ,
         \PG_Network[0][1][26] , \PG_Network[0][1][25] ,
         \PG_Network[0][1][24] , \PG_Network[0][1][23] ,
         \PG_Network[0][1][22] , \PG_Network[0][1][21] ,
         \PG_Network[0][1][20] , \PG_Network[0][1][19] ,
         \PG_Network[0][1][18] , \PG_Network[0][1][17] ,
         \PG_Network[0][1][16] , \PG_Network[0][1][15] ,
         \PG_Network[0][1][14] , \PG_Network[0][1][13] ,
         \PG_Network[0][1][12] , \PG_Network[0][1][11] ,
         \PG_Network[0][1][10] , \PG_Network[0][1][9] , \PG_Network[0][1][8] ,
         \PG_Network[0][1][7] , \PG_Network[0][1][6] , \PG_Network[0][1][5] ,
         \PG_Network[0][1][4] , \PG_Network[0][1][3] , \PG_Network[0][1][2] ,
         \PG_Network[0][1][1] , \PG_Network[0][0][63] , \PG_Network[0][0][62] ,
         \PG_Network[0][0][61] , \PG_Network[0][0][60] ,
         \PG_Network[0][0][59] , \PG_Network[0][0][58] ,
         \PG_Network[0][0][57] , \PG_Network[0][0][56] ,
         \PG_Network[0][0][55] , \PG_Network[0][0][54] ,
         \PG_Network[0][0][53] , \PG_Network[0][0][52] ,
         \PG_Network[0][0][51] , \PG_Network[0][0][50] ,
         \PG_Network[0][0][49] , \PG_Network[0][0][48] ,
         \PG_Network[0][0][47] , \PG_Network[0][0][46] ,
         \PG_Network[0][0][45] , \PG_Network[0][0][44] ,
         \PG_Network[0][0][43] , \PG_Network[0][0][42] ,
         \PG_Network[0][0][41] , \PG_Network[0][0][40] ,
         \PG_Network[0][0][39] , \PG_Network[0][0][38] ,
         \PG_Network[0][0][37] , \PG_Network[0][0][36] ,
         \PG_Network[0][0][35] , \PG_Network[0][0][34] ,
         \PG_Network[0][0][33] , \PG_Network[0][0][32] ,
         \PG_Network[0][0][31] , \PG_Network[0][0][30] ,
         \PG_Network[0][0][29] , \PG_Network[0][0][28] ,
         \PG_Network[0][0][27] , \PG_Network[0][0][26] ,
         \PG_Network[0][0][25] , \PG_Network[0][0][24] ,
         \PG_Network[0][0][23] , \PG_Network[0][0][22] ,
         \PG_Network[0][0][21] , \PG_Network[0][0][20] ,
         \PG_Network[0][0][19] , \PG_Network[0][0][18] ,
         \PG_Network[0][0][17] , \PG_Network[0][0][16] ,
         \PG_Network[0][0][15] , \PG_Network[0][0][14] ,
         \PG_Network[0][0][13] , \PG_Network[0][0][12] ,
         \PG_Network[0][0][11] , \PG_Network[0][0][10] , \PG_Network[0][0][9] ,
         \PG_Network[0][0][8] , \PG_Network[0][0][7] , \PG_Network[0][0][6] ,
         \PG_Network[0][0][5] , \PG_Network[0][0][4] , \PG_Network[0][0][3] ,
         \PG_Network[0][0][2] , \PG_Network[0][0][1] , n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18;

  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(\PG_Network[0][0][9] ) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(\PG_Network[0][0][8] ) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(\PG_Network[0][0][7] ) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(\PG_Network[0][0][6] ) );
  XOR2_X1 U72 ( .A(B[63]), .B(A[63]), .Z(\PG_Network[0][0][63] ) );
  XOR2_X1 U73 ( .A(B[62]), .B(A[62]), .Z(\PG_Network[0][0][62] ) );
  XOR2_X1 U74 ( .A(B[61]), .B(A[61]), .Z(\PG_Network[0][0][61] ) );
  XOR2_X1 U75 ( .A(B[60]), .B(A[60]), .Z(\PG_Network[0][0][60] ) );
  XOR2_X1 U76 ( .A(B[5]), .B(A[5]), .Z(\PG_Network[0][0][5] ) );
  XOR2_X1 U78 ( .A(B[58]), .B(A[58]), .Z(\PG_Network[0][0][58] ) );
  XOR2_X1 U80 ( .A(B[56]), .B(A[56]), .Z(\PG_Network[0][0][56] ) );
  XOR2_X1 U82 ( .A(B[54]), .B(A[54]), .Z(\PG_Network[0][0][54] ) );
  XOR2_X1 U84 ( .A(B[52]), .B(A[52]), .Z(\PG_Network[0][0][52] ) );
  XOR2_X1 U86 ( .A(B[50]), .B(A[50]), .Z(\PG_Network[0][0][50] ) );
  XOR2_X1 U87 ( .A(B[4]), .B(A[4]), .Z(\PG_Network[0][0][4] ) );
  XOR2_X1 U88 ( .A(B[49]), .B(A[49]), .Z(\PG_Network[0][0][49] ) );
  XOR2_X1 U89 ( .A(B[48]), .B(A[48]), .Z(\PG_Network[0][0][48] ) );
  XOR2_X1 U91 ( .A(B[46]), .B(A[46]), .Z(\PG_Network[0][0][46] ) );
  XOR2_X1 U92 ( .A(B[45]), .B(A[45]), .Z(\PG_Network[0][0][45] ) );
  XOR2_X1 U93 ( .A(B[44]), .B(A[44]), .Z(\PG_Network[0][0][44] ) );
  XOR2_X1 U95 ( .A(B[42]), .B(A[42]), .Z(\PG_Network[0][0][42] ) );
  XOR2_X1 U96 ( .A(B[41]), .B(A[41]), .Z(\PG_Network[0][0][41] ) );
  XOR2_X1 U97 ( .A(B[40]), .B(A[40]), .Z(\PG_Network[0][0][40] ) );
  XOR2_X1 U98 ( .A(B[3]), .B(A[3]), .Z(\PG_Network[0][0][3] ) );
  XOR2_X1 U99 ( .A(B[39]), .B(A[39]), .Z(\PG_Network[0][0][39] ) );
  XOR2_X1 U100 ( .A(B[38]), .B(A[38]), .Z(\PG_Network[0][0][38] ) );
  XOR2_X1 U101 ( .A(B[37]), .B(A[37]), .Z(\PG_Network[0][0][37] ) );
  XOR2_X1 U102 ( .A(B[36]), .B(A[36]), .Z(\PG_Network[0][0][36] ) );
  XOR2_X1 U103 ( .A(B[35]), .B(A[35]), .Z(\PG_Network[0][0][35] ) );
  XOR2_X1 U104 ( .A(B[34]), .B(A[34]), .Z(\PG_Network[0][0][34] ) );
  XOR2_X1 U105 ( .A(B[33]), .B(A[33]), .Z(\PG_Network[0][0][33] ) );
  XOR2_X1 U106 ( .A(B[32]), .B(A[32]), .Z(\PG_Network[0][0][32] ) );
  XOR2_X1 U107 ( .A(B[31]), .B(A[31]), .Z(\PG_Network[0][0][31] ) );
  XOR2_X1 U108 ( .A(B[30]), .B(A[30]), .Z(\PG_Network[0][0][30] ) );
  XOR2_X1 U109 ( .A(B[2]), .B(A[2]), .Z(\PG_Network[0][0][2] ) );
  XOR2_X1 U110 ( .A(B[29]), .B(A[29]), .Z(\PG_Network[0][0][29] ) );
  XOR2_X1 U111 ( .A(B[28]), .B(A[28]), .Z(\PG_Network[0][0][28] ) );
  XOR2_X1 U112 ( .A(B[27]), .B(A[27]), .Z(\PG_Network[0][0][27] ) );
  XOR2_X1 U113 ( .A(B[26]), .B(A[26]), .Z(\PG_Network[0][0][26] ) );
  XOR2_X1 U114 ( .A(B[25]), .B(A[25]), .Z(\PG_Network[0][0][25] ) );
  XOR2_X1 U115 ( .A(B[24]), .B(A[24]), .Z(\PG_Network[0][0][24] ) );
  XOR2_X1 U116 ( .A(B[23]), .B(A[23]), .Z(\PG_Network[0][0][23] ) );
  XOR2_X1 U117 ( .A(B[22]), .B(A[22]), .Z(\PG_Network[0][0][22] ) );
  XOR2_X1 U118 ( .A(B[21]), .B(A[21]), .Z(\PG_Network[0][0][21] ) );
  XOR2_X1 U119 ( .A(B[20]), .B(A[20]), .Z(\PG_Network[0][0][20] ) );
  XOR2_X1 U120 ( .A(B[1]), .B(A[1]), .Z(\PG_Network[0][0][1] ) );
  XOR2_X1 U121 ( .A(B[19]), .B(A[19]), .Z(\PG_Network[0][0][19] ) );
  XOR2_X1 U122 ( .A(B[18]), .B(A[18]), .Z(\PG_Network[0][0][18] ) );
  XOR2_X1 U123 ( .A(B[17]), .B(A[17]), .Z(\PG_Network[0][0][17] ) );
  XOR2_X1 U124 ( .A(B[16]), .B(A[16]), .Z(\PG_Network[0][0][16] ) );
  XOR2_X1 U125 ( .A(B[15]), .B(A[15]), .Z(\PG_Network[0][0][15] ) );
  XOR2_X1 U126 ( .A(B[14]), .B(A[14]), .Z(\PG_Network[0][0][14] ) );
  XOR2_X1 U127 ( .A(B[13]), .B(A[13]), .Z(\PG_Network[0][0][13] ) );
  XOR2_X1 U128 ( .A(B[12]), .B(A[12]), .Z(\PG_Network[0][0][12] ) );
  XOR2_X1 U129 ( .A(B[11]), .B(A[11]), .Z(\PG_Network[0][0][11] ) );
  XOR2_X1 U130 ( .A(B[10]), .B(A[10]), .Z(\PG_Network[0][0][10] ) );
  G_17 GJ_0_0_0 ( .G_IK(\PG_Network[0][1][1] ), .P_IK(\PG_Network[0][0][1] ), 
        .G_K_1(n15), .Gx(\PG_Network[1][1][1] ) );
  PG_63 PGJ_0_1_0 ( .G_IK(\PG_Network[0][1][3] ), .P_IK(\PG_Network[0][0][3] ), 
        .G_K_1(\PG_Network[0][1][2] ), .P_K_1(\PG_Network[0][0][2] ), .Gx(
        \PG_Network[1][1][3] ), .Px(\PG_Network[1][0][3] ) );
  PG_62 PGJ_0_2_0 ( .G_IK(\PG_Network[0][1][5] ), .P_IK(\PG_Network[0][0][5] ), 
        .G_K_1(\PG_Network[0][1][4] ), .P_K_1(\PG_Network[0][0][4] ), .Gx(
        \PG_Network[1][1][5] ), .Px(\PG_Network[1][0][5] ) );
  PG_61 PGJ_0_3_0 ( .G_IK(\PG_Network[0][1][7] ), .P_IK(\PG_Network[0][0][7] ), 
        .G_K_1(\PG_Network[0][1][6] ), .P_K_1(\PG_Network[0][0][6] ), .Gx(
        \PG_Network[1][1][7] ), .Px(\PG_Network[1][0][7] ) );
  PG_60 PGJ_0_4_0 ( .G_IK(\PG_Network[0][1][9] ), .P_IK(\PG_Network[0][0][9] ), 
        .G_K_1(\PG_Network[0][1][8] ), .P_K_1(\PG_Network[0][0][8] ), .Gx(
        \PG_Network[1][1][9] ), .Px(\PG_Network[1][0][9] ) );
  PG_59 PGJ_0_5_0 ( .G_IK(\PG_Network[0][1][11] ), .P_IK(
        \PG_Network[0][0][11] ), .G_K_1(\PG_Network[0][1][10] ), .P_K_1(
        \PG_Network[0][0][10] ), .Gx(\PG_Network[1][1][11] ), .Px(
        \PG_Network[1][0][11] ) );
  PG_58 PGJ_0_6_0 ( .G_IK(\PG_Network[0][1][13] ), .P_IK(
        \PG_Network[0][0][13] ), .G_K_1(\PG_Network[0][1][12] ), .P_K_1(
        \PG_Network[0][0][12] ), .Gx(\PG_Network[1][1][13] ), .Px(
        \PG_Network[1][0][13] ) );
  PG_57 PGJ_0_7_0 ( .G_IK(\PG_Network[0][1][15] ), .P_IK(
        \PG_Network[0][0][15] ), .G_K_1(\PG_Network[0][1][14] ), .P_K_1(
        \PG_Network[0][0][14] ), .Gx(\PG_Network[1][1][15] ), .Px(
        \PG_Network[1][0][15] ) );
  PG_56 PGJ_0_8_0 ( .G_IK(\PG_Network[0][1][17] ), .P_IK(
        \PG_Network[0][0][17] ), .G_K_1(\PG_Network[0][1][16] ), .P_K_1(
        \PG_Network[0][0][16] ), .Gx(\PG_Network[1][1][17] ), .Px(
        \PG_Network[1][0][17] ) );
  PG_55 PGJ_0_9_0 ( .G_IK(\PG_Network[0][1][19] ), .P_IK(
        \PG_Network[0][0][19] ), .G_K_1(\PG_Network[0][1][18] ), .P_K_1(
        \PG_Network[0][0][18] ), .Gx(\PG_Network[1][1][19] ), .Px(
        \PG_Network[1][0][19] ) );
  PG_54 PGJ_0_10_0 ( .G_IK(\PG_Network[0][1][21] ), .P_IK(
        \PG_Network[0][0][21] ), .G_K_1(\PG_Network[0][1][20] ), .P_K_1(
        \PG_Network[0][0][20] ), .Gx(\PG_Network[1][1][21] ), .Px(
        \PG_Network[1][0][21] ) );
  PG_53 PGJ_0_11_0 ( .G_IK(\PG_Network[0][1][23] ), .P_IK(
        \PG_Network[0][0][23] ), .G_K_1(\PG_Network[0][1][22] ), .P_K_1(
        \PG_Network[0][0][22] ), .Gx(\PG_Network[1][1][23] ), .Px(
        \PG_Network[1][0][23] ) );
  PG_52 PGJ_0_12_0 ( .G_IK(\PG_Network[0][1][25] ), .P_IK(
        \PG_Network[0][0][25] ), .G_K_1(\PG_Network[0][1][24] ), .P_K_1(
        \PG_Network[0][0][24] ), .Gx(\PG_Network[1][1][25] ), .Px(
        \PG_Network[1][0][25] ) );
  PG_51 PGJ_0_13_0 ( .G_IK(\PG_Network[0][1][27] ), .P_IK(
        \PG_Network[0][0][27] ), .G_K_1(\PG_Network[0][1][26] ), .P_K_1(
        \PG_Network[0][0][26] ), .Gx(\PG_Network[1][1][27] ), .Px(
        \PG_Network[1][0][27] ) );
  PG_50 PGJ_0_14_0 ( .G_IK(\PG_Network[0][1][29] ), .P_IK(
        \PG_Network[0][0][29] ), .G_K_1(\PG_Network[0][1][28] ), .P_K_1(
        \PG_Network[0][0][28] ), .Gx(\PG_Network[1][1][29] ), .Px(
        \PG_Network[1][0][29] ) );
  PG_49 PGJ_0_15_0 ( .G_IK(\PG_Network[0][1][31] ), .P_IK(
        \PG_Network[0][0][31] ), .G_K_1(\PG_Network[0][1][30] ), .P_K_1(
        \PG_Network[0][0][30] ), .Gx(\PG_Network[1][1][31] ), .Px(
        \PG_Network[1][0][31] ) );
  PG_48 PGJ_0_16_0 ( .G_IK(\PG_Network[0][1][33] ), .P_IK(
        \PG_Network[0][0][33] ), .G_K_1(\PG_Network[0][1][32] ), .P_K_1(
        \PG_Network[0][0][32] ), .Gx(\PG_Network[1][1][33] ), .Px(
        \PG_Network[1][0][33] ) );
  PG_47 PGJ_0_17_0 ( .G_IK(\PG_Network[0][1][35] ), .P_IK(
        \PG_Network[0][0][35] ), .G_K_1(\PG_Network[0][1][34] ), .P_K_1(
        \PG_Network[0][0][34] ), .Gx(\PG_Network[1][1][35] ), .Px(
        \PG_Network[1][0][35] ) );
  PG_46 PGJ_0_18_0 ( .G_IK(\PG_Network[0][1][37] ), .P_IK(
        \PG_Network[0][0][37] ), .G_K_1(\PG_Network[0][1][36] ), .P_K_1(
        \PG_Network[0][0][36] ), .Gx(\PG_Network[1][1][37] ), .Px(
        \PG_Network[1][0][37] ) );
  PG_45 PGJ_0_19_0 ( .G_IK(\PG_Network[0][1][39] ), .P_IK(
        \PG_Network[0][0][39] ), .G_K_1(\PG_Network[0][1][38] ), .P_K_1(
        \PG_Network[0][0][38] ), .Gx(\PG_Network[1][1][39] ), .Px(
        \PG_Network[1][0][39] ) );
  PG_44 PGJ_0_20_0 ( .G_IK(\PG_Network[0][1][41] ), .P_IK(
        \PG_Network[0][0][41] ), .G_K_1(\PG_Network[0][1][40] ), .P_K_1(
        \PG_Network[0][0][40] ), .Gx(\PG_Network[1][1][41] ), .Px(
        \PG_Network[1][0][41] ) );
  PG_43 PGJ_0_21_0 ( .G_IK(\PG_Network[0][1][43] ), .P_IK(
        \PG_Network[0][0][43] ), .G_K_1(\PG_Network[0][1][42] ), .P_K_1(
        \PG_Network[0][0][42] ), .Gx(\PG_Network[1][1][43] ), .Px(
        \PG_Network[1][0][43] ) );
  PG_42 PGJ_0_22_0 ( .G_IK(\PG_Network[0][1][45] ), .P_IK(
        \PG_Network[0][0][45] ), .G_K_1(\PG_Network[0][1][44] ), .P_K_1(
        \PG_Network[0][0][44] ), .Gx(\PG_Network[1][1][45] ), .Px(
        \PG_Network[1][0][45] ) );
  PG_41 PGJ_0_23_0 ( .G_IK(\PG_Network[0][1][47] ), .P_IK(
        \PG_Network[0][0][47] ), .G_K_1(\PG_Network[0][1][46] ), .P_K_1(
        \PG_Network[0][0][46] ), .Gx(\PG_Network[1][1][47] ), .Px(
        \PG_Network[1][0][47] ) );
  PG_40 PGJ_0_24_0 ( .G_IK(\PG_Network[0][1][49] ), .P_IK(
        \PG_Network[0][0][49] ), .G_K_1(\PG_Network[0][1][48] ), .P_K_1(
        \PG_Network[0][0][48] ), .Gx(\PG_Network[1][1][49] ), .Px(
        \PG_Network[1][0][49] ) );
  PG_39 PGJ_0_25_0 ( .G_IK(\PG_Network[0][1][51] ), .P_IK(
        \PG_Network[0][0][51] ), .G_K_1(\PG_Network[0][1][50] ), .P_K_1(
        \PG_Network[0][0][50] ), .Gx(\PG_Network[1][1][51] ), .Px(
        \PG_Network[1][0][51] ) );
  PG_38 PGJ_0_26_0 ( .G_IK(\PG_Network[0][1][53] ), .P_IK(
        \PG_Network[0][0][53] ), .G_K_1(\PG_Network[0][1][52] ), .P_K_1(
        \PG_Network[0][0][52] ), .Gx(\PG_Network[1][1][53] ), .Px(
        \PG_Network[1][0][53] ) );
  PG_37 PGJ_0_27_0 ( .G_IK(\PG_Network[0][1][55] ), .P_IK(
        \PG_Network[0][0][55] ), .G_K_1(\PG_Network[0][1][54] ), .P_K_1(
        \PG_Network[0][0][54] ), .Gx(\PG_Network[1][1][55] ), .Px(
        \PG_Network[1][0][55] ) );
  PG_36 PGJ_0_28_0 ( .G_IK(\PG_Network[0][1][57] ), .P_IK(
        \PG_Network[0][0][57] ), .G_K_1(\PG_Network[0][1][56] ), .P_K_1(
        \PG_Network[0][0][56] ), .Gx(\PG_Network[1][1][57] ), .Px(
        \PG_Network[1][0][57] ) );
  PG_35 PGJ_0_29_0 ( .G_IK(\PG_Network[0][1][59] ), .P_IK(
        \PG_Network[0][0][59] ), .G_K_1(\PG_Network[0][1][58] ), .P_K_1(
        \PG_Network[0][0][58] ), .Gx(\PG_Network[1][1][59] ), .Px(
        \PG_Network[1][0][59] ) );
  PG_34 PGJ_0_30_0 ( .G_IK(\PG_Network[0][1][61] ), .P_IK(
        \PG_Network[0][0][61] ), .G_K_1(\PG_Network[0][1][60] ), .P_K_1(
        \PG_Network[0][0][60] ), .Gx(\PG_Network[1][1][61] ), .Px(
        \PG_Network[1][0][61] ) );
  PG_33 PGJ_0_31_0 ( .G_IK(\PG_Network[0][1][63] ), .P_IK(
        \PG_Network[0][0][63] ), .G_K_1(\PG_Network[0][1][62] ), .P_K_1(
        \PG_Network[0][0][62] ), .Gx(\PG_Network[1][1][63] ), .Px(
        \PG_Network[1][0][63] ) );
  G_16 GJ_1_0_0 ( .G_IK(\PG_Network[1][1][3] ), .P_IK(\PG_Network[1][0][3] ), 
        .G_K_1(\PG_Network[1][1][1] ), .Gx(Co[0]) );
  PG_32 PGJ_1_1_0 ( .G_IK(\PG_Network[1][1][7] ), .P_IK(\PG_Network[1][0][7] ), 
        .G_K_1(\PG_Network[1][1][5] ), .P_K_1(\PG_Network[1][0][5] ), .Gx(
        \PG_Network[2][1][7] ), .Px(\PG_Network[2][0][7] ) );
  PG_31 PGJ_1_2_0 ( .G_IK(\PG_Network[1][1][11] ), .P_IK(
        \PG_Network[1][0][11] ), .G_K_1(\PG_Network[1][1][9] ), .P_K_1(
        \PG_Network[1][0][9] ), .Gx(\PG_Network[2][1][11] ), .Px(
        \PG_Network[2][0][11] ) );
  PG_30 PGJ_1_3_0 ( .G_IK(\PG_Network[1][1][15] ), .P_IK(
        \PG_Network[1][0][15] ), .G_K_1(\PG_Network[1][1][13] ), .P_K_1(
        \PG_Network[1][0][13] ), .Gx(\PG_Network[2][1][15] ), .Px(
        \PG_Network[2][0][15] ) );
  PG_29 PGJ_1_4_0 ( .G_IK(\PG_Network[1][1][19] ), .P_IK(
        \PG_Network[1][0][19] ), .G_K_1(\PG_Network[1][1][17] ), .P_K_1(
        \PG_Network[1][0][17] ), .Gx(\PG_Network[2][1][19] ), .Px(
        \PG_Network[2][0][19] ) );
  PG_28 PGJ_1_5_0 ( .G_IK(\PG_Network[1][1][23] ), .P_IK(
        \PG_Network[1][0][23] ), .G_K_1(\PG_Network[1][1][21] ), .P_K_1(
        \PG_Network[1][0][21] ), .Gx(\PG_Network[2][1][23] ), .Px(
        \PG_Network[2][0][23] ) );
  PG_27 PGJ_1_6_0 ( .G_IK(\PG_Network[1][1][27] ), .P_IK(
        \PG_Network[1][0][27] ), .G_K_1(\PG_Network[1][1][25] ), .P_K_1(
        \PG_Network[1][0][25] ), .Gx(\PG_Network[2][1][27] ), .Px(
        \PG_Network[2][0][27] ) );
  PG_26 PGJ_1_7_0 ( .G_IK(\PG_Network[1][1][31] ), .P_IK(
        \PG_Network[1][0][31] ), .G_K_1(\PG_Network[1][1][29] ), .P_K_1(
        \PG_Network[1][0][29] ), .Gx(\PG_Network[2][1][31] ), .Px(
        \PG_Network[2][0][31] ) );
  PG_25 PGJ_1_8_0 ( .G_IK(\PG_Network[1][1][35] ), .P_IK(
        \PG_Network[1][0][35] ), .G_K_1(\PG_Network[1][1][33] ), .P_K_1(
        \PG_Network[1][0][33] ), .Gx(\PG_Network[2][1][35] ), .Px(
        \PG_Network[2][0][35] ) );
  PG_24 PGJ_1_9_0 ( .G_IK(\PG_Network[1][1][39] ), .P_IK(
        \PG_Network[1][0][39] ), .G_K_1(\PG_Network[1][1][37] ), .P_K_1(
        \PG_Network[1][0][37] ), .Gx(\PG_Network[2][1][39] ), .Px(
        \PG_Network[2][0][39] ) );
  PG_23 PGJ_1_10_0 ( .G_IK(\PG_Network[1][1][43] ), .P_IK(
        \PG_Network[1][0][43] ), .G_K_1(\PG_Network[1][1][41] ), .P_K_1(
        \PG_Network[1][0][41] ), .Gx(\PG_Network[2][1][43] ), .Px(
        \PG_Network[2][0][43] ) );
  PG_22 PGJ_1_11_0 ( .G_IK(\PG_Network[1][1][47] ), .P_IK(
        \PG_Network[1][0][47] ), .G_K_1(\PG_Network[1][1][45] ), .P_K_1(
        \PG_Network[1][0][45] ), .Gx(\PG_Network[2][1][47] ), .Px(
        \PG_Network[2][0][47] ) );
  PG_21 PGJ_1_12_0 ( .G_IK(\PG_Network[1][1][51] ), .P_IK(
        \PG_Network[1][0][51] ), .G_K_1(\PG_Network[1][1][49] ), .P_K_1(
        \PG_Network[1][0][49] ), .Gx(\PG_Network[2][1][51] ), .Px(
        \PG_Network[2][0][51] ) );
  PG_20 PGJ_1_13_0 ( .G_IK(\PG_Network[1][1][55] ), .P_IK(
        \PG_Network[1][0][55] ), .G_K_1(\PG_Network[1][1][53] ), .P_K_1(
        \PG_Network[1][0][53] ), .Gx(\PG_Network[2][1][55] ), .Px(
        \PG_Network[2][0][55] ) );
  PG_19 PGJ_1_14_0 ( .G_IK(\PG_Network[1][1][59] ), .P_IK(
        \PG_Network[1][0][59] ), .G_K_1(\PG_Network[1][1][57] ), .P_K_1(
        \PG_Network[1][0][57] ), .Gx(\PG_Network[2][1][59] ), .Px(
        \PG_Network[2][0][59] ) );
  PG_18 PGJ_1_15_0 ( .G_IK(\PG_Network[1][1][63] ), .P_IK(
        \PG_Network[1][0][63] ), .G_K_1(\PG_Network[1][1][61] ), .P_K_1(
        \PG_Network[1][0][61] ), .Gx(\PG_Network[2][1][63] ), .Px(
        \PG_Network[2][0][63] ) );
  G_15 GJ_2_0_0 ( .G_IK(\PG_Network[2][1][7] ), .P_IK(\PG_Network[2][0][7] ), 
        .G_K_1(Co[0]), .Gx(Co[1]) );
  PG_17 PGJ_2_1_0 ( .G_IK(\PG_Network[2][1][15] ), .P_IK(
        \PG_Network[2][0][15] ), .G_K_1(\PG_Network[2][1][11] ), .P_K_1(
        \PG_Network[2][0][11] ), .Gx(\PG_Network[3][1][15] ), .Px(
        \PG_Network[3][0][15] ) );
  PG_16 PGJ_2_2_0 ( .G_IK(\PG_Network[2][1][23] ), .P_IK(
        \PG_Network[2][0][23] ), .G_K_1(\PG_Network[2][1][19] ), .P_K_1(
        \PG_Network[2][0][19] ), .Gx(\PG_Network[3][1][23] ), .Px(
        \PG_Network[3][0][23] ) );
  PG_15 PGJ_2_3_0 ( .G_IK(\PG_Network[2][1][31] ), .P_IK(
        \PG_Network[2][0][31] ), .G_K_1(\PG_Network[2][1][27] ), .P_K_1(
        \PG_Network[2][0][27] ), .Gx(\PG_Network[3][1][31] ), .Px(
        \PG_Network[3][0][31] ) );
  PG_14 PGJ_2_4_0 ( .G_IK(\PG_Network[2][1][39] ), .P_IK(
        \PG_Network[2][0][39] ), .G_K_1(\PG_Network[2][1][35] ), .P_K_1(
        \PG_Network[2][0][35] ), .Gx(\PG_Network[3][1][39] ), .Px(
        \PG_Network[3][0][39] ) );
  PG_13 PGJ_2_5_0 ( .G_IK(\PG_Network[2][1][47] ), .P_IK(
        \PG_Network[2][0][47] ), .G_K_1(\PG_Network[2][1][43] ), .P_K_1(
        \PG_Network[2][0][43] ), .Gx(\PG_Network[3][1][47] ), .Px(
        \PG_Network[3][0][47] ) );
  PG_12 PGJ_2_6_0 ( .G_IK(\PG_Network[2][1][55] ), .P_IK(
        \PG_Network[2][0][55] ), .G_K_1(\PG_Network[2][1][51] ), .P_K_1(
        \PG_Network[2][0][51] ), .Gx(\PG_Network[3][1][55] ), .Px(
        \PG_Network[3][0][55] ) );
  PG_11 PGJ_2_7_0 ( .G_IK(\PG_Network[2][1][63] ), .P_IK(
        \PG_Network[2][0][63] ), .G_K_1(n5), .P_K_1(\PG_Network[2][0][59] ), 
        .Gx(\PG_Network[3][1][63] ), .Px(\PG_Network[3][0][63] ) );
  G_14 GJ_3_0_0 ( .G_IK(\PG_Network[3][1][15] ), .P_IK(\PG_Network[3][0][15] ), 
        .G_K_1(Co[1]), .Gx(Co[3]) );
  G_13 GJ_3_0_1 ( .G_IK(\PG_Network[2][1][11] ), .P_IK(\PG_Network[2][0][11] ), 
        .G_K_1(Co[1]), .Gx(Co[2]) );
  PG_10 PGJ_3_1_0 ( .G_IK(\PG_Network[3][1][31] ), .P_IK(
        \PG_Network[3][0][31] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(
        \PG_Network[3][0][23] ), .Gx(\PG_Network[4][1][31] ), .Px(
        \PG_Network[4][0][31] ) );
  PG_9 PGJ_3_1_1 ( .G_IK(\PG_Network[2][1][27] ), .P_IK(\PG_Network[2][0][27] ), .G_K_1(\PG_Network[3][1][23] ), .P_K_1(\PG_Network[3][0][23] ), .Gx(
        \PG_Network[4][1][27] ), .Px(\PG_Network[4][0][27] ) );
  PG_8 PGJ_3_2_0 ( .G_IK(\PG_Network[3][1][47] ), .P_IK(\PG_Network[3][0][47] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(\PG_Network[3][0][39] ), .Gx(
        \PG_Network[4][1][47] ), .Px(\PG_Network[4][0][47] ) );
  PG_7 PGJ_3_2_1 ( .G_IK(\PG_Network[2][1][43] ), .P_IK(\PG_Network[2][0][43] ), .G_K_1(\PG_Network[3][1][39] ), .P_K_1(\PG_Network[3][0][39] ), .Gx(
        \PG_Network[4][1][43] ), .Px(\PG_Network[4][0][43] ) );
  PG_6 PGJ_3_3_0 ( .G_IK(\PG_Network[3][1][63] ), .P_IK(\PG_Network[3][0][63] ), .G_K_1(n7), .P_K_1(\PG_Network[3][0][55] ), .Gx(\PG_Network[4][1][63] ), 
        .Px(\PG_Network[4][0][63] ) );
  PG_5 PGJ_3_3_1 ( .G_IK(\PG_Network[2][1][59] ), .P_IK(\PG_Network[2][0][59] ), .G_K_1(\PG_Network[3][1][55] ), .P_K_1(\PG_Network[3][0][55] ), .Gx(
        \PG_Network[4][1][59] ), .Px(\PG_Network[4][0][59] ) );
  G_12 GJ_4_0_0 ( .G_IK(\PG_Network[4][1][31] ), .P_IK(\PG_Network[4][0][31] ), 
        .G_K_1(Co[3]), .Gx(Co[7]) );
  G_11 GJ_4_0_1 ( .G_IK(\PG_Network[4][1][27] ), .P_IK(\PG_Network[4][0][27] ), 
        .G_K_1(Co[3]), .Gx(Co[6]) );
  G_10 GJ_4_0_2 ( .G_IK(\PG_Network[3][1][23] ), .P_IK(\PG_Network[3][0][23] ), 
        .G_K_1(Co[3]), .Gx(Co[5]) );
  G_9 GJ_4_0_3 ( .G_IK(\PG_Network[2][1][19] ), .P_IK(\PG_Network[2][0][19] ), 
        .G_K_1(Co[3]), .Gx(Co[4]) );
  PG_4 PGJ_4_1_0 ( .G_IK(\PG_Network[4][1][63] ), .P_IK(\PG_Network[4][0][63] ), .G_K_1(n6), .P_K_1(\PG_Network[4][0][47] ), .Gx(\PG_Network[5][1][63] ), 
        .Px(\PG_Network[5][0][63] ) );
  PG_3 PGJ_4_1_1 ( .G_IK(\PG_Network[4][1][59] ), .P_IK(\PG_Network[4][0][59] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(\PG_Network[4][0][47] ), .Gx(
        \PG_Network[5][1][59] ), .Px(\PG_Network[5][0][59] ) );
  PG_2 PGJ_4_1_2 ( .G_IK(n7), .P_IK(\PG_Network[3][0][55] ), .G_K_1(
        \PG_Network[4][1][47] ), .P_K_1(\PG_Network[4][0][47] ), .Gx(
        \PG_Network[5][1][55] ), .Px(\PG_Network[5][0][55] ) );
  PG_1 PGJ_4_1_3 ( .G_IK(\PG_Network[2][1][51] ), .P_IK(\PG_Network[2][0][51] ), .G_K_1(\PG_Network[4][1][47] ), .P_K_1(\PG_Network[4][0][47] ), .Gx(
        \PG_Network[5][1][51] ), .Px(\PG_Network[5][0][51] ) );
  G_8 GJ_5_0_0 ( .G_IK(\PG_Network[5][1][63] ), .P_IK(\PG_Network[5][0][63] ), 
        .G_K_1(Co[7]), .Gx(Co[15]) );
  G_7 GJ_5_0_1 ( .G_IK(\PG_Network[5][1][59] ), .P_IK(\PG_Network[5][0][59] ), 
        .G_K_1(Co[7]), .Gx(Co[14]) );
  G_6 GJ_5_0_2 ( .G_IK(\PG_Network[5][1][55] ), .P_IK(\PG_Network[5][0][55] ), 
        .G_K_1(Co[7]), .Gx(Co[13]) );
  G_5 GJ_5_0_3 ( .G_IK(\PG_Network[5][1][51] ), .P_IK(\PG_Network[5][0][51] ), 
        .G_K_1(Co[7]), .Gx(Co[12]) );
  G_4 GJ_5_0_4 ( .G_IK(n6), .P_IK(\PG_Network[4][0][47] ), .G_K_1(Co[7]), .Gx(
        Co[11]) );
  G_3 GJ_5_0_5 ( .G_IK(\PG_Network[4][1][43] ), .P_IK(\PG_Network[4][0][43] ), 
        .G_K_1(Co[7]), .Gx(Co[10]) );
  G_2 GJ_5_0_6 ( .G_IK(\PG_Network[3][1][39] ), .P_IK(\PG_Network[3][0][39] ), 
        .G_K_1(Co[7]), .Gx(Co[9]) );
  G_1 GJ_5_0_7 ( .G_IK(\PG_Network[2][1][35] ), .P_IK(\PG_Network[2][0][35] ), 
        .G_K_1(Co[7]), .Gx(Co[8]) );
  CLKBUF_X1 U1 ( .A(\PG_Network[3][1][55] ), .Z(n7) );
  CLKBUF_X1 U2 ( .A(\PG_Network[2][1][59] ), .Z(n5) );
  INV_X1 U3 ( .A(A[53]), .ZN(n9) );
  INV_X1 U4 ( .A(A[47]), .ZN(n10) );
  INV_X1 U5 ( .A(A[43]), .ZN(n8) );
  INV_X1 U6 ( .A(A[57]), .ZN(n11) );
  INV_X1 U7 ( .A(A[55]), .ZN(n14) );
  INV_X1 U8 ( .A(A[51]), .ZN(n13) );
  INV_X1 U9 ( .A(A[59]), .ZN(n12) );
  CLKBUF_X1 U10 ( .A(\PG_Network[4][1][47] ), .Z(n6) );
  XNOR2_X1 U11 ( .A(B[43]), .B(n8), .ZN(\PG_Network[0][0][43] ) );
  XNOR2_X1 U12 ( .A(B[53]), .B(n9), .ZN(\PG_Network[0][0][53] ) );
  XNOR2_X1 U13 ( .A(B[47]), .B(n10), .ZN(\PG_Network[0][0][47] ) );
  XNOR2_X1 U14 ( .A(B[57]), .B(n11), .ZN(\PG_Network[0][0][57] ) );
  XNOR2_X1 U15 ( .A(B[59]), .B(n12), .ZN(\PG_Network[0][0][59] ) );
  XNOR2_X1 U16 ( .A(B[51]), .B(n13), .ZN(\PG_Network[0][0][51] ) );
  XNOR2_X1 U17 ( .A(B[55]), .B(n14), .ZN(\PG_Network[0][0][55] ) );
  AND2_X1 U18 ( .A1(A[46]), .A2(B[46]), .ZN(\PG_Network[0][1][46] ) );
  AND2_X1 U19 ( .A1(A[47]), .A2(B[47]), .ZN(\PG_Network[0][1][47] ) );
  AND2_X1 U20 ( .A1(A[44]), .A2(B[44]), .ZN(\PG_Network[0][1][44] ) );
  AND2_X1 U21 ( .A1(A[45]), .A2(B[45]), .ZN(\PG_Network[0][1][45] ) );
  AND2_X1 U22 ( .A1(A[58]), .A2(B[58]), .ZN(\PG_Network[0][1][58] ) );
  AND2_X1 U23 ( .A1(A[54]), .A2(B[54]), .ZN(\PG_Network[0][1][54] ) );
  AND2_X1 U24 ( .A1(B[55]), .A2(A[55]), .ZN(\PG_Network[0][1][55] ) );
  AND2_X1 U25 ( .A1(B[52]), .A2(A[52]), .ZN(\PG_Network[0][1][52] ) );
  AND2_X1 U26 ( .A1(A[53]), .A2(B[53]), .ZN(\PG_Network[0][1][53] ) );
  AND2_X1 U27 ( .A1(B[56]), .A2(A[56]), .ZN(\PG_Network[0][1][56] ) );
  AND2_X1 U28 ( .A1(B[57]), .A2(A[57]), .ZN(\PG_Network[0][1][57] ) );
  AND2_X1 U29 ( .A1(A[30]), .A2(B[30]), .ZN(\PG_Network[0][1][30] ) );
  AND2_X1 U30 ( .A1(A[31]), .A2(B[31]), .ZN(\PG_Network[0][1][31] ) );
  AND2_X1 U31 ( .A1(A[42]), .A2(B[42]), .ZN(\PG_Network[0][1][42] ) );
  AND2_X1 U32 ( .A1(B[43]), .A2(A[43]), .ZN(\PG_Network[0][1][43] ) );
  AND2_X1 U33 ( .A1(A[40]), .A2(B[40]), .ZN(\PG_Network[0][1][40] ) );
  AND2_X1 U34 ( .A1(A[41]), .A2(B[41]), .ZN(\PG_Network[0][1][41] ) );
  AND2_X1 U35 ( .A1(A[34]), .A2(B[34]), .ZN(\PG_Network[0][1][34] ) );
  AND2_X1 U36 ( .A1(A[35]), .A2(B[35]), .ZN(\PG_Network[0][1][35] ) );
  AND2_X1 U37 ( .A1(A[33]), .A2(B[33]), .ZN(\PG_Network[0][1][33] ) );
  AND2_X1 U38 ( .A1(A[32]), .A2(B[32]), .ZN(\PG_Network[0][1][32] ) );
  AND2_X1 U39 ( .A1(A[50]), .A2(B[50]), .ZN(\PG_Network[0][1][50] ) );
  AND2_X1 U40 ( .A1(B[51]), .A2(A[51]), .ZN(\PG_Network[0][1][51] ) );
  AND2_X1 U41 ( .A1(A[48]), .A2(B[48]), .ZN(\PG_Network[0][1][48] ) );
  AND2_X1 U42 ( .A1(A[49]), .A2(B[49]), .ZN(\PG_Network[0][1][49] ) );
  AND2_X1 U43 ( .A1(A[36]), .A2(B[36]), .ZN(\PG_Network[0][1][36] ) );
  AND2_X1 U44 ( .A1(A[37]), .A2(B[37]), .ZN(\PG_Network[0][1][37] ) );
  AND2_X1 U45 ( .A1(A[38]), .A2(B[38]), .ZN(\PG_Network[0][1][38] ) );
  AND2_X1 U46 ( .A1(A[39]), .A2(B[39]), .ZN(\PG_Network[0][1][39] ) );
  AND2_X1 U47 ( .A1(A[62]), .A2(B[62]), .ZN(\PG_Network[0][1][62] ) );
  AND2_X1 U48 ( .A1(A[17]), .A2(B[17]), .ZN(\PG_Network[0][1][17] ) );
  AND2_X1 U49 ( .A1(A[16]), .A2(B[16]), .ZN(\PG_Network[0][1][16] ) );
  AND2_X1 U50 ( .A1(A[19]), .A2(B[19]), .ZN(\PG_Network[0][1][19] ) );
  AND2_X1 U51 ( .A1(A[18]), .A2(B[18]), .ZN(\PG_Network[0][1][18] ) );
  AND2_X1 U52 ( .A1(A[9]), .A2(B[9]), .ZN(\PG_Network[0][1][9] ) );
  AND2_X1 U53 ( .A1(A[8]), .A2(B[8]), .ZN(\PG_Network[0][1][8] ) );
  AND2_X1 U54 ( .A1(A[11]), .A2(B[11]), .ZN(\PG_Network[0][1][11] ) );
  AND2_X1 U55 ( .A1(A[10]), .A2(B[10]), .ZN(\PG_Network[0][1][10] ) );
  AND2_X1 U56 ( .A1(A[15]), .A2(B[15]), .ZN(\PG_Network[0][1][15] ) );
  AND2_X1 U57 ( .A1(A[14]), .A2(B[14]), .ZN(\PG_Network[0][1][14] ) );
  AND2_X1 U58 ( .A1(A[25]), .A2(B[25]), .ZN(\PG_Network[0][1][25] ) );
  AND2_X1 U59 ( .A1(A[24]), .A2(B[24]), .ZN(\PG_Network[0][1][24] ) );
  AND2_X1 U60 ( .A1(A[27]), .A2(B[27]), .ZN(\PG_Network[0][1][27] ) );
  AND2_X1 U61 ( .A1(A[26]), .A2(B[26]), .ZN(\PG_Network[0][1][26] ) );
  AND2_X1 U62 ( .A1(A[61]), .A2(B[61]), .ZN(\PG_Network[0][1][61] ) );
  AND2_X1 U63 ( .A1(A[5]), .A2(B[5]), .ZN(\PG_Network[0][1][5] ) );
  AND2_X1 U64 ( .A1(A[4]), .A2(B[4]), .ZN(\PG_Network[0][1][4] ) );
  AND2_X1 U65 ( .A1(A[3]), .A2(B[3]), .ZN(\PG_Network[0][1][3] ) );
  AND2_X1 U66 ( .A1(A[2]), .A2(B[2]), .ZN(\PG_Network[0][1][2] ) );
  INV_X1 U67 ( .A(n18), .ZN(n15) );
  AND2_X1 U77 ( .A1(A[1]), .A2(B[1]), .ZN(\PG_Network[0][1][1] ) );
  AND2_X1 U79 ( .A1(A[28]), .A2(B[28]), .ZN(\PG_Network[0][1][28] ) );
  AND2_X1 U81 ( .A1(A[6]), .A2(B[6]), .ZN(\PG_Network[0][1][6] ) );
  AND2_X1 U83 ( .A1(A[29]), .A2(B[29]), .ZN(\PG_Network[0][1][29] ) );
  AND2_X1 U85 ( .A1(A[7]), .A2(B[7]), .ZN(\PG_Network[0][1][7] ) );
  AND2_X1 U90 ( .A1(A[21]), .A2(B[21]), .ZN(\PG_Network[0][1][21] ) );
  AND2_X1 U94 ( .A1(A[20]), .A2(B[20]), .ZN(\PG_Network[0][1][20] ) );
  AND2_X1 U131 ( .A1(A[13]), .A2(B[13]), .ZN(\PG_Network[0][1][13] ) );
  AND2_X1 U132 ( .A1(A[12]), .A2(B[12]), .ZN(\PG_Network[0][1][12] ) );
  AND2_X1 U133 ( .A1(A[23]), .A2(B[23]), .ZN(\PG_Network[0][1][23] ) );
  AND2_X1 U134 ( .A1(A[22]), .A2(B[22]), .ZN(\PG_Network[0][1][22] ) );
  AOI21_X1 U135 ( .B1(A[0]), .B2(B[0]), .A(n16), .ZN(n18) );
  INV_X1 U136 ( .A(n17), .ZN(n16) );
  OAI21_X1 U137 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n17) );
  AND2_X1 U138 ( .A1(A[63]), .A2(B[63]), .ZN(\PG_Network[0][1][63] ) );
  AND2_X1 U139 ( .A1(A[60]), .A2(B[60]), .ZN(\PG_Network[0][1][60] ) );
  AND2_X1 U140 ( .A1(B[59]), .A2(A[59]), .ZN(\PG_Network[0][1][59] ) );
endmodule


module FA_128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_32 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_128 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_127 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_126 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_125 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_123 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_122 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_121 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_31 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_124 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_123 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_122 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_121 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_16 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U2 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U4 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U5 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U7 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U9 ( .A(sel), .ZN(n13) );
endmodule


module carry_select_block_NPB4_16 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_32 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_31 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_16 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_30 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_120 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_119 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_118 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_117 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_29 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_116 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_115 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_114 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_113 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_15 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_15 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_30 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_29 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_15 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_28 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_112 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_111 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_110 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_109 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_27 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_108 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_107 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_106 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_105 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_14 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_14 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_28 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_27 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_14 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_26 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_104 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_103 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_102 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_101 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_25 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_100 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_99 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_98 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_97 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_13 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_13 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_26 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_25 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_13 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_24 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_96 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_95 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_94 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_93 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_23 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_92 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_91 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_90 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_89 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_12 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_12 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_24 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_23 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_12 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_22 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_88 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_87 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_86 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_85 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_21 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_84 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_83 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_82 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_81 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_11 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_11 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_22 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_21 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_11 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_20 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_80 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_79 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_78 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_77 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_19 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_76 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_75 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_74 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_73 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_10 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_10 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_20 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_19 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_10 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_18 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_72 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_71 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_70 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_69 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_17 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_68 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_67 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_66 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_65 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_9 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_9 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_18 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_17 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_9 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_16 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_64 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_8 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_8 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_16 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_15 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_8 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_7 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_14 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_13 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_7 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_6 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_12 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_11 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_6 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_5 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_10 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_9 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_5 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_4 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n13), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[3]), .B1(B[3]), .B2(n13), .ZN(n17) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n13), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n13), .ZN(n14) );
endmodule


module carry_select_block_NPB4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_8 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_7 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_4 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_3 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  BUF_X1 U1 ( .A(sel), .Z(n5) );
  INV_X1 U2 ( .A(sel), .ZN(n14) );
  INV_X1 U3 ( .A(n17), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n14), .ZN(n17) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U6 ( .A(n16), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n5), .B1(B[1]), .B2(n14), .ZN(n16) );
  INV_X1 U8 ( .A(n15), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(n5), .A2(A[0]), .B1(B[0]), .B2(n14), .ZN(n15) );
  AOI22_X1 U10 ( .A1(n5), .A2(A[3]), .B1(B[3]), .B2(n14), .ZN(n18) );
endmodule


module carry_select_block_NPB4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_6 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_5 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_3 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_2 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(sel), .ZN(n5) );
  INV_X1 U2 ( .A(sel), .ZN(n14) );
  INV_X1 U3 ( .A(n17), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(sel), .B1(B[2]), .B2(n14), .ZN(n17) );
  INV_X1 U5 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U6 ( .A(n16), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(sel), .B1(B[1]), .B2(n14), .ZN(n16) );
  INV_X1 U8 ( .A(n15), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(sel), .B1(B[0]), .B2(n5), .ZN(n15) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n5), .ZN(n18) );
endmodule


module carry_select_block_NPB4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_4 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_3 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_2 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net67632, n4, n5, n6, n7, n8;
  assign Co = net67632;

  INV_X1 U1 ( .A(Ci), .ZN(n8) );
  AND2_X1 U2 ( .A1(n7), .A2(n8), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
  XNOR2_X1 U6 ( .A(Ci), .B(n5), .ZN(S) );
  AOI21_X1 U7 ( .B1(n6), .B2(n7), .A(n4), .ZN(net67632) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n7, n8;

  XOR2_X1 U3 ( .A(n4), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n4) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n5) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n7), .ZN(n8) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(n4), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module RCA_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6, n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n8), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n6) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  CLKBUF_X1 U4 ( .A(n8), .Z(n5) );
  XNOR2_X1 U5 ( .A(B), .B(n6), .ZN(n8) );
  INV_X1 U6 ( .A(n9), .ZN(Co) );
  AOI22_X1 U7 ( .A1(n4), .A2(A), .B1(n5), .B2(Ci), .ZN(n9) );
endmodule


module RCA_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_generic_N4_1 ( A, B, sel, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input sel;
  wire   n5, n14, n15, n16, n17, n18;

  INV_X1 U1 ( .A(sel), .ZN(n5) );
  INV_X1 U2 ( .A(n15), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n18), .ZN(Y[3]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(sel), .A2(A[2]), .B1(n5), .B2(B[2]), .ZN(n17) );
  AOI22_X1 U6 ( .A1(sel), .A2(A[0]), .B1(n5), .B2(B[0]), .ZN(n15) );
  AOI22_X1 U7 ( .A1(sel), .A2(A[1]), .B1(n14), .B2(B[1]), .ZN(n16) );
  INV_X1 U8 ( .A(sel), .ZN(n14) );
  INV_X1 U9 ( .A(n17), .ZN(Y[2]) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(sel), .B1(B[3]), .B2(n14), .ZN(n18) );
endmodule


module carry_select_block_NPB4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_N4_2 UADDER1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  RCA_N4_1 UADDER2 ( .A(A), .B(B), .Ci(1'b0), .S(S2) );
  MUX21_generic_N4_1 mux ( .A(S1), .B(S2), .sel(Ci), .Y(S) );
endmodule


module sum_generator_N64_NPB4_1 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  input [16:0] Ci;
  output [63:0] S;
  output Co;

  assign Co = Ci[16];

  carry_select_block_NPB4_16 csbi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(
        S[3:0]) );
  carry_select_block_NPB4_15 csbi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(
        S[7:4]) );
  carry_select_block_NPB4_14 csbi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), 
        .S(S[11:8]) );
  carry_select_block_NPB4_13 csbi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), 
        .S(S[15:12]) );
  carry_select_block_NPB4_12 csbi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), 
        .S(S[19:16]) );
  carry_select_block_NPB4_11 csbi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), 
        .S(S[23:20]) );
  carry_select_block_NPB4_10 csbi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), 
        .S(S[27:24]) );
  carry_select_block_NPB4_9 csbi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), 
        .S(S[31:28]) );
  carry_select_block_NPB4_8 csbi_8 ( .A(A[35:32]), .B(B[35:32]), .Ci(Ci[8]), 
        .S(S[35:32]) );
  carry_select_block_NPB4_7 csbi_9 ( .A(A[39:36]), .B(B[39:36]), .Ci(Ci[9]), 
        .S(S[39:36]) );
  carry_select_block_NPB4_6 csbi_10 ( .A(A[43:40]), .B(B[43:40]), .Ci(Ci[10]), 
        .S(S[43:40]) );
  carry_select_block_NPB4_5 csbi_11 ( .A(A[47:44]), .B(B[47:44]), .Ci(Ci[11]), 
        .S(S[47:44]) );
  carry_select_block_NPB4_4 csbi_12 ( .A(A[51:48]), .B(B[51:48]), .Ci(Ci[12]), 
        .S(S[51:48]) );
  carry_select_block_NPB4_3 csbi_13 ( .A(A[55:52]), .B(B[55:52]), .Ci(Ci[13]), 
        .S(S[55:52]) );
  carry_select_block_NPB4_2 csbi_14 ( .A(A[59:56]), .B(B[59:56]), .Ci(Ci[14]), 
        .S(S[59:56]) );
  carry_select_block_NPB4_1 csbi_15 ( .A(A[63:60]), .B(B[63:60]), .Ci(Ci[15]), 
        .S(S[63:60]) );
endmodule


module P4_ADDER_N64_1 ( A, B, Cin, S, Cout );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [16:1] CoutCgen;

  carry_generator_N64_NPB4_1 CGEN ( .A(A), .B({B[63], n2, n13, n14, B[59:0]}), 
        .Cin(Cin), .Co(CoutCgen) );
  sum_generator_N64_NPB4_1 SGEN ( .A(A), .B({B[63:60], n10, n8, n12, B[56], 
        n11, n3, n7, B[52], n9, B[50], n6, B[48], n5, B[46], n4, B[44], n1, 
        B[42:0]}), .Ci({CoutCgen, Cin}), .S(S), .Co(Cout) );
  CLKBUF_X1 U1 ( .A(B[43]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(B[62]), .Z(n2) );
  CLKBUF_X1 U3 ( .A(B[57]), .Z(n12) );
  CLKBUF_X1 U4 ( .A(B[54]), .Z(n3) );
  CLKBUF_X1 U5 ( .A(B[45]), .Z(n4) );
  CLKBUF_X1 U6 ( .A(B[47]), .Z(n5) );
  CLKBUF_X1 U7 ( .A(B[49]), .Z(n6) );
  CLKBUF_X1 U8 ( .A(B[53]), .Z(n7) );
  CLKBUF_X1 U9 ( .A(B[58]), .Z(n8) );
  CLKBUF_X1 U10 ( .A(B[51]), .Z(n9) );
  CLKBUF_X1 U11 ( .A(B[59]), .Z(n10) );
  CLKBUF_X1 U12 ( .A(B[55]), .Z(n11) );
  CLKBUF_X1 U13 ( .A(B[61]), .Z(n13) );
  CLKBUF_X1 U14 ( .A(B[60]), .Z(n14) );
endmodule


module booth_mul_N32_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n98, n99, n101, n102, n103, n106, n107, n109, n110, n111,
         n114, n117, n118, n121, n123, n125, n127, n128, n96, n97, n100, n104,
         n105, n108, n112, n113, n115, n116, n119, n120, n122, n124, n126,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U44 ( .A(n101), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U45 ( .A(n103), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U51 ( .A(n111), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U56 ( .A(n117), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U59 ( .A(n121), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U60 ( .A(n123), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U62 ( .A(n140), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U63 ( .A(n127), .B(B[3]), .Z(DIFF[3]) );
  OR2_X1 U1 ( .A1(n153), .A2(n158), .ZN(n160) );
  OR3_X1 U2 ( .A1(n137), .A2(B[4]), .A3(B[3]), .ZN(n140) );
  OR3_X1 U3 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n137) );
  OR2_X1 U4 ( .A1(n113), .A2(n133), .ZN(n121) );
  NAND2_X1 U5 ( .A1(n124), .A2(n126), .ZN(DIFF[21]) );
  INV_X1 U6 ( .A(n139), .ZN(n96) );
  NAND2_X1 U7 ( .A1(n138), .A2(n97), .ZN(n98) );
  NOR2_X1 U8 ( .A1(n152), .A2(n96), .ZN(n97) );
  NAND2_X1 U9 ( .A1(n130), .A2(n131), .ZN(n100) );
  OR2_X1 U10 ( .A1(n100), .A2(n104), .ZN(n103) );
  OR2_X1 U11 ( .A1(n105), .A2(n166), .ZN(n104) );
  INV_X1 U12 ( .A(n115), .ZN(n105) );
  OR2_X1 U13 ( .A1(n132), .A2(n155), .ZN(n108) );
  OR2_X1 U14 ( .A1(n132), .A2(n155), .ZN(n123) );
  NOR2_X1 U15 ( .A1(n132), .A2(n112), .ZN(n146) );
  OR2_X1 U16 ( .A1(n155), .A2(B[7]), .ZN(n112) );
  OR3_X1 U17 ( .A1(n136), .A2(B[4]), .A3(B[3]), .ZN(n113) );
  NOR2_X1 U18 ( .A1(B[25]), .A2(B[26]), .ZN(n115) );
  NOR2_X1 U19 ( .A1(B[27]), .A2(B[28]), .ZN(n116) );
  XNOR2_X1 U20 ( .A(n119), .B(B[11]), .ZN(DIFF[11]) );
  NOR2_X1 U21 ( .A1(n134), .A2(n147), .ZN(n119) );
  NAND2_X1 U22 ( .A1(n109), .A2(n122), .ZN(n124) );
  NAND2_X1 U23 ( .A1(n120), .A2(B[21]), .ZN(n126) );
  INV_X1 U24 ( .A(n109), .ZN(n120) );
  INV_X1 U25 ( .A(B[21]), .ZN(n122) );
  OR3_X2 U26 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n127) );
  XNOR2_X1 U27 ( .A(n129), .B(B[15]), .ZN(DIFF[15]) );
  NOR2_X1 U28 ( .A1(n108), .A2(n160), .ZN(n129) );
  NAND2_X1 U29 ( .A1(n130), .A2(n131), .ZN(n107) );
  NOR2_X1 U30 ( .A1(n145), .A2(n148), .ZN(n130) );
  NOR2_X1 U31 ( .A1(n161), .A2(n165), .ZN(n131) );
  OR2_X2 U32 ( .A1(B[7]), .A2(B[8]), .ZN(n163) );
  OR3_X2 U33 ( .A1(n141), .A2(B[4]), .A3(B[3]), .ZN(n125) );
  OR3_X2 U34 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n136) );
  OR3_X2 U35 ( .A1(n136), .A2(B[4]), .A3(B[3]), .ZN(n132) );
  OR2_X2 U36 ( .A1(n125), .A2(n155), .ZN(n134) );
  XNOR2_X1 U37 ( .A(n143), .B(B[6]), .ZN(DIFF[6]) );
  OR2_X1 U38 ( .A1(n155), .A2(n163), .ZN(n133) );
  NOR2_X1 U39 ( .A1(n108), .A2(n135), .ZN(n118) );
  OR2_X1 U40 ( .A1(n147), .A2(B[11]), .ZN(n135) );
  NOR2_X1 U41 ( .A1(n107), .A2(n166), .ZN(n138) );
  NAND2_X1 U42 ( .A1(n138), .A2(n139), .ZN(n101) );
  AND2_X1 U43 ( .A1(n116), .A2(n115), .ZN(n139) );
  OR2_X2 U46 ( .A1(n134), .A2(n160), .ZN(n145) );
  OR3_X2 U47 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n141) );
  XNOR2_X1 U48 ( .A(n142), .B(B[17]), .ZN(DIFF[17]) );
  NOR2_X1 U49 ( .A1(n144), .A2(n167), .ZN(n142) );
  NOR2_X1 U50 ( .A1(n140), .A2(B[5]), .ZN(n143) );
  OR2_X1 U52 ( .A1(n134), .A2(n160), .ZN(n144) );
  XNOR2_X1 U53 ( .A(n146), .B(B[8]), .ZN(DIFF[8]) );
  OR2_X1 U54 ( .A1(n168), .A2(n163), .ZN(n147) );
  OR2_X1 U55 ( .A1(n154), .A2(n167), .ZN(n148) );
  XNOR2_X1 U57 ( .A(n149), .B(B[25]), .ZN(DIFF[25]) );
  NOR2_X1 U58 ( .A1(n166), .A2(n107), .ZN(n149) );
  OR2_X1 U61 ( .A1(n166), .A2(n107), .ZN(n150) );
  XNOR2_X1 U64 ( .A(n151), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U65 ( .A1(n121), .A2(B[9]), .ZN(n151) );
  OR2_X1 U66 ( .A1(B[29]), .A2(B[30]), .ZN(n152) );
  INV_X1 U67 ( .A(B[23]), .ZN(n159) );
  OR2_X1 U68 ( .A1(n168), .A2(n169), .ZN(n153) );
  OR2_X1 U69 ( .A1(B[17]), .A2(B[18]), .ZN(n154) );
  OR2_X2 U70 ( .A1(n145), .A2(n148), .ZN(n111) );
  OR2_X1 U71 ( .A1(B[5]), .A2(B[6]), .ZN(n155) );
  OR2_X1 U72 ( .A1(n167), .A2(n145), .ZN(n156) );
  AND2_X1 U73 ( .A1(n98), .A2(n176), .ZN(DIFF[32]) );
  OR2_X1 U74 ( .A1(n163), .A2(n164), .ZN(n158) );
  OR2_X1 U75 ( .A1(n162), .A2(n134), .ZN(n117) );
  XNOR2_X1 U76 ( .A(n107), .B(n159), .ZN(DIFF[23]) );
  OR2_X2 U77 ( .A1(n111), .A2(n165), .ZN(n109) );
  OR2_X1 U78 ( .A1(B[21]), .A2(B[22]), .ZN(n161) );
  OR2_X1 U79 ( .A1(n163), .A2(n153), .ZN(n162) );
  OR2_X1 U80 ( .A1(B[14]), .A2(B[13]), .ZN(n164) );
  OR2_X1 U81 ( .A1(B[19]), .A2(B[20]), .ZN(n165) );
  OR2_X1 U82 ( .A1(B[23]), .A2(B[24]), .ZN(n166) );
  OR2_X1 U83 ( .A1(B[15]), .A2(B[16]), .ZN(n167) );
  OR2_X1 U84 ( .A1(B[10]), .A2(B[9]), .ZN(n168) );
  OR2_X1 U85 ( .A1(B[12]), .A2(B[11]), .ZN(n169) );
  XOR2_X1 U86 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XNOR2_X1 U87 ( .A(n170), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U88 ( .A1(n150), .A2(B[25]), .ZN(n170) );
  XNOR2_X1 U89 ( .A(n171), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U90 ( .A1(n101), .A2(B[29]), .ZN(n171) );
  XNOR2_X1 U91 ( .A(n110), .B(B[20]), .ZN(DIFF[20]) );
  XNOR2_X1 U92 ( .A(B[24]), .B(n106), .ZN(DIFF[24]) );
  XNOR2_X1 U93 ( .A(n172), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U94 ( .A1(n109), .A2(B[21]), .ZN(n172) );
  XOR2_X1 U95 ( .A(B[4]), .B(n173), .Z(DIFF[4]) );
  OR2_X1 U96 ( .A1(n127), .A2(B[3]), .ZN(n173) );
  XNOR2_X1 U97 ( .A(n174), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U98 ( .A1(n117), .A2(B[13]), .ZN(n174) );
  XNOR2_X1 U99 ( .A(n175), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U100 ( .A1(n156), .A2(B[17]), .ZN(n175) );
  XNOR2_X1 U101 ( .A(n118), .B(B[12]), .ZN(DIFF[12]) );
  XNOR2_X1 U102 ( .A(B[16]), .B(n114), .ZN(DIFF[16]) );
  XNOR2_X1 U103 ( .A(n102), .B(B[28]), .ZN(DIFF[28]) );
  NOR2_X1 U104 ( .A1(B[27]), .A2(n103), .ZN(n102) );
  NOR2_X1 U105 ( .A1(\B[0] ), .A2(B[1]), .ZN(n128) );
  NOR2_X1 U106 ( .A1(B[15]), .A2(n144), .ZN(n114) );
  NOR2_X1 U107 ( .A1(B[23]), .A2(n107), .ZN(n106) );
  NOR2_X1 U108 ( .A1(B[19]), .A2(n111), .ZN(n110) );
  XNOR2_X1 U109 ( .A(B[2]), .B(n128), .ZN(DIFF[2]) );
  NAND2_X1 U110 ( .A1(n98), .A2(n176), .ZN(n99) );
  OAI21_X1 U111 ( .B1(n98), .B2(n176), .A(n99), .ZN(DIFF[31]) );
  INV_X1 U112 ( .A(B[32]), .ZN(n176) );
endmodule


module booth_mul_N32 ( A, B, S );
  input [31:0] A;
  input [31:0] B;
  output [63:0] S;
  wire   minus_A_63, \select_array[15][2] , \select_array[15][1] ,
         \select_array[15][0] , \select_array[14][2] , \select_array[14][1] ,
         \select_array[14][0] , \select_array[13][2] , \select_array[13][1] ,
         \select_array[13][0] , \select_array[12][2] , \select_array[12][1] ,
         \select_array[12][0] , \select_array[11][2] , \select_array[11][1] ,
         \select_array[11][0] , \select_array[10][2] , \select_array[10][1] ,
         \select_array[10][0] , \select_array[9][2] , \select_array[9][1] ,
         \select_array[9][0] , \select_array[8][2] , \select_array[8][1] ,
         \select_array[8][0] , \select_array[7][2] , \select_array[7][1] ,
         \select_array[7][0] , \select_array[6][2] , \select_array[6][1] ,
         \select_array[6][0] , \select_array[5][2] , \select_array[5][1] ,
         \select_array[5][0] , \select_array[4][2] , \select_array[4][1] ,
         \select_array[4][0] , \select_array[3][2] , \select_array[3][1] ,
         \select_array[3][0] , \select_array[2][2] , \select_array[2][1] ,
         \select_array[2][0] , \select_array[1][2] , \select_array[1][1] ,
         \select_array[1][0] , \select_array[0][2] , \select_array[0][1] ,
         \select_array[0][0] , \result_array[7][63] , \result_array[7][62] ,
         \result_array[7][61] , \result_array[7][60] , \result_array[7][59] ,
         \result_array[7][58] , \result_array[7][57] , \result_array[7][56] ,
         \result_array[7][55] , \result_array[7][54] , \result_array[7][53] ,
         \result_array[7][52] , \result_array[7][51] , \result_array[7][50] ,
         \result_array[7][49] , \result_array[7][48] , \result_array[7][47] ,
         \result_array[7][46] , \result_array[7][45] , \result_array[7][44] ,
         \result_array[7][43] , \result_array[7][42] , \result_array[7][41] ,
         \result_array[7][40] , \result_array[7][39] , \result_array[7][38] ,
         \result_array[7][37] , \result_array[7][36] , \result_array[7][35] ,
         \result_array[7][34] , \result_array[7][33] , \result_array[7][32] ,
         \result_array[7][31] , \result_array[7][30] , \result_array[7][29] ,
         \result_array[7][28] , \result_array[7][27] , \result_array[7][26] ,
         \result_array[7][25] , \result_array[7][24] , \result_array[7][23] ,
         \result_array[7][22] , \result_array[7][21] , \result_array[7][20] ,
         \result_array[7][19] , \result_array[7][18] , \result_array[7][17] ,
         \result_array[7][16] , \result_array[7][15] , \result_array[7][14] ,
         \result_array[7][13] , \result_array[7][12] , \result_array[7][11] ,
         \result_array[7][10] , \result_array[7][9] , \result_array[7][8] ,
         \result_array[7][7] , \result_array[7][6] , \result_array[7][5] ,
         \result_array[7][4] , \result_array[7][3] , \result_array[7][2] ,
         \result_array[7][1] , \result_array[7][0] , \result_array[6][63] ,
         \result_array[6][62] , \result_array[6][61] , \result_array[6][60] ,
         \result_array[6][59] , \result_array[6][58] , \result_array[6][57] ,
         \result_array[6][56] , \result_array[6][55] , \result_array[6][54] ,
         \result_array[6][53] , \result_array[6][52] , \result_array[6][51] ,
         \result_array[6][50] , \result_array[6][49] , \result_array[6][48] ,
         \result_array[6][47] , \result_array[6][46] , \result_array[6][45] ,
         \result_array[6][44] , \result_array[6][43] , \result_array[6][42] ,
         \result_array[6][41] , \result_array[6][40] , \result_array[6][39] ,
         \result_array[6][38] , \result_array[6][37] , \result_array[6][36] ,
         \result_array[6][35] , \result_array[6][34] , \result_array[6][33] ,
         \result_array[6][32] , \result_array[6][31] , \result_array[6][30] ,
         \result_array[6][29] , \result_array[6][28] , \result_array[6][27] ,
         \result_array[6][26] , \result_array[6][25] , \result_array[6][24] ,
         \result_array[6][23] , \result_array[6][22] , \result_array[6][21] ,
         \result_array[6][20] , \result_array[6][19] , \result_array[6][18] ,
         \result_array[6][17] , \result_array[6][16] , \result_array[6][15] ,
         \result_array[6][14] , \result_array[6][13] , \result_array[6][12] ,
         \result_array[6][11] , \result_array[6][10] , \result_array[6][9] ,
         \result_array[6][8] , \result_array[6][7] , \result_array[6][6] ,
         \result_array[6][5] , \result_array[6][4] , \result_array[6][3] ,
         \result_array[6][2] , \result_array[6][1] , \result_array[6][0] ,
         \result_array[5][63] , \result_array[5][62] , \result_array[5][61] ,
         \result_array[5][60] , \result_array[5][59] , \result_array[5][58] ,
         \result_array[5][57] , \result_array[5][56] , \result_array[5][55] ,
         \result_array[5][54] , \result_array[5][53] , \result_array[5][52] ,
         \result_array[5][51] , \result_array[5][50] , \result_array[5][49] ,
         \result_array[5][48] , \result_array[5][47] , \result_array[5][46] ,
         \result_array[5][45] , \result_array[5][44] , \result_array[5][43] ,
         \result_array[5][42] , \result_array[5][41] , \result_array[5][40] ,
         \result_array[5][39] , \result_array[5][38] , \result_array[5][37] ,
         \result_array[5][36] , \result_array[5][35] , \result_array[5][34] ,
         \result_array[5][33] , \result_array[5][32] , \result_array[5][31] ,
         \result_array[5][30] , \result_array[5][29] , \result_array[5][28] ,
         \result_array[5][27] , \result_array[5][26] , \result_array[5][25] ,
         \result_array[5][24] , \result_array[5][23] , \result_array[5][22] ,
         \result_array[5][21] , \result_array[5][20] , \result_array[5][19] ,
         \result_array[5][18] , \result_array[5][17] , \result_array[5][16] ,
         \result_array[5][15] , \result_array[5][14] , \result_array[5][13] ,
         \result_array[5][12] , \result_array[5][11] , \result_array[5][10] ,
         \result_array[5][9] , \result_array[5][8] , \result_array[5][7] ,
         \result_array[5][6] , \result_array[5][5] , \result_array[5][4] ,
         \result_array[5][3] , \result_array[5][2] , \result_array[5][1] ,
         \result_array[5][0] , \result_array[4][63] , \result_array[4][62] ,
         \result_array[4][61] , \result_array[4][60] , \result_array[4][59] ,
         \result_array[4][58] , \result_array[4][57] , \result_array[4][56] ,
         \result_array[4][55] , \result_array[4][54] , \result_array[4][53] ,
         \result_array[4][52] , \result_array[4][51] , \result_array[4][50] ,
         \result_array[4][49] , \result_array[4][48] , \result_array[4][47] ,
         \result_array[4][46] , \result_array[4][45] , \result_array[4][44] ,
         \result_array[4][43] , \result_array[4][42] , \result_array[4][41] ,
         \result_array[4][40] , \result_array[4][39] , \result_array[4][38] ,
         \result_array[4][37] , \result_array[4][36] , \result_array[4][35] ,
         \result_array[4][34] , \result_array[4][33] , \result_array[4][32] ,
         \result_array[4][31] , \result_array[4][30] , \result_array[4][29] ,
         \result_array[4][28] , \result_array[4][27] , \result_array[4][26] ,
         \result_array[4][25] , \result_array[4][24] , \result_array[4][23] ,
         \result_array[4][22] , \result_array[4][21] , \result_array[4][20] ,
         \result_array[4][19] , \result_array[4][18] , \result_array[4][17] ,
         \result_array[4][16] , \result_array[4][15] , \result_array[4][14] ,
         \result_array[4][13] , \result_array[4][12] , \result_array[4][11] ,
         \result_array[4][10] , \result_array[4][9] , \result_array[4][8] ,
         \result_array[4][7] , \result_array[4][6] , \result_array[4][5] ,
         \result_array[4][4] , \result_array[4][3] , \result_array[4][2] ,
         \result_array[4][1] , \result_array[4][0] , \result_array[3][63] ,
         \result_array[3][62] , \result_array[3][61] , \result_array[3][60] ,
         \result_array[3][59] , \result_array[3][58] , \result_array[3][57] ,
         \result_array[3][56] , \result_array[3][55] , \result_array[3][54] ,
         \result_array[3][53] , \result_array[3][52] , \result_array[3][51] ,
         \result_array[3][50] , \result_array[3][49] , \result_array[3][48] ,
         \result_array[3][47] , \result_array[3][46] , \result_array[3][45] ,
         \result_array[3][44] , \result_array[3][43] , \result_array[3][42] ,
         \result_array[3][41] , \result_array[3][40] , \result_array[3][39] ,
         \result_array[3][38] , \result_array[3][37] , \result_array[3][36] ,
         \result_array[3][35] , \result_array[3][34] , \result_array[3][33] ,
         \result_array[3][32] , \result_array[3][31] , \result_array[3][30] ,
         \result_array[3][29] , \result_array[3][28] , \result_array[3][27] ,
         \result_array[3][26] , \result_array[3][25] , \result_array[3][24] ,
         \result_array[3][23] , \result_array[3][22] , \result_array[3][21] ,
         \result_array[3][20] , \result_array[3][19] , \result_array[3][18] ,
         \result_array[3][17] , \result_array[3][16] , \result_array[3][15] ,
         \result_array[3][14] , \result_array[3][13] , \result_array[3][12] ,
         \result_array[3][11] , \result_array[3][10] , \result_array[3][9] ,
         \result_array[3][8] , \result_array[3][7] , \result_array[3][6] ,
         \result_array[3][5] , \result_array[3][4] , \result_array[3][3] ,
         \result_array[3][2] , \result_array[3][1] , \result_array[3][0] ,
         \result_array[2][63] , \result_array[2][62] , \result_array[2][61] ,
         \result_array[2][60] , \result_array[2][59] , \result_array[2][58] ,
         \result_array[2][57] , \result_array[2][56] , \result_array[2][55] ,
         \result_array[2][54] , \result_array[2][53] , \result_array[2][52] ,
         \result_array[2][51] , \result_array[2][50] , \result_array[2][49] ,
         \result_array[2][48] , \result_array[2][47] , \result_array[2][46] ,
         \result_array[2][45] , \result_array[2][44] , \result_array[2][43] ,
         \result_array[2][42] , \result_array[2][41] , \result_array[2][40] ,
         \result_array[2][39] , \result_array[2][38] , \result_array[2][37] ,
         \result_array[2][36] , \result_array[2][35] , \result_array[2][34] ,
         \result_array[2][33] , \result_array[2][32] , \result_array[2][31] ,
         \result_array[2][30] , \result_array[2][29] , \result_array[2][28] ,
         \result_array[2][27] , \result_array[2][26] , \result_array[2][25] ,
         \result_array[2][24] , \result_array[2][23] , \result_array[2][22] ,
         \result_array[2][21] , \result_array[2][20] , \result_array[2][19] ,
         \result_array[2][18] , \result_array[2][17] , \result_array[2][16] ,
         \result_array[2][15] , \result_array[2][14] , \result_array[2][13] ,
         \result_array[2][12] , \result_array[2][11] , \result_array[2][10] ,
         \result_array[2][9] , \result_array[2][8] , \result_array[2][7] ,
         \result_array[2][6] , \result_array[2][5] , \result_array[2][4] ,
         \result_array[2][3] , \result_array[2][2] , \result_array[2][1] ,
         \result_array[2][0] , \result_array[1][63] , \result_array[1][62] ,
         \result_array[1][61] , \result_array[1][60] , \result_array[1][59] ,
         \result_array[1][58] , \result_array[1][57] , \result_array[1][56] ,
         \result_array[1][55] , \result_array[1][54] , \result_array[1][53] ,
         \result_array[1][52] , \result_array[1][51] , \result_array[1][50] ,
         \result_array[1][49] , \result_array[1][48] , \result_array[1][47] ,
         \result_array[1][46] , \result_array[1][45] , \result_array[1][44] ,
         \result_array[1][43] , \result_array[1][42] , \result_array[1][41] ,
         \result_array[1][40] , \result_array[1][39] , \result_array[1][38] ,
         \result_array[1][37] , \result_array[1][36] , \result_array[1][35] ,
         \result_array[1][34] , \result_array[1][33] , \result_array[1][32] ,
         \result_array[1][31] , \result_array[1][30] , \result_array[1][29] ,
         \result_array[1][28] , \result_array[1][27] , \result_array[1][26] ,
         \result_array[1][25] , \result_array[1][24] , \result_array[1][23] ,
         \result_array[1][22] , \result_array[1][21] , \result_array[1][20] ,
         \result_array[1][19] , \result_array[1][18] , \result_array[1][17] ,
         \result_array[1][16] , \result_array[1][15] , \result_array[1][14] ,
         \result_array[1][13] , \result_array[1][12] , \result_array[1][11] ,
         \result_array[1][10] , \result_array[1][9] , \result_array[1][8] ,
         \result_array[1][7] , \result_array[1][6] , \result_array[1][5] ,
         \result_array[1][4] , \result_array[1][3] , \result_array[1][2] ,
         \result_array[1][1] , \result_array[1][0] , \result_array[0][63] ,
         \result_array[0][62] , \result_array[0][61] , \result_array[0][60] ,
         \result_array[0][59] , \result_array[0][58] , \result_array[0][57] ,
         \result_array[0][56] , \result_array[0][55] , \result_array[0][54] ,
         \result_array[0][53] , \result_array[0][52] , \result_array[0][51] ,
         \result_array[0][50] , \result_array[0][49] , \result_array[0][48] ,
         \result_array[0][47] , \result_array[0][46] , \result_array[0][45] ,
         \result_array[0][44] , \result_array[0][43] , \result_array[0][42] ,
         \result_array[0][41] , \result_array[0][40] , \result_array[0][39] ,
         \result_array[0][38] , \result_array[0][37] , \result_array[0][36] ,
         \result_array[0][35] , \result_array[0][34] , \result_array[0][33] ,
         \result_array[0][32] , \result_array[0][31] , \result_array[0][30] ,
         \result_array[0][29] , \result_array[0][28] , \result_array[0][27] ,
         \result_array[0][26] , \result_array[0][25] , \result_array[0][24] ,
         \result_array[0][23] , \result_array[0][22] , \result_array[0][21] ,
         \result_array[0][20] , \result_array[0][19] , \result_array[0][18] ,
         \result_array[0][17] , \result_array[0][16] , \result_array[0][15] ,
         \result_array[0][14] , \result_array[0][13] , \result_array[0][12] ,
         \result_array[0][11] , \result_array[0][10] , \result_array[0][9] ,
         \result_array[0][8] , \result_array[0][7] , \result_array[0][6] ,
         \result_array[0][5] , \result_array[0][4] , \result_array[0][3] ,
         \result_array[0][2] , \result_array[0][1] , \result_array[0][0] ,
         \array_mux_out[7][63] , \array_mux_out[7][62] ,
         \array_mux_out[7][61] , \array_mux_out[7][60] ,
         \array_mux_out[7][59] , \array_mux_out[7][58] ,
         \array_mux_out[7][57] , \array_mux_out[7][56] ,
         \array_mux_out[7][55] , \array_mux_out[7][54] ,
         \array_mux_out[7][53] , \array_mux_out[7][52] ,
         \array_mux_out[7][51] , \array_mux_out[7][50] ,
         \array_mux_out[7][49] , \array_mux_out[7][48] ,
         \array_mux_out[7][47] , \array_mux_out[7][46] ,
         \array_mux_out[7][45] , \array_mux_out[7][44] ,
         \array_mux_out[7][43] , \array_mux_out[7][42] ,
         \array_mux_out[7][41] , \array_mux_out[7][40] ,
         \array_mux_out[7][39] , \array_mux_out[7][38] ,
         \array_mux_out[7][37] , \array_mux_out[7][36] ,
         \array_mux_out[7][35] , \array_mux_out[7][34] ,
         \array_mux_out[7][33] , \array_mux_out[7][32] ,
         \array_mux_out[7][31] , \array_mux_out[7][30] ,
         \array_mux_out[7][29] , \array_mux_out[7][28] ,
         \array_mux_out[7][27] , \array_mux_out[7][26] ,
         \array_mux_out[7][25] , \array_mux_out[7][24] ,
         \array_mux_out[7][23] , \array_mux_out[7][22] ,
         \array_mux_out[7][21] , \array_mux_out[7][20] ,
         \array_mux_out[7][19] , \array_mux_out[7][18] ,
         \array_mux_out[7][17] , \array_mux_out[7][16] ,
         \array_mux_out[7][15] , \array_mux_out[7][14] ,
         \array_mux_out[7][13] , \array_mux_out[7][12] ,
         \array_mux_out[7][11] , \array_mux_out[7][10] , \array_mux_out[7][9] ,
         \array_mux_out[7][8] , \array_mux_out[7][7] , \array_mux_out[7][6] ,
         \array_mux_out[7][5] , \array_mux_out[7][4] , \array_mux_out[7][3] ,
         \array_mux_out[7][2] , \array_mux_out[7][1] , \array_mux_out[7][0] ,
         \array_mux_out[6][63] , \array_mux_out[6][62] ,
         \array_mux_out[6][61] , \array_mux_out[6][60] ,
         \array_mux_out[6][59] , \array_mux_out[6][58] ,
         \array_mux_out[6][57] , \array_mux_out[6][56] ,
         \array_mux_out[6][55] , \array_mux_out[6][54] ,
         \array_mux_out[6][53] , \array_mux_out[6][52] ,
         \array_mux_out[6][51] , \array_mux_out[6][50] ,
         \array_mux_out[6][49] , \array_mux_out[6][48] ,
         \array_mux_out[6][47] , \array_mux_out[6][46] ,
         \array_mux_out[6][45] , \array_mux_out[6][44] ,
         \array_mux_out[6][43] , \array_mux_out[6][42] ,
         \array_mux_out[6][41] , \array_mux_out[6][40] ,
         \array_mux_out[6][39] , \array_mux_out[6][38] ,
         \array_mux_out[6][37] , \array_mux_out[6][36] ,
         \array_mux_out[6][35] , \array_mux_out[6][34] ,
         \array_mux_out[6][33] , \array_mux_out[6][32] ,
         \array_mux_out[6][31] , \array_mux_out[6][30] ,
         \array_mux_out[6][29] , \array_mux_out[6][28] ,
         \array_mux_out[6][27] , \array_mux_out[6][26] ,
         \array_mux_out[6][25] , \array_mux_out[6][24] ,
         \array_mux_out[6][23] , \array_mux_out[6][22] ,
         \array_mux_out[6][21] , \array_mux_out[6][20] ,
         \array_mux_out[6][19] , \array_mux_out[6][18] ,
         \array_mux_out[6][17] , \array_mux_out[6][16] ,
         \array_mux_out[6][15] , \array_mux_out[6][14] ,
         \array_mux_out[6][13] , \array_mux_out[6][12] ,
         \array_mux_out[6][11] , \array_mux_out[6][10] , \array_mux_out[6][9] ,
         \array_mux_out[6][8] , \array_mux_out[6][7] , \array_mux_out[6][6] ,
         \array_mux_out[6][5] , \array_mux_out[6][4] , \array_mux_out[6][3] ,
         \array_mux_out[6][2] , \array_mux_out[6][1] , \array_mux_out[6][0] ,
         \array_mux_out[5][63] , \array_mux_out[5][62] ,
         \array_mux_out[5][61] , \array_mux_out[5][60] ,
         \array_mux_out[5][59] , \array_mux_out[5][58] ,
         \array_mux_out[5][57] , \array_mux_out[5][56] ,
         \array_mux_out[5][55] , \array_mux_out[5][54] ,
         \array_mux_out[5][53] , \array_mux_out[5][52] ,
         \array_mux_out[5][51] , \array_mux_out[5][50] ,
         \array_mux_out[5][49] , \array_mux_out[5][48] ,
         \array_mux_out[5][47] , \array_mux_out[5][46] ,
         \array_mux_out[5][45] , \array_mux_out[5][44] ,
         \array_mux_out[5][43] , \array_mux_out[5][42] ,
         \array_mux_out[5][41] , \array_mux_out[5][40] ,
         \array_mux_out[5][39] , \array_mux_out[5][38] ,
         \array_mux_out[5][37] , \array_mux_out[5][36] ,
         \array_mux_out[5][35] , \array_mux_out[5][34] ,
         \array_mux_out[5][33] , \array_mux_out[5][32] ,
         \array_mux_out[5][31] , \array_mux_out[5][30] ,
         \array_mux_out[5][29] , \array_mux_out[5][28] ,
         \array_mux_out[5][27] , \array_mux_out[5][26] ,
         \array_mux_out[5][25] , \array_mux_out[5][24] ,
         \array_mux_out[5][23] , \array_mux_out[5][22] ,
         \array_mux_out[5][21] , \array_mux_out[5][20] ,
         \array_mux_out[5][19] , \array_mux_out[5][18] ,
         \array_mux_out[5][17] , \array_mux_out[5][16] ,
         \array_mux_out[5][15] , \array_mux_out[5][14] ,
         \array_mux_out[5][13] , \array_mux_out[5][12] ,
         \array_mux_out[5][11] , \array_mux_out[5][10] , \array_mux_out[5][9] ,
         \array_mux_out[5][8] , \array_mux_out[5][7] , \array_mux_out[5][6] ,
         \array_mux_out[5][5] , \array_mux_out[5][4] , \array_mux_out[5][3] ,
         \array_mux_out[5][2] , \array_mux_out[5][1] , \array_mux_out[5][0] ,
         \array_mux_out[4][63] , \array_mux_out[4][62] ,
         \array_mux_out[4][61] , \array_mux_out[4][60] ,
         \array_mux_out[4][59] , \array_mux_out[4][58] ,
         \array_mux_out[4][57] , \array_mux_out[4][56] ,
         \array_mux_out[4][55] , \array_mux_out[4][54] ,
         \array_mux_out[4][53] , \array_mux_out[4][52] ,
         \array_mux_out[4][51] , \array_mux_out[4][50] ,
         \array_mux_out[4][49] , \array_mux_out[4][48] ,
         \array_mux_out[4][47] , \array_mux_out[4][46] ,
         \array_mux_out[4][45] , \array_mux_out[4][44] ,
         \array_mux_out[4][43] , \array_mux_out[4][42] ,
         \array_mux_out[4][41] , \array_mux_out[4][40] ,
         \array_mux_out[4][39] , \array_mux_out[4][38] ,
         \array_mux_out[4][37] , \array_mux_out[4][36] ,
         \array_mux_out[4][35] , \array_mux_out[4][34] ,
         \array_mux_out[4][33] , \array_mux_out[4][32] ,
         \array_mux_out[4][31] , \array_mux_out[4][30] ,
         \array_mux_out[4][29] , \array_mux_out[4][28] ,
         \array_mux_out[4][27] , \array_mux_out[4][26] ,
         \array_mux_out[4][25] , \array_mux_out[4][24] ,
         \array_mux_out[4][23] , \array_mux_out[4][22] ,
         \array_mux_out[4][21] , \array_mux_out[4][20] ,
         \array_mux_out[4][19] , \array_mux_out[4][18] ,
         \array_mux_out[4][17] , \array_mux_out[4][16] ,
         \array_mux_out[4][15] , \array_mux_out[4][14] ,
         \array_mux_out[4][13] , \array_mux_out[4][12] ,
         \array_mux_out[4][11] , \array_mux_out[4][10] , \array_mux_out[4][9] ,
         \array_mux_out[4][8] , \array_mux_out[4][7] , \array_mux_out[4][6] ,
         \array_mux_out[4][5] , \array_mux_out[4][4] , \array_mux_out[4][3] ,
         \array_mux_out[4][2] , \array_mux_out[4][1] , \array_mux_out[4][0] ,
         \array_mux_out[3][63] , \array_mux_out[3][62] ,
         \array_mux_out[3][61] , \array_mux_out[3][60] ,
         \array_mux_out[3][59] , \array_mux_out[3][58] ,
         \array_mux_out[3][57] , \array_mux_out[3][56] ,
         \array_mux_out[3][55] , \array_mux_out[3][54] ,
         \array_mux_out[3][53] , \array_mux_out[3][52] ,
         \array_mux_out[3][51] , \array_mux_out[3][50] ,
         \array_mux_out[3][49] , \array_mux_out[3][48] ,
         \array_mux_out[3][47] , \array_mux_out[3][46] ,
         \array_mux_out[3][45] , \array_mux_out[3][44] ,
         \array_mux_out[3][43] , \array_mux_out[3][42] ,
         \array_mux_out[3][41] , \array_mux_out[3][40] ,
         \array_mux_out[3][39] , \array_mux_out[3][38] ,
         \array_mux_out[3][37] , \array_mux_out[3][36] ,
         \array_mux_out[3][35] , \array_mux_out[3][34] ,
         \array_mux_out[3][33] , \array_mux_out[3][32] ,
         \array_mux_out[3][31] , \array_mux_out[3][30] ,
         \array_mux_out[3][29] , \array_mux_out[3][28] ,
         \array_mux_out[3][27] , \array_mux_out[3][26] ,
         \array_mux_out[3][25] , \array_mux_out[3][24] ,
         \array_mux_out[3][23] , \array_mux_out[3][22] ,
         \array_mux_out[3][21] , \array_mux_out[3][20] ,
         \array_mux_out[3][19] , \array_mux_out[3][18] ,
         \array_mux_out[3][17] , \array_mux_out[3][16] ,
         \array_mux_out[3][15] , \array_mux_out[3][14] ,
         \array_mux_out[3][13] , \array_mux_out[3][12] ,
         \array_mux_out[3][11] , \array_mux_out[3][10] , \array_mux_out[3][9] ,
         \array_mux_out[3][8] , \array_mux_out[3][7] , \array_mux_out[3][6] ,
         \array_mux_out[3][5] , \array_mux_out[3][4] , \array_mux_out[3][3] ,
         \array_mux_out[3][2] , \array_mux_out[3][1] , \array_mux_out[3][0] ,
         \array_mux_out[2][63] , \array_mux_out[2][62] ,
         \array_mux_out[2][61] , \array_mux_out[2][60] ,
         \array_mux_out[2][59] , \array_mux_out[2][58] ,
         \array_mux_out[2][57] , \array_mux_out[2][56] ,
         \array_mux_out[2][55] , \array_mux_out[2][54] ,
         \array_mux_out[2][53] , \array_mux_out[2][52] ,
         \array_mux_out[2][51] , \array_mux_out[2][50] ,
         \array_mux_out[2][49] , \array_mux_out[2][48] ,
         \array_mux_out[2][47] , \array_mux_out[2][46] ,
         \array_mux_out[2][45] , \array_mux_out[2][44] ,
         \array_mux_out[2][43] , \array_mux_out[2][42] ,
         \array_mux_out[2][41] , \array_mux_out[2][40] ,
         \array_mux_out[2][39] , \array_mux_out[2][38] ,
         \array_mux_out[2][37] , \array_mux_out[2][36] ,
         \array_mux_out[2][35] , \array_mux_out[2][34] ,
         \array_mux_out[2][33] , \array_mux_out[2][32] ,
         \array_mux_out[2][31] , \array_mux_out[2][30] ,
         \array_mux_out[2][29] , \array_mux_out[2][28] ,
         \array_mux_out[2][27] , \array_mux_out[2][26] ,
         \array_mux_out[2][25] , \array_mux_out[2][24] ,
         \array_mux_out[2][23] , \array_mux_out[2][22] ,
         \array_mux_out[2][21] , \array_mux_out[2][20] ,
         \array_mux_out[2][19] , \array_mux_out[2][18] ,
         \array_mux_out[2][17] , \array_mux_out[2][16] ,
         \array_mux_out[2][15] , \array_mux_out[2][14] ,
         \array_mux_out[2][13] , \array_mux_out[2][12] ,
         \array_mux_out[2][11] , \array_mux_out[2][10] , \array_mux_out[2][9] ,
         \array_mux_out[2][8] , \array_mux_out[2][7] , \array_mux_out[2][6] ,
         \array_mux_out[2][5] , \array_mux_out[2][4] , \array_mux_out[2][3] ,
         \array_mux_out[2][2] , \array_mux_out[2][1] , \array_mux_out[2][0] ,
         \array_mux_out[1][63] , \array_mux_out[1][62] ,
         \array_mux_out[1][61] , \array_mux_out[1][60] ,
         \array_mux_out[1][59] , \array_mux_out[1][58] ,
         \array_mux_out[1][57] , \array_mux_out[1][56] ,
         \array_mux_out[1][55] , \array_mux_out[1][54] ,
         \array_mux_out[1][53] , \array_mux_out[1][52] ,
         \array_mux_out[1][51] , \array_mux_out[1][50] ,
         \array_mux_out[1][49] , \array_mux_out[1][48] ,
         \array_mux_out[1][47] , \array_mux_out[1][46] ,
         \array_mux_out[1][45] , \array_mux_out[1][44] ,
         \array_mux_out[1][43] , \array_mux_out[1][42] ,
         \array_mux_out[1][41] , \array_mux_out[1][40] ,
         \array_mux_out[1][39] , \array_mux_out[1][38] ,
         \array_mux_out[1][37] , \array_mux_out[1][36] ,
         \array_mux_out[1][35] , \array_mux_out[1][34] ,
         \array_mux_out[1][33] , \array_mux_out[1][32] ,
         \array_mux_out[1][31] , \array_mux_out[1][30] ,
         \array_mux_out[1][29] , \array_mux_out[1][28] ,
         \array_mux_out[1][27] , \array_mux_out[1][26] ,
         \array_mux_out[1][25] , \array_mux_out[1][24] ,
         \array_mux_out[1][23] , \array_mux_out[1][22] ,
         \array_mux_out[1][21] , \array_mux_out[1][20] ,
         \array_mux_out[1][19] , \array_mux_out[1][18] ,
         \array_mux_out[1][17] , \array_mux_out[1][16] ,
         \array_mux_out[1][15] , \array_mux_out[1][14] ,
         \array_mux_out[1][13] , \array_mux_out[1][12] ,
         \array_mux_out[1][11] , \array_mux_out[1][10] , \array_mux_out[1][9] ,
         \array_mux_out[1][8] , \array_mux_out[1][7] , \array_mux_out[1][6] ,
         \array_mux_out[1][5] , \array_mux_out[1][4] , \array_mux_out[1][3] ,
         \array_mux_out[1][2] , \array_mux_out[1][1] , \array_mux_out[1][0] ,
         \array_mux_out[15][63] , \array_mux_out[15][62] ,
         \array_mux_out[15][61] , \array_mux_out[15][60] ,
         \array_mux_out[15][59] , \array_mux_out[15][58] ,
         \array_mux_out[15][57] , \array_mux_out[15][56] ,
         \array_mux_out[15][55] , \array_mux_out[15][54] ,
         \array_mux_out[15][53] , \array_mux_out[15][52] ,
         \array_mux_out[15][51] , \array_mux_out[15][50] ,
         \array_mux_out[15][49] , \array_mux_out[15][48] ,
         \array_mux_out[15][47] , \array_mux_out[15][46] ,
         \array_mux_out[15][45] , \array_mux_out[15][44] ,
         \array_mux_out[15][43] , \array_mux_out[15][42] ,
         \array_mux_out[15][41] , \array_mux_out[15][40] ,
         \array_mux_out[15][39] , \array_mux_out[15][38] ,
         \array_mux_out[15][37] , \array_mux_out[15][36] ,
         \array_mux_out[15][35] , \array_mux_out[15][34] ,
         \array_mux_out[15][33] , \array_mux_out[15][32] ,
         \array_mux_out[15][31] , \array_mux_out[15][30] ,
         \array_mux_out[15][29] , \array_mux_out[15][28] ,
         \array_mux_out[15][27] , \array_mux_out[15][26] ,
         \array_mux_out[15][25] , \array_mux_out[15][24] ,
         \array_mux_out[15][23] , \array_mux_out[15][22] ,
         \array_mux_out[15][21] , \array_mux_out[15][20] ,
         \array_mux_out[15][19] , \array_mux_out[15][18] ,
         \array_mux_out[15][17] , \array_mux_out[15][16] ,
         \array_mux_out[15][15] , \array_mux_out[15][14] ,
         \array_mux_out[15][13] , \array_mux_out[15][12] ,
         \array_mux_out[15][11] , \array_mux_out[15][10] ,
         \array_mux_out[15][9] , \array_mux_out[15][8] ,
         \array_mux_out[15][7] , \array_mux_out[15][6] ,
         \array_mux_out[15][5] , \array_mux_out[15][4] ,
         \array_mux_out[15][3] , \array_mux_out[15][2] ,
         \array_mux_out[15][1] , \array_mux_out[15][0] ,
         \array_mux_out[14][63] , \array_mux_out[14][62] ,
         \array_mux_out[14][61] , \array_mux_out[14][60] ,
         \array_mux_out[14][59] , \array_mux_out[14][58] ,
         \array_mux_out[14][57] , \array_mux_out[14][56] ,
         \array_mux_out[14][55] , \array_mux_out[14][54] ,
         \array_mux_out[14][53] , \array_mux_out[14][52] ,
         \array_mux_out[14][51] , \array_mux_out[14][50] ,
         \array_mux_out[14][49] , \array_mux_out[14][48] ,
         \array_mux_out[14][47] , \array_mux_out[14][46] ,
         \array_mux_out[14][45] , \array_mux_out[14][44] ,
         \array_mux_out[14][43] , \array_mux_out[14][42] ,
         \array_mux_out[14][41] , \array_mux_out[14][40] ,
         \array_mux_out[14][39] , \array_mux_out[14][38] ,
         \array_mux_out[14][37] , \array_mux_out[14][36] ,
         \array_mux_out[14][35] , \array_mux_out[14][34] ,
         \array_mux_out[14][33] , \array_mux_out[14][32] ,
         \array_mux_out[14][31] , \array_mux_out[14][30] ,
         \array_mux_out[14][29] , \array_mux_out[14][28] ,
         \array_mux_out[14][27] , \array_mux_out[14][26] ,
         \array_mux_out[14][25] , \array_mux_out[14][24] ,
         \array_mux_out[14][23] , \array_mux_out[14][22] ,
         \array_mux_out[14][21] , \array_mux_out[14][20] ,
         \array_mux_out[14][19] , \array_mux_out[14][18] ,
         \array_mux_out[14][17] , \array_mux_out[14][16] ,
         \array_mux_out[14][15] , \array_mux_out[14][14] ,
         \array_mux_out[14][13] , \array_mux_out[14][12] ,
         \array_mux_out[14][11] , \array_mux_out[14][10] ,
         \array_mux_out[14][9] , \array_mux_out[14][8] ,
         \array_mux_out[14][7] , \array_mux_out[14][6] ,
         \array_mux_out[14][5] , \array_mux_out[14][4] ,
         \array_mux_out[14][3] , \array_mux_out[14][2] ,
         \array_mux_out[14][1] , \array_mux_out[14][0] ,
         \array_mux_out[13][63] , \array_mux_out[13][62] ,
         \array_mux_out[13][61] , \array_mux_out[13][60] ,
         \array_mux_out[13][59] , \array_mux_out[13][58] ,
         \array_mux_out[13][57] , \array_mux_out[13][56] ,
         \array_mux_out[13][55] , \array_mux_out[13][54] ,
         \array_mux_out[13][53] , \array_mux_out[13][52] ,
         \array_mux_out[13][51] , \array_mux_out[13][50] ,
         \array_mux_out[13][49] , \array_mux_out[13][48] ,
         \array_mux_out[13][47] , \array_mux_out[13][46] ,
         \array_mux_out[13][45] , \array_mux_out[13][44] ,
         \array_mux_out[13][43] , \array_mux_out[13][42] ,
         \array_mux_out[13][41] , \array_mux_out[13][40] ,
         \array_mux_out[13][39] , \array_mux_out[13][38] ,
         \array_mux_out[13][37] , \array_mux_out[13][36] ,
         \array_mux_out[13][35] , \array_mux_out[13][34] ,
         \array_mux_out[13][33] , \array_mux_out[13][32] ,
         \array_mux_out[13][31] , \array_mux_out[13][30] ,
         \array_mux_out[13][29] , \array_mux_out[13][28] ,
         \array_mux_out[13][27] , \array_mux_out[13][26] ,
         \array_mux_out[13][25] , \array_mux_out[13][24] ,
         \array_mux_out[13][23] , \array_mux_out[13][22] ,
         \array_mux_out[13][21] , \array_mux_out[13][20] ,
         \array_mux_out[13][19] , \array_mux_out[13][18] ,
         \array_mux_out[13][17] , \array_mux_out[13][16] ,
         \array_mux_out[13][15] , \array_mux_out[13][14] ,
         \array_mux_out[13][13] , \array_mux_out[13][12] ,
         \array_mux_out[13][11] , \array_mux_out[13][10] ,
         \array_mux_out[13][9] , \array_mux_out[13][8] ,
         \array_mux_out[13][7] , \array_mux_out[13][6] ,
         \array_mux_out[13][5] , \array_mux_out[13][4] ,
         \array_mux_out[13][3] , \array_mux_out[13][2] ,
         \array_mux_out[13][1] , \array_mux_out[13][0] ,
         \array_mux_out[12][63] , \array_mux_out[12][62] ,
         \array_mux_out[12][61] , \array_mux_out[12][60] ,
         \array_mux_out[12][59] , \array_mux_out[12][58] ,
         \array_mux_out[12][57] , \array_mux_out[12][56] ,
         \array_mux_out[12][55] , \array_mux_out[12][54] ,
         \array_mux_out[12][53] , \array_mux_out[12][52] ,
         \array_mux_out[12][51] , \array_mux_out[12][50] ,
         \array_mux_out[12][49] , \array_mux_out[12][48] ,
         \array_mux_out[12][47] , \array_mux_out[12][46] ,
         \array_mux_out[12][45] , \array_mux_out[12][44] ,
         \array_mux_out[12][43] , \array_mux_out[12][42] ,
         \array_mux_out[12][41] , \array_mux_out[12][40] ,
         \array_mux_out[12][39] , \array_mux_out[12][38] ,
         \array_mux_out[12][37] , \array_mux_out[12][36] ,
         \array_mux_out[12][35] , \array_mux_out[12][34] ,
         \array_mux_out[12][33] , \array_mux_out[12][32] ,
         \array_mux_out[12][31] , \array_mux_out[12][30] ,
         \array_mux_out[12][29] , \array_mux_out[12][28] ,
         \array_mux_out[12][27] , \array_mux_out[12][26] ,
         \array_mux_out[12][25] , \array_mux_out[12][24] ,
         \array_mux_out[12][23] , \array_mux_out[12][22] ,
         \array_mux_out[12][21] , \array_mux_out[12][20] ,
         \array_mux_out[12][19] , \array_mux_out[12][18] ,
         \array_mux_out[12][17] , \array_mux_out[12][16] ,
         \array_mux_out[12][15] , \array_mux_out[12][14] ,
         \array_mux_out[12][13] , \array_mux_out[12][12] ,
         \array_mux_out[12][11] , \array_mux_out[12][10] ,
         \array_mux_out[12][9] , \array_mux_out[12][8] ,
         \array_mux_out[12][7] , \array_mux_out[12][6] ,
         \array_mux_out[12][5] , \array_mux_out[12][4] ,
         \array_mux_out[12][3] , \array_mux_out[12][2] ,
         \array_mux_out[12][1] , \array_mux_out[12][0] ,
         \array_mux_out[11][63] , \array_mux_out[11][62] ,
         \array_mux_out[11][61] , \array_mux_out[11][60] ,
         \array_mux_out[11][59] , \array_mux_out[11][58] ,
         \array_mux_out[11][57] , \array_mux_out[11][56] ,
         \array_mux_out[11][55] , \array_mux_out[11][54] ,
         \array_mux_out[11][53] , \array_mux_out[11][52] ,
         \array_mux_out[11][51] , \array_mux_out[11][50] ,
         \array_mux_out[11][49] , \array_mux_out[11][48] ,
         \array_mux_out[11][47] , \array_mux_out[11][46] ,
         \array_mux_out[11][45] , \array_mux_out[11][44] ,
         \array_mux_out[11][43] , \array_mux_out[11][42] ,
         \array_mux_out[11][41] , \array_mux_out[11][40] ,
         \array_mux_out[11][39] , \array_mux_out[11][38] ,
         \array_mux_out[11][37] , \array_mux_out[11][36] ,
         \array_mux_out[11][35] , \array_mux_out[11][34] ,
         \array_mux_out[11][33] , \array_mux_out[11][32] ,
         \array_mux_out[11][31] , \array_mux_out[11][30] ,
         \array_mux_out[11][29] , \array_mux_out[11][28] ,
         \array_mux_out[11][27] , \array_mux_out[11][26] ,
         \array_mux_out[11][25] , \array_mux_out[11][24] ,
         \array_mux_out[11][23] , \array_mux_out[11][22] ,
         \array_mux_out[11][21] , \array_mux_out[11][20] ,
         \array_mux_out[11][19] , \array_mux_out[11][18] ,
         \array_mux_out[11][17] , \array_mux_out[11][16] ,
         \array_mux_out[11][15] , \array_mux_out[11][14] ,
         \array_mux_out[11][13] , \array_mux_out[11][12] ,
         \array_mux_out[11][11] , \array_mux_out[11][10] ,
         \array_mux_out[11][9] , \array_mux_out[11][8] ,
         \array_mux_out[11][7] , \array_mux_out[11][6] ,
         \array_mux_out[11][5] , \array_mux_out[11][4] ,
         \array_mux_out[11][3] , \array_mux_out[11][2] ,
         \array_mux_out[11][1] , \array_mux_out[11][0] ,
         \array_mux_out[10][63] , \array_mux_out[10][62] ,
         \array_mux_out[10][61] , \array_mux_out[10][60] ,
         \array_mux_out[10][59] , \array_mux_out[10][58] ,
         \array_mux_out[10][57] , \array_mux_out[10][56] ,
         \array_mux_out[10][55] , \array_mux_out[10][54] ,
         \array_mux_out[10][53] , \array_mux_out[10][52] ,
         \array_mux_out[10][51] , \array_mux_out[10][50] ,
         \array_mux_out[10][49] , \array_mux_out[10][48] ,
         \array_mux_out[10][47] , \array_mux_out[10][46] ,
         \array_mux_out[10][45] , \array_mux_out[10][44] ,
         \array_mux_out[10][43] , \array_mux_out[10][42] ,
         \array_mux_out[10][41] , \array_mux_out[10][40] ,
         \array_mux_out[10][39] , \array_mux_out[10][38] ,
         \array_mux_out[10][37] , \array_mux_out[10][36] ,
         \array_mux_out[10][35] , \array_mux_out[10][34] ,
         \array_mux_out[10][33] , \array_mux_out[10][32] ,
         \array_mux_out[10][31] , \array_mux_out[10][30] ,
         \array_mux_out[10][29] , \array_mux_out[10][28] ,
         \array_mux_out[10][27] , \array_mux_out[10][26] ,
         \array_mux_out[10][25] , \array_mux_out[10][24] ,
         \array_mux_out[10][23] , \array_mux_out[10][22] ,
         \array_mux_out[10][21] , \array_mux_out[10][20] ,
         \array_mux_out[10][19] , \array_mux_out[10][18] ,
         \array_mux_out[10][17] , \array_mux_out[10][16] ,
         \array_mux_out[10][15] , \array_mux_out[10][14] ,
         \array_mux_out[10][13] , \array_mux_out[10][12] ,
         \array_mux_out[10][11] , \array_mux_out[10][10] ,
         \array_mux_out[10][9] , \array_mux_out[10][8] ,
         \array_mux_out[10][7] , \array_mux_out[10][6] ,
         \array_mux_out[10][5] , \array_mux_out[10][4] ,
         \array_mux_out[10][3] , \array_mux_out[10][2] ,
         \array_mux_out[10][1] , \array_mux_out[10][0] ,
         \array_mux_out[9][63] , \array_mux_out[9][62] ,
         \array_mux_out[9][61] , \array_mux_out[9][60] ,
         \array_mux_out[9][59] , \array_mux_out[9][58] ,
         \array_mux_out[9][57] , \array_mux_out[9][56] ,
         \array_mux_out[9][55] , \array_mux_out[9][54] ,
         \array_mux_out[9][53] , \array_mux_out[9][52] ,
         \array_mux_out[9][51] , \array_mux_out[9][50] ,
         \array_mux_out[9][49] , \array_mux_out[9][48] ,
         \array_mux_out[9][47] , \array_mux_out[9][46] ,
         \array_mux_out[9][45] , \array_mux_out[9][44] ,
         \array_mux_out[9][43] , \array_mux_out[9][42] ,
         \array_mux_out[9][41] , \array_mux_out[9][40] ,
         \array_mux_out[9][39] , \array_mux_out[9][38] ,
         \array_mux_out[9][37] , \array_mux_out[9][36] ,
         \array_mux_out[9][35] , \array_mux_out[9][34] ,
         \array_mux_out[9][33] , \array_mux_out[9][32] ,
         \array_mux_out[9][31] , \array_mux_out[9][30] ,
         \array_mux_out[9][29] , \array_mux_out[9][28] ,
         \array_mux_out[9][27] , \array_mux_out[9][26] ,
         \array_mux_out[9][25] , \array_mux_out[9][24] ,
         \array_mux_out[9][23] , \array_mux_out[9][22] ,
         \array_mux_out[9][21] , \array_mux_out[9][20] ,
         \array_mux_out[9][19] , \array_mux_out[9][18] ,
         \array_mux_out[9][17] , \array_mux_out[9][16] ,
         \array_mux_out[9][15] , \array_mux_out[9][14] ,
         \array_mux_out[9][13] , \array_mux_out[9][12] ,
         \array_mux_out[9][11] , \array_mux_out[9][10] , \array_mux_out[9][9] ,
         \array_mux_out[9][8] , \array_mux_out[9][7] , \array_mux_out[9][6] ,
         \array_mux_out[9][5] , \array_mux_out[9][4] , \array_mux_out[9][3] ,
         \array_mux_out[9][2] , \array_mux_out[9][1] , \array_mux_out[9][0] ,
         \array_mux_out[8][63] , \array_mux_out[8][62] ,
         \array_mux_out[8][61] , \array_mux_out[8][60] ,
         \array_mux_out[8][59] , \array_mux_out[8][58] ,
         \array_mux_out[8][57] , \array_mux_out[8][56] ,
         \array_mux_out[8][55] , \array_mux_out[8][54] ,
         \array_mux_out[8][53] , \array_mux_out[8][52] ,
         \array_mux_out[8][51] , \array_mux_out[8][50] ,
         \array_mux_out[8][49] , \array_mux_out[8][48] ,
         \array_mux_out[8][47] , \array_mux_out[8][46] ,
         \array_mux_out[8][45] , \array_mux_out[8][44] ,
         \array_mux_out[8][43] , \array_mux_out[8][42] ,
         \array_mux_out[8][41] , \array_mux_out[8][40] ,
         \array_mux_out[8][39] , \array_mux_out[8][38] ,
         \array_mux_out[8][37] , \array_mux_out[8][36] ,
         \array_mux_out[8][35] , \array_mux_out[8][34] ,
         \array_mux_out[8][33] , \array_mux_out[8][32] ,
         \array_mux_out[8][31] , \array_mux_out[8][30] ,
         \array_mux_out[8][29] , \array_mux_out[8][28] ,
         \array_mux_out[8][27] , \array_mux_out[8][26] ,
         \array_mux_out[8][25] , \array_mux_out[8][24] ,
         \array_mux_out[8][23] , \array_mux_out[8][22] ,
         \array_mux_out[8][21] , \array_mux_out[8][20] ,
         \array_mux_out[8][19] , \array_mux_out[8][18] ,
         \array_mux_out[8][17] , \array_mux_out[8][16] ,
         \array_mux_out[8][15] , \array_mux_out[8][14] ,
         \array_mux_out[8][13] , \array_mux_out[8][12] ,
         \array_mux_out[8][11] , \array_mux_out[8][10] , \array_mux_out[8][9] ,
         \array_mux_out[8][8] , \array_mux_out[8][7] , \array_mux_out[8][6] ,
         \array_mux_out[8][5] , \array_mux_out[8][4] , \array_mux_out[8][3] ,
         \array_mux_out[8][2] , \array_mux_out[8][1] , \array_mux_out[8][0] ,
         \result_array[14][63] , \result_array[14][62] ,
         \result_array[14][61] , \result_array[14][60] ,
         \result_array[14][59] , \result_array[14][58] ,
         \result_array[14][57] , \result_array[14][56] ,
         \result_array[14][55] , \result_array[14][54] ,
         \result_array[14][53] , \result_array[14][52] ,
         \result_array[14][51] , \result_array[14][50] ,
         \result_array[14][49] , \result_array[14][48] ,
         \result_array[14][47] , \result_array[14][46] ,
         \result_array[14][45] , \result_array[14][44] ,
         \result_array[14][43] , \result_array[14][42] ,
         \result_array[14][41] , \result_array[14][40] ,
         \result_array[14][39] , \result_array[14][38] ,
         \result_array[14][37] , \result_array[14][36] ,
         \result_array[14][35] , \result_array[14][34] ,
         \result_array[14][33] , \result_array[14][32] ,
         \result_array[14][31] , \result_array[14][30] ,
         \result_array[14][29] , \result_array[14][28] ,
         \result_array[14][27] , \result_array[14][26] ,
         \result_array[14][25] , \result_array[14][24] ,
         \result_array[14][23] , \result_array[14][22] ,
         \result_array[14][21] , \result_array[14][20] ,
         \result_array[14][19] , \result_array[14][18] ,
         \result_array[14][17] , \result_array[14][16] ,
         \result_array[14][15] , \result_array[14][14] ,
         \result_array[14][13] , \result_array[14][12] ,
         \result_array[14][11] , \result_array[14][10] , \result_array[14][9] ,
         \result_array[14][8] , \result_array[14][7] , \result_array[14][6] ,
         \result_array[14][5] , \result_array[14][4] , \result_array[14][3] ,
         \result_array[14][2] , \result_array[14][1] , \result_array[14][0] ,
         \result_array[13][63] , \result_array[13][62] ,
         \result_array[13][61] , \result_array[13][60] ,
         \result_array[13][59] , \result_array[13][58] ,
         \result_array[13][57] , \result_array[13][56] ,
         \result_array[13][55] , \result_array[13][54] ,
         \result_array[13][53] , \result_array[13][52] ,
         \result_array[13][51] , \result_array[13][50] ,
         \result_array[13][49] , \result_array[13][48] ,
         \result_array[13][47] , \result_array[13][46] ,
         \result_array[13][45] , \result_array[13][44] ,
         \result_array[13][43] , \result_array[13][42] ,
         \result_array[13][41] , \result_array[13][40] ,
         \result_array[13][39] , \result_array[13][38] ,
         \result_array[13][37] , \result_array[13][36] ,
         \result_array[13][35] , \result_array[13][34] ,
         \result_array[13][33] , \result_array[13][32] ,
         \result_array[13][31] , \result_array[13][30] ,
         \result_array[13][29] , \result_array[13][28] ,
         \result_array[13][27] , \result_array[13][26] ,
         \result_array[13][25] , \result_array[13][24] ,
         \result_array[13][23] , \result_array[13][22] ,
         \result_array[13][21] , \result_array[13][20] ,
         \result_array[13][19] , \result_array[13][18] ,
         \result_array[13][17] , \result_array[13][16] ,
         \result_array[13][15] , \result_array[13][14] ,
         \result_array[13][13] , \result_array[13][12] ,
         \result_array[13][11] , \result_array[13][10] , \result_array[13][9] ,
         \result_array[13][8] , \result_array[13][7] , \result_array[13][6] ,
         \result_array[13][5] , \result_array[13][4] , \result_array[13][3] ,
         \result_array[13][2] , \result_array[13][1] , \result_array[13][0] ,
         \result_array[12][63] , \result_array[12][62] ,
         \result_array[12][61] , \result_array[12][60] ,
         \result_array[12][59] , \result_array[12][58] ,
         \result_array[12][57] , \result_array[12][56] ,
         \result_array[12][55] , \result_array[12][54] ,
         \result_array[12][53] , \result_array[12][52] ,
         \result_array[12][51] , \result_array[12][50] ,
         \result_array[12][49] , \result_array[12][48] ,
         \result_array[12][47] , \result_array[12][46] ,
         \result_array[12][45] , \result_array[12][44] ,
         \result_array[12][43] , \result_array[12][42] ,
         \result_array[12][41] , \result_array[12][40] ,
         \result_array[12][39] , \result_array[12][38] ,
         \result_array[12][37] , \result_array[12][36] ,
         \result_array[12][35] , \result_array[12][34] ,
         \result_array[12][33] , \result_array[12][32] ,
         \result_array[12][31] , \result_array[12][30] ,
         \result_array[12][29] , \result_array[12][28] ,
         \result_array[12][27] , \result_array[12][26] ,
         \result_array[12][25] , \result_array[12][24] ,
         \result_array[12][23] , \result_array[12][22] ,
         \result_array[12][21] , \result_array[12][20] ,
         \result_array[12][19] , \result_array[12][18] ,
         \result_array[12][17] , \result_array[12][16] ,
         \result_array[12][15] , \result_array[12][14] ,
         \result_array[12][13] , \result_array[12][12] ,
         \result_array[12][11] , \result_array[12][10] , \result_array[12][9] ,
         \result_array[12][8] , \result_array[12][7] , \result_array[12][6] ,
         \result_array[12][5] , \result_array[12][4] , \result_array[12][3] ,
         \result_array[12][2] , \result_array[12][1] , \result_array[12][0] ,
         \result_array[11][63] , \result_array[11][62] ,
         \result_array[11][61] , \result_array[11][60] ,
         \result_array[11][59] , \result_array[11][58] ,
         \result_array[11][57] , \result_array[11][56] ,
         \result_array[11][55] , \result_array[11][54] ,
         \result_array[11][53] , \result_array[11][52] ,
         \result_array[11][51] , \result_array[11][50] ,
         \result_array[11][49] , \result_array[11][48] ,
         \result_array[11][47] , \result_array[11][46] ,
         \result_array[11][45] , \result_array[11][44] ,
         \result_array[11][43] , \result_array[11][42] ,
         \result_array[11][41] , \result_array[11][40] ,
         \result_array[11][39] , \result_array[11][38] ,
         \result_array[11][37] , \result_array[11][36] ,
         \result_array[11][35] , \result_array[11][34] ,
         \result_array[11][33] , \result_array[11][32] ,
         \result_array[11][31] , \result_array[11][30] ,
         \result_array[11][29] , \result_array[11][28] ,
         \result_array[11][27] , \result_array[11][26] ,
         \result_array[11][25] , \result_array[11][24] ,
         \result_array[11][23] , \result_array[11][22] ,
         \result_array[11][21] , \result_array[11][20] ,
         \result_array[11][19] , \result_array[11][18] ,
         \result_array[11][17] , \result_array[11][16] ,
         \result_array[11][15] , \result_array[11][14] ,
         \result_array[11][13] , \result_array[11][12] ,
         \result_array[11][11] , \result_array[11][10] , \result_array[11][9] ,
         \result_array[11][8] , \result_array[11][7] , \result_array[11][6] ,
         \result_array[11][5] , \result_array[11][4] , \result_array[11][3] ,
         \result_array[11][2] , \result_array[11][1] , \result_array[11][0] ,
         \result_array[10][63] , \result_array[10][62] ,
         \result_array[10][61] , \result_array[10][60] ,
         \result_array[10][59] , \result_array[10][58] ,
         \result_array[10][57] , \result_array[10][56] ,
         \result_array[10][55] , \result_array[10][54] ,
         \result_array[10][53] , \result_array[10][52] ,
         \result_array[10][51] , \result_array[10][50] ,
         \result_array[10][49] , \result_array[10][48] ,
         \result_array[10][47] , \result_array[10][46] ,
         \result_array[10][45] , \result_array[10][44] ,
         \result_array[10][43] , \result_array[10][42] ,
         \result_array[10][41] , \result_array[10][40] ,
         \result_array[10][39] , \result_array[10][38] ,
         \result_array[10][37] , \result_array[10][36] ,
         \result_array[10][35] , \result_array[10][34] ,
         \result_array[10][33] , \result_array[10][32] ,
         \result_array[10][31] , \result_array[10][30] ,
         \result_array[10][29] , \result_array[10][28] ,
         \result_array[10][27] , \result_array[10][26] ,
         \result_array[10][25] , \result_array[10][24] ,
         \result_array[10][23] , \result_array[10][22] ,
         \result_array[10][21] , \result_array[10][20] ,
         \result_array[10][19] , \result_array[10][18] ,
         \result_array[10][17] , \result_array[10][16] ,
         \result_array[10][15] , \result_array[10][14] ,
         \result_array[10][13] , \result_array[10][12] ,
         \result_array[10][11] , \result_array[10][10] , \result_array[10][9] ,
         \result_array[10][8] , \result_array[10][7] , \result_array[10][6] ,
         \result_array[10][5] , \result_array[10][4] , \result_array[10][3] ,
         \result_array[10][2] , \result_array[10][1] , \result_array[10][0] ,
         \result_array[9][63] , \result_array[9][62] , \result_array[9][61] ,
         \result_array[9][60] , \result_array[9][59] , \result_array[9][58] ,
         \result_array[9][57] , \result_array[9][56] , \result_array[9][55] ,
         \result_array[9][54] , \result_array[9][53] , \result_array[9][52] ,
         \result_array[9][51] , \result_array[9][50] , \result_array[9][49] ,
         \result_array[9][48] , \result_array[9][47] , \result_array[9][46] ,
         \result_array[9][45] , \result_array[9][44] , \result_array[9][43] ,
         \result_array[9][42] , \result_array[9][41] , \result_array[9][40] ,
         \result_array[9][39] , \result_array[9][38] , \result_array[9][37] ,
         \result_array[9][36] , \result_array[9][35] , \result_array[9][34] ,
         \result_array[9][33] , \result_array[9][32] , \result_array[9][31] ,
         \result_array[9][30] , \result_array[9][29] , \result_array[9][28] ,
         \result_array[9][27] , \result_array[9][26] , \result_array[9][25] ,
         \result_array[9][24] , \result_array[9][23] , \result_array[9][22] ,
         \result_array[9][21] , \result_array[9][20] , \result_array[9][19] ,
         \result_array[9][18] , \result_array[9][17] , \result_array[9][16] ,
         \result_array[9][15] , \result_array[9][14] , \result_array[9][13] ,
         \result_array[9][12] , \result_array[9][11] , \result_array[9][10] ,
         \result_array[9][9] , \result_array[9][8] , \result_array[9][7] ,
         \result_array[9][6] , \result_array[9][5] , \result_array[9][4] ,
         \result_array[9][3] , \result_array[9][2] , \result_array[9][1] ,
         \result_array[9][0] , \result_array[8][63] , \result_array[8][62] ,
         \result_array[8][61] , \result_array[8][60] , \result_array[8][59] ,
         \result_array[8][58] , \result_array[8][57] , \result_array[8][56] ,
         \result_array[8][55] , \result_array[8][54] , \result_array[8][53] ,
         \result_array[8][52] , \result_array[8][51] , \result_array[8][50] ,
         \result_array[8][49] , \result_array[8][48] , \result_array[8][47] ,
         \result_array[8][46] , \result_array[8][45] , \result_array[8][44] ,
         \result_array[8][43] , \result_array[8][42] , \result_array[8][41] ,
         \result_array[8][40] , \result_array[8][39] , \result_array[8][38] ,
         \result_array[8][37] , \result_array[8][36] , \result_array[8][35] ,
         \result_array[8][34] , \result_array[8][33] , \result_array[8][32] ,
         \result_array[8][31] , \result_array[8][30] , \result_array[8][29] ,
         \result_array[8][28] , \result_array[8][27] , \result_array[8][26] ,
         \result_array[8][25] , \result_array[8][24] , \result_array[8][23] ,
         \result_array[8][22] , \result_array[8][21] , \result_array[8][20] ,
         \result_array[8][19] , \result_array[8][18] , \result_array[8][17] ,
         \result_array[8][16] , \result_array[8][15] , \result_array[8][14] ,
         \result_array[8][13] , \result_array[8][12] , \result_array[8][11] ,
         \result_array[8][10] , \result_array[8][9] , \result_array[8][8] ,
         \result_array[8][7] , \result_array[8][6] , \result_array[8][5] ,
         \result_array[8][4] , \result_array[8][3] , \result_array[8][2] ,
         \result_array[8][1] , \result_array[8][0] , n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334;
  wire   [31:0] minus_A;

  Booth_Encoder_0 booth_o_0 ( .i({B[1:0], 1'b0}), .o({\select_array[0][2] , 
        \select_array[0][1] , \select_array[0][0] }) );
  MUX_booth_N64_0 mux_0_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n311, n302, n303, 
        n302, n302, n303, n303, n303, n304, n303, n303, n304, n306, n304, n304, 
        n304, n305, n306, n306, n306, n306, n306, n308, n308, n308, n308, n308, 
        n308, n308, n308, n310, n310, n310, n278, n276, n273, n271, n268, n266, 
        n263, n261, n258, n256, n253, n251, n248, n246, n243, n241, n238, n237, 
        n235, n234, n71, n229, n228, n227, n224, n223, n76, n220, n96, n216, 
        n97}), .C({n173, n182, n181, n180, n180, n180, n181, n180, n180, n180, 
        n181, n180, n179, n179, n180, n179, n178, n177, n177, n177, n177, n177, 
        n177, n177, n177, n175, n175, n175, n210, n205, n204, n209, 
        minus_A[31:30], n154, n151, minus_A[27], n148, n146, n143, n141, 
        minus_A[22:20], n134, n58, n131, minus_A[16], n126, n125, 
        minus_A[13:12], n59, n118, n116, minus_A[8], n61, n112, minus_A[5], 
        n108, n105, n102, n99, n212}), .D({n299, n299, n299, n299, n299, n299, 
        n299, n299, n298, n298, n298, n298, n298, n298, n298, n298, n298, n298, 
        n297, n297, n297, n297, n297, n297, n297, n296, n296, n296, n300, n296, 
        n295, n295, n277, n275, n272, n270, n267, n265, n262, n260, n257, n255, 
        n252, n250, n247, n245, n242, n240, n238, n236, n235, n233, n72, n229, 
        n228, n226, A[6], n222, n78, n219, n96, n215, n97, 1'b0}), .E({n183, 
        n184, n184, n184, n184, n184, n185, n185, n185, n185, n185, n185, n185, 
        n185, n186, n186, n186, n186, n186, n186, n186, n186, n186, n187, n187, 
        n187, n187, n183, n187, n188, n188, n161, minus_A[30], n154, n151, 
        minus_A[27:25], n143, minus_A[23:16], n128, minus_A[14:10], n116, 
        minus_A[8:4], n107, n104, n101, n214, 1'b0}), .sel({
        \select_array[0][2] , \select_array[0][1] , \select_array[0][0] }), 
        .Y({\result_array[0][63] , \result_array[0][62] , 
        \result_array[0][61] , \result_array[0][60] , \result_array[0][59] , 
        \result_array[0][58] , \result_array[0][57] , \result_array[0][56] , 
        \result_array[0][55] , \result_array[0][54] , \result_array[0][53] , 
        \result_array[0][52] , \result_array[0][51] , \result_array[0][50] , 
        \result_array[0][49] , \result_array[0][48] , \result_array[0][47] , 
        \result_array[0][46] , \result_array[0][45] , \result_array[0][44] , 
        \result_array[0][43] , \result_array[0][42] , \result_array[0][41] , 
        \result_array[0][40] , \result_array[0][39] , \result_array[0][38] , 
        \result_array[0][37] , \result_array[0][36] , \result_array[0][35] , 
        \result_array[0][34] , \result_array[0][33] , \result_array[0][32] , 
        \result_array[0][31] , \result_array[0][30] , \result_array[0][29] , 
        \result_array[0][28] , \result_array[0][27] , \result_array[0][26] , 
        \result_array[0][25] , \result_array[0][24] , \result_array[0][23] , 
        \result_array[0][22] , \result_array[0][21] , \result_array[0][20] , 
        \result_array[0][19] , \result_array[0][18] , \result_array[0][17] , 
        \result_array[0][16] , \result_array[0][15] , \result_array[0][14] , 
        \result_array[0][13] , \result_array[0][12] , \result_array[0][11] , 
        \result_array[0][10] , \result_array[0][9] , \result_array[0][8] , 
        \result_array[0][7] , \result_array[0][6] , \result_array[0][5] , 
        \result_array[0][4] , \result_array[0][3] , \result_array[0][2] , 
        \result_array[0][1] , \result_array[0][0] }) );
  Booth_Encoder_15 booth_j_1 ( .i(B[3:1]), .o({\select_array[1][2] , 
        \select_array[1][1] , \select_array[1][0] }) );
  MUX_booth_N64_15 mux_j_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n310, n310, 
        n310, n310, n310, n311, n311, n311, n311, n302, n310, n310, n310, n310, 
        n310, n309, n309, n309, n309, n309, n309, n309, n309, n309, n309, n309, 
        n309, n309, n308, n308, n308, n278, n276, n273, n271, n268, n266, n263, 
        n261, n258, n256, n253, n251, n248, n246, n243, n241, n238, n237, n235, 
        n234, n72, n230, n228, n227, n224, n223, n79, n220, n96, n98, A[0], 
        1'b0, 1'b0}), .C({n173, n173, n173, n174, n173, n173, n173, n173, n173, 
        n172, n174, n174, n178, n174, n174, n174, n174, n174, n174, n174, n174, 
        n174, n175, n175, n175, n175, n175, n175, n175, n175, n160, n158, n154, 
        n152, n94, n148, n147, n144, n141, minus_A[22:21], n136, n134, 
        minus_A[18], n132, n129, n127, n125, n64, n121, n119, minus_A[10], 
        n116, n115, n63, n112, minus_A[5], n109, n106, n103, n100, n213, 1'b0, 
        1'b0}), .D({n292, n292, n292, n292, n292, n292, n292, n292, n292, n292, 
        n292, n292, n293, n293, n293, n293, n293, n293, n293, n293, n293, n293, 
        n293, n293, n294, n294, n294, n294, n279, n279, n277, n275, n272, n270, 
        n267, n265, n262, n260, n257, n255, n252, n250, n247, n245, n242, n240, 
        n238, n236, n235, n233, n72, n230, n228, n226, A[6], n222, n77, n219, 
        n96, n217, n67, 1'b0, 1'b0, 1'b0}), .E({n191, n191, n191, n191, n191, 
        n191, n191, n191, n190, n190, n190, n190, n190, n190, n190, n190, n190, 
        n190, n190, n190, n189, n189, n189, n189, n189, n189, n196, n187, n189, 
        n161, n157, n155, n151, n94, n148, minus_A[25], n143, n141, 
        minus_A[22:20], n134, minus_A[18:16], n128, n125, minus_A[13:8], n61, 
        n112, minus_A[5:4], n107, n104, n101, n214, 1'b0, 1'b0, 1'b0}), .sel({
        \select_array[1][2] , \select_array[1][1] , \select_array[1][0] }), 
        .Y({\array_mux_out[1][63] , \array_mux_out[1][62] , 
        \array_mux_out[1][61] , \array_mux_out[1][60] , \array_mux_out[1][59] , 
        \array_mux_out[1][58] , \array_mux_out[1][57] , \array_mux_out[1][56] , 
        \array_mux_out[1][55] , \array_mux_out[1][54] , \array_mux_out[1][53] , 
        \array_mux_out[1][52] , \array_mux_out[1][51] , \array_mux_out[1][50] , 
        \array_mux_out[1][49] , \array_mux_out[1][48] , \array_mux_out[1][47] , 
        \array_mux_out[1][46] , \array_mux_out[1][45] , \array_mux_out[1][44] , 
        \array_mux_out[1][43] , \array_mux_out[1][42] , \array_mux_out[1][41] , 
        \array_mux_out[1][40] , \array_mux_out[1][39] , \array_mux_out[1][38] , 
        \array_mux_out[1][37] , \array_mux_out[1][36] , \array_mux_out[1][35] , 
        \array_mux_out[1][34] , \array_mux_out[1][33] , \array_mux_out[1][32] , 
        \array_mux_out[1][31] , \array_mux_out[1][30] , \array_mux_out[1][29] , 
        \array_mux_out[1][28] , \array_mux_out[1][27] , \array_mux_out[1][26] , 
        \array_mux_out[1][25] , \array_mux_out[1][24] , \array_mux_out[1][23] , 
        \array_mux_out[1][22] , \array_mux_out[1][21] , \array_mux_out[1][20] , 
        \array_mux_out[1][19] , \array_mux_out[1][18] , \array_mux_out[1][17] , 
        \array_mux_out[1][16] , \array_mux_out[1][15] , \array_mux_out[1][14] , 
        \array_mux_out[1][13] , \array_mux_out[1][12] , \array_mux_out[1][11] , 
        \array_mux_out[1][10] , \array_mux_out[1][9] , \array_mux_out[1][8] , 
        \array_mux_out[1][7] , \array_mux_out[1][6] , \array_mux_out[1][5] , 
        \array_mux_out[1][4] , \array_mux_out[1][3] , \array_mux_out[1][2] , 
        \array_mux_out[1][1] , \array_mux_out[1][0] }) );
  P4_ADDER_N64_0 adder_1 ( .A({\array_mux_out[1][63] , \array_mux_out[1][62] , 
        \array_mux_out[1][61] , \array_mux_out[1][60] , \array_mux_out[1][59] , 
        \array_mux_out[1][58] , \array_mux_out[1][57] , \array_mux_out[1][56] , 
        \array_mux_out[1][55] , \array_mux_out[1][54] , \array_mux_out[1][53] , 
        \array_mux_out[1][52] , \array_mux_out[1][51] , \array_mux_out[1][50] , 
        \array_mux_out[1][49] , \array_mux_out[1][48] , \array_mux_out[1][47] , 
        \array_mux_out[1][46] , \array_mux_out[1][45] , \array_mux_out[1][44] , 
        \array_mux_out[1][43] , \array_mux_out[1][42] , \array_mux_out[1][41] , 
        \array_mux_out[1][40] , \array_mux_out[1][39] , \array_mux_out[1][38] , 
        \array_mux_out[1][37] , \array_mux_out[1][36] , \array_mux_out[1][35] , 
        \array_mux_out[1][34] , \array_mux_out[1][33] , \array_mux_out[1][32] , 
        \array_mux_out[1][31] , \array_mux_out[1][30] , \array_mux_out[1][29] , 
        \array_mux_out[1][28] , \array_mux_out[1][27] , \array_mux_out[1][26] , 
        \array_mux_out[1][25] , \array_mux_out[1][24] , \array_mux_out[1][23] , 
        \array_mux_out[1][22] , \array_mux_out[1][21] , \array_mux_out[1][20] , 
        \array_mux_out[1][19] , \array_mux_out[1][18] , \array_mux_out[1][17] , 
        \array_mux_out[1][16] , \array_mux_out[1][15] , \array_mux_out[1][14] , 
        \array_mux_out[1][13] , \array_mux_out[1][12] , \array_mux_out[1][11] , 
        \array_mux_out[1][10] , \array_mux_out[1][9] , \array_mux_out[1][8] , 
        \array_mux_out[1][7] , \array_mux_out[1][6] , \array_mux_out[1][5] , 
        \array_mux_out[1][4] , \array_mux_out[1][3] , \array_mux_out[1][2] , 
        \array_mux_out[1][1] , \array_mux_out[1][0] }), .B({
        \result_array[0][63] , \result_array[0][62] , \result_array[0][61] , 
        \result_array[0][60] , \result_array[0][59] , \result_array[0][58] , 
        \result_array[0][57] , \result_array[0][56] , \result_array[0][55] , 
        \result_array[0][54] , \result_array[0][53] , \result_array[0][52] , 
        \result_array[0][51] , \result_array[0][50] , \result_array[0][49] , 
        \result_array[0][48] , \result_array[0][47] , \result_array[0][46] , 
        \result_array[0][45] , \result_array[0][44] , \result_array[0][43] , 
        \result_array[0][42] , \result_array[0][41] , \result_array[0][40] , 
        \result_array[0][39] , \result_array[0][38] , \result_array[0][37] , 
        \result_array[0][36] , \result_array[0][35] , \result_array[0][34] , 
        \result_array[0][33] , \result_array[0][32] , \result_array[0][31] , 
        \result_array[0][30] , \result_array[0][29] , \result_array[0][28] , 
        \result_array[0][27] , \result_array[0][26] , \result_array[0][25] , 
        \result_array[0][24] , \result_array[0][23] , \result_array[0][22] , 
        \result_array[0][21] , \result_array[0][20] , \result_array[0][19] , 
        \result_array[0][18] , \result_array[0][17] , \result_array[0][16] , 
        \result_array[0][15] , \result_array[0][14] , \result_array[0][13] , 
        \result_array[0][12] , \result_array[0][11] , \result_array[0][10] , 
        \result_array[0][9] , \result_array[0][8] , \result_array[0][7] , 
        \result_array[0][6] , \result_array[0][5] , \result_array[0][4] , 
        \result_array[0][3] , \result_array[0][2] , \result_array[0][1] , 
        \result_array[0][0] }), .Cin(1'b0), .S({\result_array[1][63] , 
        \result_array[1][62] , \result_array[1][61] , \result_array[1][60] , 
        \result_array[1][59] , \result_array[1][58] , \result_array[1][57] , 
        \result_array[1][56] , \result_array[1][55] , \result_array[1][54] , 
        \result_array[1][53] , \result_array[1][52] , \result_array[1][51] , 
        \result_array[1][50] , \result_array[1][49] , \result_array[1][48] , 
        \result_array[1][47] , \result_array[1][46] , \result_array[1][45] , 
        \result_array[1][44] , \result_array[1][43] , \result_array[1][42] , 
        \result_array[1][41] , \result_array[1][40] , \result_array[1][39] , 
        \result_array[1][38] , \result_array[1][37] , \result_array[1][36] , 
        \result_array[1][35] , \result_array[1][34] , \result_array[1][33] , 
        \result_array[1][32] , \result_array[1][31] , \result_array[1][30] , 
        \result_array[1][29] , \result_array[1][28] , \result_array[1][27] , 
        \result_array[1][26] , \result_array[1][25] , \result_array[1][24] , 
        \result_array[1][23] , \result_array[1][22] , \result_array[1][21] , 
        \result_array[1][20] , \result_array[1][19] , \result_array[1][18] , 
        \result_array[1][17] , \result_array[1][16] , \result_array[1][15] , 
        \result_array[1][14] , \result_array[1][13] , \result_array[1][12] , 
        \result_array[1][11] , \result_array[1][10] , \result_array[1][9] , 
        \result_array[1][8] , \result_array[1][7] , \result_array[1][6] , 
        \result_array[1][5] , \result_array[1][4] , \result_array[1][3] , 
        \result_array[1][2] , \result_array[1][1] , \result_array[1][0] }) );
  Booth_Encoder_14 booth_j_2 ( .i(B[5:3]), .o({\select_array[2][2] , 
        \select_array[2][1] , \select_array[2][0] }) );
  MUX_booth_N64_14 mux_j_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n305, n305, 
        n305, n305, n305, n305, n305, n306, n306, n306, n306, n306, n306, n306, 
        n307, n307, n307, n307, n307, n307, n307, n307, n307, n307, n307, n307, 
        n307, n308, n308, n278, n276, n273, n271, n268, n266, n263, n261, n258, 
        n256, n253, n251, n248, n246, n243, n241, n238, n237, n235, n234, n71, 
        n229, n228, n227, n224, n223, n80, n220, n96, n217, n67, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n179, n178, n178, n178, n178, n178, n178, n178, n178, 
        n178, n178, n177, n177, n177, n177, n176, n176, n176, n176, n176, n176, 
        n176, n176, n176, n176, n176, n176, n175, n160, n158, n155, n153, n94, 
        n149, n147, n145, n142, n139, n70, n69, n135, n133, n132, n129, n127, 
        n124, n122, n121, n119, n118, n116, n114, n113, n111, n110, n109, n106, 
        n103, n100, n213, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n289, n289, n289, n289, 
        n290, n290, n290, n290, n290, n290, n290, n290, n290, n290, n290, n290, 
        n291, n291, n291, n291, n291, n291, n291, n291, n291, n291, n291, n291, 
        n277, n274, n272, n269, n267, n264, n262, n259, n257, n254, n252, n249, 
        n247, n244, n242, n239, n238, n236, n235, n232, n71, n229, n228, n225, 
        A[6], n221, n81, n218, n96, n216, n67, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .E({n193, n193, n193, n193, n193, n193, n193, n193, n193, n193, n193, 
        n192, n192, n192, n192, n192, n192, n192, n192, n192, n192, n192, n192, 
        n191, n191, n191, n191, n161, n157, n155, n153, n94, n149, n147, n144, 
        n142, n140, n70, n137, n135, n133, n62, n130, n128, n124, n123, n120, 
        n119, n117, n91, n114, n113, n111, n110, n109, n107, n104, n101, n214, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[2][2] , 
        \select_array[2][1] , \select_array[2][0] }), .Y({
        \array_mux_out[2][63] , \array_mux_out[2][62] , \array_mux_out[2][61] , 
        \array_mux_out[2][60] , \array_mux_out[2][59] , \array_mux_out[2][58] , 
        \array_mux_out[2][57] , \array_mux_out[2][56] , \array_mux_out[2][55] , 
        \array_mux_out[2][54] , \array_mux_out[2][53] , \array_mux_out[2][52] , 
        \array_mux_out[2][51] , \array_mux_out[2][50] , \array_mux_out[2][49] , 
        \array_mux_out[2][48] , \array_mux_out[2][47] , \array_mux_out[2][46] , 
        \array_mux_out[2][45] , \array_mux_out[2][44] , \array_mux_out[2][43] , 
        \array_mux_out[2][42] , \array_mux_out[2][41] , \array_mux_out[2][40] , 
        \array_mux_out[2][39] , \array_mux_out[2][38] , \array_mux_out[2][37] , 
        \array_mux_out[2][36] , \array_mux_out[2][35] , \array_mux_out[2][34] , 
        \array_mux_out[2][33] , \array_mux_out[2][32] , \array_mux_out[2][31] , 
        \array_mux_out[2][30] , \array_mux_out[2][29] , \array_mux_out[2][28] , 
        \array_mux_out[2][27] , \array_mux_out[2][26] , \array_mux_out[2][25] , 
        \array_mux_out[2][24] , \array_mux_out[2][23] , \array_mux_out[2][22] , 
        \array_mux_out[2][21] , \array_mux_out[2][20] , \array_mux_out[2][19] , 
        \array_mux_out[2][18] , \array_mux_out[2][17] , \array_mux_out[2][16] , 
        \array_mux_out[2][15] , \array_mux_out[2][14] , \array_mux_out[2][13] , 
        \array_mux_out[2][12] , \array_mux_out[2][11] , \array_mux_out[2][10] , 
        \array_mux_out[2][9] , \array_mux_out[2][8] , \array_mux_out[2][7] , 
        \array_mux_out[2][6] , \array_mux_out[2][5] , \array_mux_out[2][4] , 
        \array_mux_out[2][3] , \array_mux_out[2][2] , \array_mux_out[2][1] , 
        \array_mux_out[2][0] }) );
  P4_ADDER_N64_14 adder_2 ( .A({\array_mux_out[2][63] , \array_mux_out[2][62] , 
        \array_mux_out[2][61] , \array_mux_out[2][60] , \array_mux_out[2][59] , 
        \array_mux_out[2][58] , \array_mux_out[2][57] , \array_mux_out[2][56] , 
        \array_mux_out[2][55] , \array_mux_out[2][54] , \array_mux_out[2][53] , 
        \array_mux_out[2][52] , \array_mux_out[2][51] , \array_mux_out[2][50] , 
        \array_mux_out[2][49] , \array_mux_out[2][48] , \array_mux_out[2][47] , 
        \array_mux_out[2][46] , \array_mux_out[2][45] , \array_mux_out[2][44] , 
        \array_mux_out[2][43] , \array_mux_out[2][42] , \array_mux_out[2][41] , 
        \array_mux_out[2][40] , \array_mux_out[2][39] , \array_mux_out[2][38] , 
        \array_mux_out[2][37] , \array_mux_out[2][36] , \array_mux_out[2][35] , 
        \array_mux_out[2][34] , \array_mux_out[2][33] , \array_mux_out[2][32] , 
        \array_mux_out[2][31] , \array_mux_out[2][30] , \array_mux_out[2][29] , 
        \array_mux_out[2][28] , \array_mux_out[2][27] , \array_mux_out[2][26] , 
        \array_mux_out[2][25] , \array_mux_out[2][24] , \array_mux_out[2][23] , 
        \array_mux_out[2][22] , \array_mux_out[2][21] , \array_mux_out[2][20] , 
        \array_mux_out[2][19] , \array_mux_out[2][18] , \array_mux_out[2][17] , 
        \array_mux_out[2][16] , \array_mux_out[2][15] , \array_mux_out[2][14] , 
        \array_mux_out[2][13] , \array_mux_out[2][12] , \array_mux_out[2][11] , 
        \array_mux_out[2][10] , \array_mux_out[2][9] , \array_mux_out[2][8] , 
        \array_mux_out[2][7] , \array_mux_out[2][6] , \array_mux_out[2][5] , 
        \array_mux_out[2][4] , \array_mux_out[2][3] , \array_mux_out[2][2] , 
        \array_mux_out[2][1] , \array_mux_out[2][0] }), .B({
        \result_array[1][63] , \result_array[1][62] , \result_array[1][61] , 
        \result_array[1][60] , \result_array[1][59] , \result_array[1][58] , 
        \result_array[1][57] , \result_array[1][56] , \result_array[1][55] , 
        \result_array[1][54] , \result_array[1][53] , \result_array[1][52] , 
        \result_array[1][51] , \result_array[1][50] , \result_array[1][49] , 
        \result_array[1][48] , \result_array[1][47] , \result_array[1][46] , 
        \result_array[1][45] , \result_array[1][44] , \result_array[1][43] , 
        \result_array[1][42] , \result_array[1][41] , \result_array[1][40] , 
        \result_array[1][39] , \result_array[1][38] , \result_array[1][37] , 
        \result_array[1][36] , \result_array[1][35] , \result_array[1][34] , 
        \result_array[1][33] , \result_array[1][32] , \result_array[1][31] , 
        \result_array[1][30] , \result_array[1][29] , \result_array[1][28] , 
        \result_array[1][27] , \result_array[1][26] , \result_array[1][25] , 
        \result_array[1][24] , \result_array[1][23] , \result_array[1][22] , 
        \result_array[1][21] , \result_array[1][20] , \result_array[1][19] , 
        \result_array[1][18] , \result_array[1][17] , \result_array[1][16] , 
        \result_array[1][15] , \result_array[1][14] , \result_array[1][13] , 
        \result_array[1][12] , \result_array[1][11] , \result_array[1][10] , 
        \result_array[1][9] , \result_array[1][8] , \result_array[1][7] , 
        \result_array[1][6] , \result_array[1][5] , \result_array[1][4] , 
        \result_array[1][3] , \result_array[1][2] , \result_array[1][1] , 
        \result_array[1][0] }), .Cin(1'b0), .S({\result_array[2][63] , 
        \result_array[2][62] , \result_array[2][61] , \result_array[2][60] , 
        \result_array[2][59] , \result_array[2][58] , \result_array[2][57] , 
        \result_array[2][56] , \result_array[2][55] , \result_array[2][54] , 
        \result_array[2][53] , \result_array[2][52] , \result_array[2][51] , 
        \result_array[2][50] , \result_array[2][49] , \result_array[2][48] , 
        \result_array[2][47] , \result_array[2][46] , \result_array[2][45] , 
        \result_array[2][44] , \result_array[2][43] , \result_array[2][42] , 
        \result_array[2][41] , \result_array[2][40] , \result_array[2][39] , 
        \result_array[2][38] , \result_array[2][37] , \result_array[2][36] , 
        \result_array[2][35] , \result_array[2][34] , \result_array[2][33] , 
        \result_array[2][32] , \result_array[2][31] , \result_array[2][30] , 
        \result_array[2][29] , \result_array[2][28] , \result_array[2][27] , 
        \result_array[2][26] , \result_array[2][25] , \result_array[2][24] , 
        \result_array[2][23] , \result_array[2][22] , \result_array[2][21] , 
        \result_array[2][20] , \result_array[2][19] , \result_array[2][18] , 
        \result_array[2][17] , \result_array[2][16] , \result_array[2][15] , 
        \result_array[2][14] , \result_array[2][13] , \result_array[2][12] , 
        \result_array[2][11] , \result_array[2][10] , \result_array[2][9] , 
        \result_array[2][8] , \result_array[2][7] , \result_array[2][6] , 
        \result_array[2][5] , \result_array[2][4] , \result_array[2][3] , 
        \result_array[2][2] , \result_array[2][1] , \result_array[2][0] }) );
  Booth_Encoder_13 booth_j_3 ( .i(B[7:5]), .o({\select_array[3][2] , 
        \select_array[3][1] , \select_array[3][0] }) );
  MUX_booth_N64_13 mux_j_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n323, n323, 
        n323, n323, n323, n321, n305, n301, n302, n301, n302, n301, n303, n301, 
        n302, n302, n302, n303, n302, n303, n302, n304, n302, n303, n305, n303, 
        n304, n278, n276, n273, n271, n268, n266, n263, n261, n258, n256, n253, 
        n251, n248, n246, n243, n241, n238, n237, n235, n234, n72, n230, n228, 
        n227, n224, n223, n84, n220, n96, n216, n95, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n164, n164, n164, n164, n164, n164, n164, n164, n164, 
        n170, n179, n182, n182, n182, n182, n181, n182, n182, n181, n182, n181, 
        n181, n181, n181, n181, n181, n160, n157, n156, n152, n94, n149, n147, 
        n145, n142, n139, n138, n68, n135, n133, n132, n129, n127, n124, n123, 
        n121, n119, n118, n116, n114, n113, n111, n110, n109, n106, n103, n100, 
        n213, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n287, n287, n287, n287, 
        n287, n287, n288, n288, n288, n288, n288, n288, n288, n288, n288, n288, 
        n288, n288, n289, n289, n289, n289, n289, n289, n289, n289, n277, n274, 
        n272, n269, n267, n264, n262, n259, n257, n254, n252, n249, n247, n244, 
        n242, n239, n238, n236, n235, n232, n72, n230, n228, n225, A[6], n221, 
        n82, n218, n96, n216, n95, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .E({n195, n195, n195, n195, n195, n195, n195, n195, n195, n195, n195, 
        n195, n194, n194, n194, n194, n194, n194, n194, n194, n194, n194, n194, 
        n194, n193, n161, n157, n155, n153, n150, n149, n147, n144, n142, n140, 
        n138, n137, n135, n133, n62, n130, n128, n124, n122, n121, n119, n117, 
        n91, n115, n113, n65, n110, n109, n107, n104, n101, n214, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[3][2] , 
        \select_array[3][1] , \select_array[3][0] }), .Y({
        \array_mux_out[3][63] , \array_mux_out[3][62] , \array_mux_out[3][61] , 
        \array_mux_out[3][60] , \array_mux_out[3][59] , \array_mux_out[3][58] , 
        \array_mux_out[3][57] , \array_mux_out[3][56] , \array_mux_out[3][55] , 
        \array_mux_out[3][54] , \array_mux_out[3][53] , \array_mux_out[3][52] , 
        \array_mux_out[3][51] , \array_mux_out[3][50] , \array_mux_out[3][49] , 
        \array_mux_out[3][48] , \array_mux_out[3][47] , \array_mux_out[3][46] , 
        \array_mux_out[3][45] , \array_mux_out[3][44] , \array_mux_out[3][43] , 
        \array_mux_out[3][42] , \array_mux_out[3][41] , \array_mux_out[3][40] , 
        \array_mux_out[3][39] , \array_mux_out[3][38] , \array_mux_out[3][37] , 
        \array_mux_out[3][36] , \array_mux_out[3][35] , \array_mux_out[3][34] , 
        \array_mux_out[3][33] , \array_mux_out[3][32] , \array_mux_out[3][31] , 
        \array_mux_out[3][30] , \array_mux_out[3][29] , \array_mux_out[3][28] , 
        \array_mux_out[3][27] , \array_mux_out[3][26] , \array_mux_out[3][25] , 
        \array_mux_out[3][24] , \array_mux_out[3][23] , \array_mux_out[3][22] , 
        \array_mux_out[3][21] , \array_mux_out[3][20] , \array_mux_out[3][19] , 
        \array_mux_out[3][18] , \array_mux_out[3][17] , \array_mux_out[3][16] , 
        \array_mux_out[3][15] , \array_mux_out[3][14] , \array_mux_out[3][13] , 
        \array_mux_out[3][12] , \array_mux_out[3][11] , \array_mux_out[3][10] , 
        \array_mux_out[3][9] , \array_mux_out[3][8] , \array_mux_out[3][7] , 
        \array_mux_out[3][6] , \array_mux_out[3][5] , \array_mux_out[3][4] , 
        \array_mux_out[3][3] , \array_mux_out[3][2] , \array_mux_out[3][1] , 
        \array_mux_out[3][0] }) );
  P4_ADDER_N64_13 adder_3 ( .A({\array_mux_out[3][63] , \array_mux_out[3][62] , 
        \array_mux_out[3][61] , \array_mux_out[3][60] , \array_mux_out[3][59] , 
        \array_mux_out[3][58] , \array_mux_out[3][57] , \array_mux_out[3][56] , 
        \array_mux_out[3][55] , \array_mux_out[3][54] , \array_mux_out[3][53] , 
        \array_mux_out[3][52] , \array_mux_out[3][51] , \array_mux_out[3][50] , 
        \array_mux_out[3][49] , \array_mux_out[3][48] , \array_mux_out[3][47] , 
        \array_mux_out[3][46] , \array_mux_out[3][45] , \array_mux_out[3][44] , 
        \array_mux_out[3][43] , \array_mux_out[3][42] , \array_mux_out[3][41] , 
        \array_mux_out[3][40] , \array_mux_out[3][39] , \array_mux_out[3][38] , 
        \array_mux_out[3][37] , \array_mux_out[3][36] , \array_mux_out[3][35] , 
        \array_mux_out[3][34] , \array_mux_out[3][33] , \array_mux_out[3][32] , 
        \array_mux_out[3][31] , \array_mux_out[3][30] , \array_mux_out[3][29] , 
        \array_mux_out[3][28] , \array_mux_out[3][27] , \array_mux_out[3][26] , 
        \array_mux_out[3][25] , \array_mux_out[3][24] , \array_mux_out[3][23] , 
        \array_mux_out[3][22] , \array_mux_out[3][21] , \array_mux_out[3][20] , 
        \array_mux_out[3][19] , \array_mux_out[3][18] , \array_mux_out[3][17] , 
        \array_mux_out[3][16] , \array_mux_out[3][15] , \array_mux_out[3][14] , 
        \array_mux_out[3][13] , \array_mux_out[3][12] , \array_mux_out[3][11] , 
        \array_mux_out[3][10] , \array_mux_out[3][9] , \array_mux_out[3][8] , 
        \array_mux_out[3][7] , \array_mux_out[3][6] , \array_mux_out[3][5] , 
        \array_mux_out[3][4] , \array_mux_out[3][3] , \array_mux_out[3][2] , 
        \array_mux_out[3][1] , \array_mux_out[3][0] }), .B({
        \result_array[2][63] , \result_array[2][62] , \result_array[2][61] , 
        \result_array[2][60] , \result_array[2][59] , \result_array[2][58] , 
        \result_array[2][57] , \result_array[2][56] , \result_array[2][55] , 
        \result_array[2][54] , \result_array[2][53] , \result_array[2][52] , 
        \result_array[2][51] , \result_array[2][50] , \result_array[2][49] , 
        \result_array[2][48] , \result_array[2][47] , \result_array[2][46] , 
        \result_array[2][45] , \result_array[2][44] , \result_array[2][43] , 
        \result_array[2][42] , \result_array[2][41] , \result_array[2][40] , 
        \result_array[2][39] , \result_array[2][38] , \result_array[2][37] , 
        \result_array[2][36] , \result_array[2][35] , \result_array[2][34] , 
        \result_array[2][33] , \result_array[2][32] , \result_array[2][31] , 
        \result_array[2][30] , \result_array[2][29] , \result_array[2][28] , 
        \result_array[2][27] , \result_array[2][26] , \result_array[2][25] , 
        \result_array[2][24] , \result_array[2][23] , \result_array[2][22] , 
        \result_array[2][21] , \result_array[2][20] , \result_array[2][19] , 
        \result_array[2][18] , \result_array[2][17] , \result_array[2][16] , 
        \result_array[2][15] , \result_array[2][14] , \result_array[2][13] , 
        \result_array[2][12] , \result_array[2][11] , \result_array[2][10] , 
        \result_array[2][9] , \result_array[2][8] , \result_array[2][7] , 
        \result_array[2][6] , \result_array[2][5] , \result_array[2][4] , 
        \result_array[2][3] , \result_array[2][2] , \result_array[2][1] , 
        \result_array[2][0] }), .Cin(1'b0), .S({\result_array[3][63] , 
        \result_array[3][62] , \result_array[3][61] , \result_array[3][60] , 
        \result_array[3][59] , \result_array[3][58] , \result_array[3][57] , 
        \result_array[3][56] , \result_array[3][55] , \result_array[3][54] , 
        \result_array[3][53] , \result_array[3][52] , \result_array[3][51] , 
        \result_array[3][50] , \result_array[3][49] , \result_array[3][48] , 
        \result_array[3][47] , \result_array[3][46] , \result_array[3][45] , 
        \result_array[3][44] , \result_array[3][43] , \result_array[3][42] , 
        \result_array[3][41] , \result_array[3][40] , \result_array[3][39] , 
        \result_array[3][38] , \result_array[3][37] , \result_array[3][36] , 
        \result_array[3][35] , \result_array[3][34] , \result_array[3][33] , 
        \result_array[3][32] , \result_array[3][31] , \result_array[3][30] , 
        \result_array[3][29] , \result_array[3][28] , \result_array[3][27] , 
        \result_array[3][26] , \result_array[3][25] , \result_array[3][24] , 
        \result_array[3][23] , \result_array[3][22] , \result_array[3][21] , 
        \result_array[3][20] , \result_array[3][19] , \result_array[3][18] , 
        \result_array[3][17] , \result_array[3][16] , \result_array[3][15] , 
        \result_array[3][14] , \result_array[3][13] , \result_array[3][12] , 
        \result_array[3][11] , \result_array[3][10] , \result_array[3][9] , 
        \result_array[3][8] , \result_array[3][7] , \result_array[3][6] , 
        \result_array[3][5] , \result_array[3][4] , \result_array[3][3] , 
        \result_array[3][2] , \result_array[3][1] , \result_array[3][0] }) );
  Booth_Encoder_12 booth_j_4 ( .i(B[9:7]), .o({\select_array[4][2] , 
        \select_array[4][1] , \select_array[4][0] }) );
  MUX_booth_N64_12 mux_j_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n320, n320, 
        n320, n320, n320, n320, n320, n321, n321, n321, n321, n321, n321, n321, 
        n321, n321, n321, n321, n321, n322, n322, n322, n322, n322, n322, n278, 
        n276, n273, n271, n268, n266, n263, n261, n258, n256, n253, n251, n248, 
        n246, n243, n241, n238, n237, n235, n234, n72, n230, n228, n227, n224, 
        n223, n83, n220, n96, n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n167, n167, n167, n167, n167, n167, n167, n167, n167, 
        n167, n166, n166, n166, n166, n166, n166, n166, n166, n166, n166, n166, 
        n166, n165, n165, n160, n158, n155, n153, n150, n149, n147, n144, n142, 
        n139, n70, n68, n135, n133, n132, n130, n127, n124, n123, n120, n119, 
        n118, n116, n114, n113, n111, n110, n109, n106, n103, n100, n213, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n285, n285, n285, n285, 
        n285, n285, n285, n286, n286, n286, n286, n286, n286, n286, n286, n286, 
        n286, n286, n287, n287, n287, n287, n287, n287, n277, n274, n272, n269, 
        n267, n264, n262, n259, n257, n254, n252, n249, n247, n244, n242, n239, 
        n238, n236, n235, n232, n71, n229, n228, n225, A[6], n221, n86, n218, 
        n96, n216, n95, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .E({n197, n197, n197, n197, n197, n197, n197, n197, n197, n197, n197, 
        n197, n180, n196, n196, n196, n196, n196, n196, n196, n196, n196, n196, 
        n160, n158, n155, n153, n150, n149, n147, n144, n142, n140, n70, n69, 
        n135, n133, n132, n130, n127, n124, n122, n120, n119, n117, n116, n114, 
        n113, n111, n110, n109, n106, n103, n100, n213, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[4][2] , 
        \select_array[4][1] , \select_array[4][0] }), .Y({
        \array_mux_out[4][63] , \array_mux_out[4][62] , \array_mux_out[4][61] , 
        \array_mux_out[4][60] , \array_mux_out[4][59] , \array_mux_out[4][58] , 
        \array_mux_out[4][57] , \array_mux_out[4][56] , \array_mux_out[4][55] , 
        \array_mux_out[4][54] , \array_mux_out[4][53] , \array_mux_out[4][52] , 
        \array_mux_out[4][51] , \array_mux_out[4][50] , \array_mux_out[4][49] , 
        \array_mux_out[4][48] , \array_mux_out[4][47] , \array_mux_out[4][46] , 
        \array_mux_out[4][45] , \array_mux_out[4][44] , \array_mux_out[4][43] , 
        \array_mux_out[4][42] , \array_mux_out[4][41] , \array_mux_out[4][40] , 
        \array_mux_out[4][39] , \array_mux_out[4][38] , \array_mux_out[4][37] , 
        \array_mux_out[4][36] , \array_mux_out[4][35] , \array_mux_out[4][34] , 
        \array_mux_out[4][33] , \array_mux_out[4][32] , \array_mux_out[4][31] , 
        \array_mux_out[4][30] , \array_mux_out[4][29] , \array_mux_out[4][28] , 
        \array_mux_out[4][27] , \array_mux_out[4][26] , \array_mux_out[4][25] , 
        \array_mux_out[4][24] , \array_mux_out[4][23] , \array_mux_out[4][22] , 
        \array_mux_out[4][21] , \array_mux_out[4][20] , \array_mux_out[4][19] , 
        \array_mux_out[4][18] , \array_mux_out[4][17] , \array_mux_out[4][16] , 
        \array_mux_out[4][15] , \array_mux_out[4][14] , \array_mux_out[4][13] , 
        \array_mux_out[4][12] , \array_mux_out[4][11] , \array_mux_out[4][10] , 
        \array_mux_out[4][9] , \array_mux_out[4][8] , \array_mux_out[4][7] , 
        \array_mux_out[4][6] , \array_mux_out[4][5] , \array_mux_out[4][4] , 
        \array_mux_out[4][3] , \array_mux_out[4][2] , \array_mux_out[4][1] , 
        \array_mux_out[4][0] }) );
  P4_ADDER_N64_12 adder_4 ( .A({\array_mux_out[4][63] , \array_mux_out[4][62] , 
        \array_mux_out[4][61] , \array_mux_out[4][60] , \array_mux_out[4][59] , 
        \array_mux_out[4][58] , \array_mux_out[4][57] , \array_mux_out[4][56] , 
        \array_mux_out[4][55] , \array_mux_out[4][54] , \array_mux_out[4][53] , 
        \array_mux_out[4][52] , \array_mux_out[4][51] , \array_mux_out[4][50] , 
        \array_mux_out[4][49] , \array_mux_out[4][48] , \array_mux_out[4][47] , 
        \array_mux_out[4][46] , \array_mux_out[4][45] , \array_mux_out[4][44] , 
        \array_mux_out[4][43] , \array_mux_out[4][42] , \array_mux_out[4][41] , 
        \array_mux_out[4][40] , \array_mux_out[4][39] , \array_mux_out[4][38] , 
        \array_mux_out[4][37] , \array_mux_out[4][36] , \array_mux_out[4][35] , 
        \array_mux_out[4][34] , \array_mux_out[4][33] , \array_mux_out[4][32] , 
        \array_mux_out[4][31] , \array_mux_out[4][30] , \array_mux_out[4][29] , 
        \array_mux_out[4][28] , \array_mux_out[4][27] , \array_mux_out[4][26] , 
        \array_mux_out[4][25] , \array_mux_out[4][24] , \array_mux_out[4][23] , 
        \array_mux_out[4][22] , \array_mux_out[4][21] , \array_mux_out[4][20] , 
        \array_mux_out[4][19] , \array_mux_out[4][18] , \array_mux_out[4][17] , 
        \array_mux_out[4][16] , \array_mux_out[4][15] , \array_mux_out[4][14] , 
        \array_mux_out[4][13] , \array_mux_out[4][12] , \array_mux_out[4][11] , 
        \array_mux_out[4][10] , \array_mux_out[4][9] , \array_mux_out[4][8] , 
        \array_mux_out[4][7] , \array_mux_out[4][6] , \array_mux_out[4][5] , 
        \array_mux_out[4][4] , \array_mux_out[4][3] , \array_mux_out[4][2] , 
        \array_mux_out[4][1] , \array_mux_out[4][0] }), .B({
        \result_array[3][63] , \result_array[3][62] , \result_array[3][61] , 
        \result_array[3][60] , \result_array[3][59] , \result_array[3][58] , 
        \result_array[3][57] , \result_array[3][56] , \result_array[3][55] , 
        \result_array[3][54] , \result_array[3][53] , \result_array[3][52] , 
        \result_array[3][51] , \result_array[3][50] , \result_array[3][49] , 
        \result_array[3][48] , \result_array[3][47] , \result_array[3][46] , 
        \result_array[3][45] , \result_array[3][44] , \result_array[3][43] , 
        \result_array[3][42] , \result_array[3][41] , \result_array[3][40] , 
        \result_array[3][39] , \result_array[3][38] , \result_array[3][37] , 
        \result_array[3][36] , \result_array[3][35] , \result_array[3][34] , 
        \result_array[3][33] , \result_array[3][32] , \result_array[3][31] , 
        \result_array[3][30] , \result_array[3][29] , \result_array[3][28] , 
        \result_array[3][27] , \result_array[3][26] , \result_array[3][25] , 
        \result_array[3][24] , \result_array[3][23] , \result_array[3][22] , 
        \result_array[3][21] , \result_array[3][20] , \result_array[3][19] , 
        \result_array[3][18] , \result_array[3][17] , \result_array[3][16] , 
        \result_array[3][15] , \result_array[3][14] , \result_array[3][13] , 
        \result_array[3][12] , \result_array[3][11] , \result_array[3][10] , 
        \result_array[3][9] , \result_array[3][8] , \result_array[3][7] , 
        \result_array[3][6] , \result_array[3][5] , \result_array[3][4] , 
        \result_array[3][3] , \result_array[3][2] , \result_array[3][1] , 
        \result_array[3][0] }), .Cin(1'b0), .S({\result_array[4][63] , 
        \result_array[4][62] , \result_array[4][61] , \result_array[4][60] , 
        \result_array[4][59] , \result_array[4][58] , \result_array[4][57] , 
        \result_array[4][56] , \result_array[4][55] , \result_array[4][54] , 
        \result_array[4][53] , \result_array[4][52] , \result_array[4][51] , 
        \result_array[4][50] , \result_array[4][49] , \result_array[4][48] , 
        \result_array[4][47] , \result_array[4][46] , \result_array[4][45] , 
        \result_array[4][44] , \result_array[4][43] , \result_array[4][42] , 
        \result_array[4][41] , \result_array[4][40] , \result_array[4][39] , 
        \result_array[4][38] , \result_array[4][37] , \result_array[4][36] , 
        \result_array[4][35] , \result_array[4][34] , \result_array[4][33] , 
        \result_array[4][32] , \result_array[4][31] , \result_array[4][30] , 
        \result_array[4][29] , \result_array[4][28] , \result_array[4][27] , 
        \result_array[4][26] , \result_array[4][25] , \result_array[4][24] , 
        \result_array[4][23] , \result_array[4][22] , \result_array[4][21] , 
        \result_array[4][20] , \result_array[4][19] , \result_array[4][18] , 
        \result_array[4][17] , \result_array[4][16] , \result_array[4][15] , 
        \result_array[4][14] , \result_array[4][13] , \result_array[4][12] , 
        \result_array[4][11] , \result_array[4][10] , \result_array[4][9] , 
        \result_array[4][8] , \result_array[4][7] , \result_array[4][6] , 
        \result_array[4][5] , \result_array[4][4] , \result_array[4][3] , 
        \result_array[4][2] , \result_array[4][1] , \result_array[4][0] }) );
  Booth_Encoder_11 booth_j_5 ( .i(B[11:9]), .o({\select_array[5][2] , 
        \select_array[5][1] , \select_array[5][0] }) );
  MUX_booth_N64_11 mux_j_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n317, n317, 
        n318, n318, n318, n318, n318, n318, n318, n318, n318, n318, n318, n318, 
        n318, n319, n319, n319, n319, n319, n319, n319, n319, n278, n276, n273, 
        n271, n268, n266, n263, n261, n258, n256, n253, n251, n248, n246, n243, 
        n241, n238, n237, n235, n234, n71, n229, n228, n227, n224, n223, n87, 
        n220, n96, n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n170, n170, n170, n170, n170, n170, n170, n170, n169, 
        n169, n169, n169, n169, n169, n169, n169, n169, n169, n169, n169, n168, 
        n168, n159, n157, n156, n152, n150, n149, n146, n144, n142, n140, n70, 
        n68, n135, n133, n131, n130, n126, n124, n123, n92, n93, n118, n91, 
        n115, n113, n111, n110, n108, n105, n102, n99, n212, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n283, n283, n283, n283, 
        n283, n284, n284, n284, n284, n284, n284, n284, n284, n284, n284, n284, 
        n284, n285, n285, n285, n285, n285, n277, n274, n272, n269, n267, n264, 
        n262, n259, n257, n254, n252, n249, n247, n244, n242, n239, n238, n236, 
        n235, n232, n231, n230, n228, n225, A[6], n221, n85, n218, n96, n216, 
        n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n199, n199, n199, n199, n199, n199, n199, n199, n199, n198, n198, n198, 
        n198, n198, n198, n198, n198, n198, n198, n198, n198, n160, n157, n156, 
        n152, n94, n149, n147, n145, n142, n140, n138, n69, n135, n133, n132, 
        n130, n127, n124, n122, n120, n119, n117, n116, n114, n113, n111, n110, 
        n109, n106, n103, n100, n213, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[5][2] , 
        \select_array[5][1] , \select_array[5][0] }), .Y({
        \array_mux_out[5][63] , \array_mux_out[5][62] , \array_mux_out[5][61] , 
        \array_mux_out[5][60] , \array_mux_out[5][59] , \array_mux_out[5][58] , 
        \array_mux_out[5][57] , \array_mux_out[5][56] , \array_mux_out[5][55] , 
        \array_mux_out[5][54] , \array_mux_out[5][53] , \array_mux_out[5][52] , 
        \array_mux_out[5][51] , \array_mux_out[5][50] , \array_mux_out[5][49] , 
        \array_mux_out[5][48] , \array_mux_out[5][47] , \array_mux_out[5][46] , 
        \array_mux_out[5][45] , \array_mux_out[5][44] , \array_mux_out[5][43] , 
        \array_mux_out[5][42] , \array_mux_out[5][41] , \array_mux_out[5][40] , 
        \array_mux_out[5][39] , \array_mux_out[5][38] , \array_mux_out[5][37] , 
        \array_mux_out[5][36] , \array_mux_out[5][35] , \array_mux_out[5][34] , 
        \array_mux_out[5][33] , \array_mux_out[5][32] , \array_mux_out[5][31] , 
        \array_mux_out[5][30] , \array_mux_out[5][29] , \array_mux_out[5][28] , 
        \array_mux_out[5][27] , \array_mux_out[5][26] , \array_mux_out[5][25] , 
        \array_mux_out[5][24] , \array_mux_out[5][23] , \array_mux_out[5][22] , 
        \array_mux_out[5][21] , \array_mux_out[5][20] , \array_mux_out[5][19] , 
        \array_mux_out[5][18] , \array_mux_out[5][17] , \array_mux_out[5][16] , 
        \array_mux_out[5][15] , \array_mux_out[5][14] , \array_mux_out[5][13] , 
        \array_mux_out[5][12] , \array_mux_out[5][11] , \array_mux_out[5][10] , 
        \array_mux_out[5][9] , \array_mux_out[5][8] , \array_mux_out[5][7] , 
        \array_mux_out[5][6] , \array_mux_out[5][5] , \array_mux_out[5][4] , 
        \array_mux_out[5][3] , \array_mux_out[5][2] , \array_mux_out[5][1] , 
        \array_mux_out[5][0] }) );
  P4_ADDER_N64_11 adder_5 ( .A({\array_mux_out[5][63] , \array_mux_out[5][62] , 
        \array_mux_out[5][61] , \array_mux_out[5][60] , \array_mux_out[5][59] , 
        \array_mux_out[5][58] , \array_mux_out[5][57] , \array_mux_out[5][56] , 
        \array_mux_out[5][55] , \array_mux_out[5][54] , \array_mux_out[5][53] , 
        \array_mux_out[5][52] , \array_mux_out[5][51] , \array_mux_out[5][50] , 
        \array_mux_out[5][49] , \array_mux_out[5][48] , \array_mux_out[5][47] , 
        \array_mux_out[5][46] , \array_mux_out[5][45] , \array_mux_out[5][44] , 
        \array_mux_out[5][43] , \array_mux_out[5][42] , \array_mux_out[5][41] , 
        \array_mux_out[5][40] , \array_mux_out[5][39] , \array_mux_out[5][38] , 
        \array_mux_out[5][37] , \array_mux_out[5][36] , \array_mux_out[5][35] , 
        \array_mux_out[5][34] , \array_mux_out[5][33] , \array_mux_out[5][32] , 
        \array_mux_out[5][31] , \array_mux_out[5][30] , \array_mux_out[5][29] , 
        \array_mux_out[5][28] , \array_mux_out[5][27] , \array_mux_out[5][26] , 
        \array_mux_out[5][25] , \array_mux_out[5][24] , \array_mux_out[5][23] , 
        \array_mux_out[5][22] , \array_mux_out[5][21] , \array_mux_out[5][20] , 
        \array_mux_out[5][19] , \array_mux_out[5][18] , \array_mux_out[5][17] , 
        \array_mux_out[5][16] , \array_mux_out[5][15] , \array_mux_out[5][14] , 
        \array_mux_out[5][13] , \array_mux_out[5][12] , \array_mux_out[5][11] , 
        \array_mux_out[5][10] , \array_mux_out[5][9] , \array_mux_out[5][8] , 
        \array_mux_out[5][7] , \array_mux_out[5][6] , \array_mux_out[5][5] , 
        \array_mux_out[5][4] , \array_mux_out[5][3] , \array_mux_out[5][2] , 
        \array_mux_out[5][1] , \array_mux_out[5][0] }), .B({
        \result_array[4][63] , \result_array[4][62] , \result_array[4][61] , 
        \result_array[4][60] , \result_array[4][59] , \result_array[4][58] , 
        \result_array[4][57] , \result_array[4][56] , \result_array[4][55] , 
        \result_array[4][54] , \result_array[4][53] , \result_array[4][52] , 
        \result_array[4][51] , \result_array[4][50] , \result_array[4][49] , 
        \result_array[4][48] , \result_array[4][47] , \result_array[4][46] , 
        \result_array[4][45] , \result_array[4][44] , \result_array[4][43] , 
        \result_array[4][42] , \result_array[4][41] , \result_array[4][40] , 
        \result_array[4][39] , \result_array[4][38] , \result_array[4][37] , 
        \result_array[4][36] , \result_array[4][35] , \result_array[4][34] , 
        \result_array[4][33] , \result_array[4][32] , \result_array[4][31] , 
        \result_array[4][30] , \result_array[4][29] , \result_array[4][28] , 
        \result_array[4][27] , \result_array[4][26] , \result_array[4][25] , 
        \result_array[4][24] , \result_array[4][23] , \result_array[4][22] , 
        \result_array[4][21] , \result_array[4][20] , \result_array[4][19] , 
        \result_array[4][18] , \result_array[4][17] , \result_array[4][16] , 
        \result_array[4][15] , \result_array[4][14] , \result_array[4][13] , 
        \result_array[4][12] , \result_array[4][11] , \result_array[4][10] , 
        \result_array[4][9] , \result_array[4][8] , \result_array[4][7] , 
        \result_array[4][6] , \result_array[4][5] , \result_array[4][4] , 
        \result_array[4][3] , \result_array[4][2] , \result_array[4][1] , 
        \result_array[4][0] }), .Cin(1'b0), .S({\result_array[5][63] , 
        \result_array[5][62] , \result_array[5][61] , \result_array[5][60] , 
        \result_array[5][59] , \result_array[5][58] , \result_array[5][57] , 
        \result_array[5][56] , \result_array[5][55] , \result_array[5][54] , 
        \result_array[5][53] , \result_array[5][52] , \result_array[5][51] , 
        \result_array[5][50] , \result_array[5][49] , \result_array[5][48] , 
        \result_array[5][47] , \result_array[5][46] , \result_array[5][45] , 
        \result_array[5][44] , \result_array[5][43] , \result_array[5][42] , 
        \result_array[5][41] , \result_array[5][40] , \result_array[5][39] , 
        \result_array[5][38] , \result_array[5][37] , \result_array[5][36] , 
        \result_array[5][35] , \result_array[5][34] , \result_array[5][33] , 
        \result_array[5][32] , \result_array[5][31] , \result_array[5][30] , 
        \result_array[5][29] , \result_array[5][28] , \result_array[5][27] , 
        \result_array[5][26] , \result_array[5][25] , \result_array[5][24] , 
        \result_array[5][23] , \result_array[5][22] , \result_array[5][21] , 
        \result_array[5][20] , \result_array[5][19] , \result_array[5][18] , 
        \result_array[5][17] , \result_array[5][16] , \result_array[5][15] , 
        \result_array[5][14] , \result_array[5][13] , \result_array[5][12] , 
        \result_array[5][11] , \result_array[5][10] , \result_array[5][9] , 
        \result_array[5][8] , \result_array[5][7] , \result_array[5][6] , 
        \result_array[5][5] , \result_array[5][4] , \result_array[5][3] , 
        \result_array[5][2] , \result_array[5][1] , \result_array[5][0] }) );
  Booth_Encoder_10 booth_j_6 ( .i(B[13:11]), .o({\select_array[6][2] , 
        \select_array[6][1] , \select_array[6][0] }) );
  MUX_booth_N64_10 mux_j_6 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n315, n315, 
        n315, n315, n315, n315, n315, n315, n315, n315, n315, n316, n316, n316, 
        n316, n316, n316, n316, n316, n316, n316, n278, n276, n273, n271, n268, 
        n266, n263, n261, n258, n256, n253, n251, n248, n246, n243, n241, n238, 
        n237, n235, n234, n71, n229, n228, n227, n224, n223, n88, n220, n96, 
        n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n173, n173, n172, n173, n172, n173, n173, n173, n173, 
        n173, n173, n173, n173, n171, n171, n171, n171, n171, n171, n171, n159, 
        n158, n155, n153, n150, n149, n146, n145, n142, n139, n70, n68, n135, 
        n133, n131, n129, n126, n124, n122, n92, n93, n118, n91, n114, n113, 
        n111, n110, n108, n105, n102, n99, n212, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n281, n282, n282, n282, 
        n282, n282, n282, n282, n282, n282, n282, n282, n282, n283, n283, n283, 
        n283, n283, n283, n283, n277, n274, n272, n269, n267, n264, n262, n259, 
        n257, n254, n252, n249, n247, n244, n242, n239, n238, n236, n235, n232, 
        n71, n230, n228, n225, A[6], n221, n89, n218, n96, n216, n97, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n201, n201, n201, n201, n200, n200, n200, n200, n200, n200, n200, n200, 
        n200, n200, n200, n200, n199, n199, n199, n160, n157, n155, n153, n150, 
        n149, n147, n145, n142, n140, n70, n69, n135, n133, n132, n130, n127, 
        n124, n122, n120, n119, n117, n116, n114, n113, n111, n110, n109, n106, 
        n103, n100, n213, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[6][2] , 
        \select_array[6][1] , \select_array[6][0] }), .Y({
        \array_mux_out[6][63] , \array_mux_out[6][62] , \array_mux_out[6][61] , 
        \array_mux_out[6][60] , \array_mux_out[6][59] , \array_mux_out[6][58] , 
        \array_mux_out[6][57] , \array_mux_out[6][56] , \array_mux_out[6][55] , 
        \array_mux_out[6][54] , \array_mux_out[6][53] , \array_mux_out[6][52] , 
        \array_mux_out[6][51] , \array_mux_out[6][50] , \array_mux_out[6][49] , 
        \array_mux_out[6][48] , \array_mux_out[6][47] , \array_mux_out[6][46] , 
        \array_mux_out[6][45] , \array_mux_out[6][44] , \array_mux_out[6][43] , 
        \array_mux_out[6][42] , \array_mux_out[6][41] , \array_mux_out[6][40] , 
        \array_mux_out[6][39] , \array_mux_out[6][38] , \array_mux_out[6][37] , 
        \array_mux_out[6][36] , \array_mux_out[6][35] , \array_mux_out[6][34] , 
        \array_mux_out[6][33] , \array_mux_out[6][32] , \array_mux_out[6][31] , 
        \array_mux_out[6][30] , \array_mux_out[6][29] , \array_mux_out[6][28] , 
        \array_mux_out[6][27] , \array_mux_out[6][26] , \array_mux_out[6][25] , 
        \array_mux_out[6][24] , \array_mux_out[6][23] , \array_mux_out[6][22] , 
        \array_mux_out[6][21] , \array_mux_out[6][20] , \array_mux_out[6][19] , 
        \array_mux_out[6][18] , \array_mux_out[6][17] , \array_mux_out[6][16] , 
        \array_mux_out[6][15] , \array_mux_out[6][14] , \array_mux_out[6][13] , 
        \array_mux_out[6][12] , \array_mux_out[6][11] , \array_mux_out[6][10] , 
        \array_mux_out[6][9] , \array_mux_out[6][8] , \array_mux_out[6][7] , 
        \array_mux_out[6][6] , \array_mux_out[6][5] , \array_mux_out[6][4] , 
        \array_mux_out[6][3] , \array_mux_out[6][2] , \array_mux_out[6][1] , 
        \array_mux_out[6][0] }) );
  P4_ADDER_N64_10 adder_6 ( .A({\array_mux_out[6][63] , \array_mux_out[6][62] , 
        \array_mux_out[6][61] , \array_mux_out[6][60] , \array_mux_out[6][59] , 
        \array_mux_out[6][58] , \array_mux_out[6][57] , \array_mux_out[6][56] , 
        \array_mux_out[6][55] , \array_mux_out[6][54] , \array_mux_out[6][53] , 
        \array_mux_out[6][52] , \array_mux_out[6][51] , \array_mux_out[6][50] , 
        \array_mux_out[6][49] , \array_mux_out[6][48] , \array_mux_out[6][47] , 
        \array_mux_out[6][46] , \array_mux_out[6][45] , \array_mux_out[6][44] , 
        \array_mux_out[6][43] , \array_mux_out[6][42] , \array_mux_out[6][41] , 
        \array_mux_out[6][40] , \array_mux_out[6][39] , \array_mux_out[6][38] , 
        \array_mux_out[6][37] , \array_mux_out[6][36] , \array_mux_out[6][35] , 
        \array_mux_out[6][34] , \array_mux_out[6][33] , \array_mux_out[6][32] , 
        \array_mux_out[6][31] , \array_mux_out[6][30] , \array_mux_out[6][29] , 
        \array_mux_out[6][28] , \array_mux_out[6][27] , \array_mux_out[6][26] , 
        \array_mux_out[6][25] , \array_mux_out[6][24] , \array_mux_out[6][23] , 
        \array_mux_out[6][22] , \array_mux_out[6][21] , \array_mux_out[6][20] , 
        \array_mux_out[6][19] , \array_mux_out[6][18] , \array_mux_out[6][17] , 
        \array_mux_out[6][16] , \array_mux_out[6][15] , \array_mux_out[6][14] , 
        \array_mux_out[6][13] , \array_mux_out[6][12] , \array_mux_out[6][11] , 
        \array_mux_out[6][10] , \array_mux_out[6][9] , \array_mux_out[6][8] , 
        \array_mux_out[6][7] , \array_mux_out[6][6] , \array_mux_out[6][5] , 
        \array_mux_out[6][4] , \array_mux_out[6][3] , \array_mux_out[6][2] , 
        \array_mux_out[6][1] , \array_mux_out[6][0] }), .B({
        \result_array[5][63] , \result_array[5][62] , \result_array[5][61] , 
        \result_array[5][60] , \result_array[5][59] , \result_array[5][58] , 
        \result_array[5][57] , \result_array[5][56] , \result_array[5][55] , 
        \result_array[5][54] , \result_array[5][53] , \result_array[5][52] , 
        \result_array[5][51] , \result_array[5][50] , \result_array[5][49] , 
        \result_array[5][48] , \result_array[5][47] , \result_array[5][46] , 
        \result_array[5][45] , \result_array[5][44] , \result_array[5][43] , 
        \result_array[5][42] , \result_array[5][41] , \result_array[5][40] , 
        \result_array[5][39] , \result_array[5][38] , \result_array[5][37] , 
        \result_array[5][36] , \result_array[5][35] , \result_array[5][34] , 
        \result_array[5][33] , \result_array[5][32] , \result_array[5][31] , 
        \result_array[5][30] , \result_array[5][29] , \result_array[5][28] , 
        \result_array[5][27] , \result_array[5][26] , \result_array[5][25] , 
        \result_array[5][24] , \result_array[5][23] , \result_array[5][22] , 
        \result_array[5][21] , \result_array[5][20] , \result_array[5][19] , 
        \result_array[5][18] , \result_array[5][17] , \result_array[5][16] , 
        \result_array[5][15] , \result_array[5][14] , \result_array[5][13] , 
        \result_array[5][12] , \result_array[5][11] , \result_array[5][10] , 
        \result_array[5][9] , \result_array[5][8] , \result_array[5][7] , 
        \result_array[5][6] , \result_array[5][5] , \result_array[5][4] , 
        \result_array[5][3] , \result_array[5][2] , \result_array[5][1] , 
        \result_array[5][0] }), .Cin(1'b0), .S({\result_array[6][63] , 
        \result_array[6][62] , \result_array[6][61] , \result_array[6][60] , 
        \result_array[6][59] , \result_array[6][58] , \result_array[6][57] , 
        \result_array[6][56] , \result_array[6][55] , \result_array[6][54] , 
        \result_array[6][53] , \result_array[6][52] , \result_array[6][51] , 
        \result_array[6][50] , \result_array[6][49] , \result_array[6][48] , 
        \result_array[6][47] , \result_array[6][46] , \result_array[6][45] , 
        \result_array[6][44] , \result_array[6][43] , \result_array[6][42] , 
        \result_array[6][41] , \result_array[6][40] , \result_array[6][39] , 
        \result_array[6][38] , \result_array[6][37] , \result_array[6][36] , 
        \result_array[6][35] , \result_array[6][34] , \result_array[6][33] , 
        \result_array[6][32] , \result_array[6][31] , \result_array[6][30] , 
        \result_array[6][29] , \result_array[6][28] , \result_array[6][27] , 
        \result_array[6][26] , \result_array[6][25] , \result_array[6][24] , 
        \result_array[6][23] , \result_array[6][22] , \result_array[6][21] , 
        \result_array[6][20] , \result_array[6][19] , \result_array[6][18] , 
        \result_array[6][17] , \result_array[6][16] , \result_array[6][15] , 
        \result_array[6][14] , \result_array[6][13] , \result_array[6][12] , 
        \result_array[6][11] , \result_array[6][10] , \result_array[6][9] , 
        \result_array[6][8] , \result_array[6][7] , \result_array[6][6] , 
        \result_array[6][5] , \result_array[6][4] , \result_array[6][3] , 
        \result_array[6][2] , \result_array[6][1] , \result_array[6][0] }) );
  Booth_Encoder_9 booth_j_7 ( .i(B[15:13]), .o({\select_array[7][2] , 
        \select_array[7][1] , \select_array[7][0] }) );
  MUX_booth_N64_9 mux_j_7 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n312, n312, n313, 
        n313, n313, n313, n313, n313, n313, n313, n313, n313, n313, n313, n313, 
        n314, n314, n314, n314, n278, n275, n272, n271, n268, n265, n262, n261, 
        n258, n255, n252, n251, n248, n245, n242, n241, n238, n236, n235, n234, 
        n72, n230, n228, n227, n224, n222, n90, n220, n96, n216, n97, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .C({n172, n172, n172, n172, n172, n173, n172, n173, n172, n173, 
        n173, n173, n173, n173, n173, n173, n173, n173, n159, n157, n156, n152, 
        n150, n149, n146, n144, n142, n140, n138, n68, n135, n133, n131, n129, 
        n126, n124, n123, n92, n93, n118, n91, n114, n113, n111, n110, n108, 
        n105, n102, n99, n212, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n280, n280, n280, n280, n280, 
        n280, n280, n281, n281, n281, n281, n281, n281, n281, n281, n281, n281, 
        n281, n277, n274, n272, n269, n267, n264, n262, n259, n257, n254, n252, 
        n249, n247, n244, n242, n239, n238, n236, n235, n232, n72, n229, n228, 
        n225, A[6], n221, n90, n218, n96, n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .E({n202, n202, n202, n202, n202, n202, n202, n202, n202, n201, n201, 
        n201, n201, n201, n201, n201, n201, n160, n158, n155, n153, n150, n149, 
        n147, n145, n142, n139, n70, n68, n135, n133, n132, n130, n127, n124, 
        n123, n120, n119, n117, n116, n115, n113, n111, n110, n109, n106, n103, 
        n100, n213, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[7][2] , 
        \select_array[7][1] , \select_array[7][0] }), .Y({
        \array_mux_out[7][63] , \array_mux_out[7][62] , \array_mux_out[7][61] , 
        \array_mux_out[7][60] , \array_mux_out[7][59] , \array_mux_out[7][58] , 
        \array_mux_out[7][57] , \array_mux_out[7][56] , \array_mux_out[7][55] , 
        \array_mux_out[7][54] , \array_mux_out[7][53] , \array_mux_out[7][52] , 
        \array_mux_out[7][51] , \array_mux_out[7][50] , \array_mux_out[7][49] , 
        \array_mux_out[7][48] , \array_mux_out[7][47] , \array_mux_out[7][46] , 
        \array_mux_out[7][45] , \array_mux_out[7][44] , \array_mux_out[7][43] , 
        \array_mux_out[7][42] , \array_mux_out[7][41] , \array_mux_out[7][40] , 
        \array_mux_out[7][39] , \array_mux_out[7][38] , \array_mux_out[7][37] , 
        \array_mux_out[7][36] , \array_mux_out[7][35] , \array_mux_out[7][34] , 
        \array_mux_out[7][33] , \array_mux_out[7][32] , \array_mux_out[7][31] , 
        \array_mux_out[7][30] , \array_mux_out[7][29] , \array_mux_out[7][28] , 
        \array_mux_out[7][27] , \array_mux_out[7][26] , \array_mux_out[7][25] , 
        \array_mux_out[7][24] , \array_mux_out[7][23] , \array_mux_out[7][22] , 
        \array_mux_out[7][21] , \array_mux_out[7][20] , \array_mux_out[7][19] , 
        \array_mux_out[7][18] , \array_mux_out[7][17] , \array_mux_out[7][16] , 
        \array_mux_out[7][15] , \array_mux_out[7][14] , \array_mux_out[7][13] , 
        \array_mux_out[7][12] , \array_mux_out[7][11] , \array_mux_out[7][10] , 
        \array_mux_out[7][9] , \array_mux_out[7][8] , \array_mux_out[7][7] , 
        \array_mux_out[7][6] , \array_mux_out[7][5] , \array_mux_out[7][4] , 
        \array_mux_out[7][3] , \array_mux_out[7][2] , \array_mux_out[7][1] , 
        \array_mux_out[7][0] }) );
  P4_ADDER_N64_9 adder_7 ( .A({\array_mux_out[7][63] , \array_mux_out[7][62] , 
        \array_mux_out[7][61] , \array_mux_out[7][60] , \array_mux_out[7][59] , 
        \array_mux_out[7][58] , \array_mux_out[7][57] , \array_mux_out[7][56] , 
        \array_mux_out[7][55] , \array_mux_out[7][54] , \array_mux_out[7][53] , 
        \array_mux_out[7][52] , \array_mux_out[7][51] , \array_mux_out[7][50] , 
        \array_mux_out[7][49] , \array_mux_out[7][48] , \array_mux_out[7][47] , 
        \array_mux_out[7][46] , \array_mux_out[7][45] , \array_mux_out[7][44] , 
        \array_mux_out[7][43] , \array_mux_out[7][42] , \array_mux_out[7][41] , 
        \array_mux_out[7][40] , \array_mux_out[7][39] , \array_mux_out[7][38] , 
        \array_mux_out[7][37] , \array_mux_out[7][36] , \array_mux_out[7][35] , 
        \array_mux_out[7][34] , \array_mux_out[7][33] , \array_mux_out[7][32] , 
        \array_mux_out[7][31] , \array_mux_out[7][30] , \array_mux_out[7][29] , 
        \array_mux_out[7][28] , \array_mux_out[7][27] , \array_mux_out[7][26] , 
        \array_mux_out[7][25] , \array_mux_out[7][24] , \array_mux_out[7][23] , 
        \array_mux_out[7][22] , \array_mux_out[7][21] , \array_mux_out[7][20] , 
        \array_mux_out[7][19] , \array_mux_out[7][18] , \array_mux_out[7][17] , 
        \array_mux_out[7][16] , \array_mux_out[7][15] , \array_mux_out[7][14] , 
        \array_mux_out[7][13] , \array_mux_out[7][12] , \array_mux_out[7][11] , 
        \array_mux_out[7][10] , \array_mux_out[7][9] , \array_mux_out[7][8] , 
        \array_mux_out[7][7] , \array_mux_out[7][6] , \array_mux_out[7][5] , 
        \array_mux_out[7][4] , \array_mux_out[7][3] , \array_mux_out[7][2] , 
        \array_mux_out[7][1] , \array_mux_out[7][0] }), .B({
        \result_array[6][63] , \result_array[6][62] , \result_array[6][61] , 
        \result_array[6][60] , \result_array[6][59] , \result_array[6][58] , 
        \result_array[6][57] , \result_array[6][56] , \result_array[6][55] , 
        \result_array[6][54] , \result_array[6][53] , \result_array[6][52] , 
        \result_array[6][51] , \result_array[6][50] , \result_array[6][49] , 
        \result_array[6][48] , \result_array[6][47] , \result_array[6][46] , 
        \result_array[6][45] , \result_array[6][44] , \result_array[6][43] , 
        \result_array[6][42] , \result_array[6][41] , \result_array[6][40] , 
        \result_array[6][39] , \result_array[6][38] , \result_array[6][37] , 
        \result_array[6][36] , \result_array[6][35] , \result_array[6][34] , 
        \result_array[6][33] , \result_array[6][32] , \result_array[6][31] , 
        \result_array[6][30] , \result_array[6][29] , \result_array[6][28] , 
        \result_array[6][27] , \result_array[6][26] , \result_array[6][25] , 
        \result_array[6][24] , \result_array[6][23] , \result_array[6][22] , 
        \result_array[6][21] , \result_array[6][20] , \result_array[6][19] , 
        \result_array[6][18] , \result_array[6][17] , \result_array[6][16] , 
        \result_array[6][15] , \result_array[6][14] , \result_array[6][13] , 
        \result_array[6][12] , \result_array[6][11] , \result_array[6][10] , 
        \result_array[6][9] , \result_array[6][8] , \result_array[6][7] , 
        \result_array[6][6] , \result_array[6][5] , \result_array[6][4] , 
        \result_array[6][3] , \result_array[6][2] , \result_array[6][1] , 
        \result_array[6][0] }), .Cin(1'b0), .S({\result_array[7][63] , 
        \result_array[7][62] , \result_array[7][61] , \result_array[7][60] , 
        \result_array[7][59] , \result_array[7][58] , \result_array[7][57] , 
        \result_array[7][56] , \result_array[7][55] , \result_array[7][54] , 
        \result_array[7][53] , \result_array[7][52] , \result_array[7][51] , 
        \result_array[7][50] , \result_array[7][49] , \result_array[7][48] , 
        \result_array[7][47] , \result_array[7][46] , \result_array[7][45] , 
        \result_array[7][44] , \result_array[7][43] , \result_array[7][42] , 
        \result_array[7][41] , \result_array[7][40] , \result_array[7][39] , 
        \result_array[7][38] , \result_array[7][37] , \result_array[7][36] , 
        \result_array[7][35] , \result_array[7][34] , \result_array[7][33] , 
        \result_array[7][32] , \result_array[7][31] , \result_array[7][30] , 
        \result_array[7][29] , \result_array[7][28] , \result_array[7][27] , 
        \result_array[7][26] , \result_array[7][25] , \result_array[7][24] , 
        \result_array[7][23] , \result_array[7][22] , \result_array[7][21] , 
        \result_array[7][20] , \result_array[7][19] , \result_array[7][18] , 
        \result_array[7][17] , \result_array[7][16] , \result_array[7][15] , 
        \result_array[7][14] , \result_array[7][13] , \result_array[7][12] , 
        \result_array[7][11] , \result_array[7][10] , \result_array[7][9] , 
        \result_array[7][8] , \result_array[7][7] , \result_array[7][6] , 
        \result_array[7][5] , \result_array[7][4] , \result_array[7][3] , 
        \result_array[7][2] , \result_array[7][1] , \result_array[7][0] }) );
  Booth_Encoder_8 booth_j_8 ( .i(B[17:15]), .o({\select_array[8][2] , 
        \select_array[8][1] , \select_array[8][0] }) );
  MUX_booth_N64_8 mux_j_8 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n302, n317, n311, 
        n311, n311, n311, n311, n311, n311, n311, n312, n312, n312, n312, n312, 
        n312, n312, n278, n275, n272, n270, n268, n265, n262, n260, n258, n255, 
        n252, n250, n248, n245, n242, n240, n238, n236, n235, n233, n71, n229, 
        n228, n226, n224, n222, n90, n219, n96, n216, n97, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .C({n172, n172, n172, n172, n173, n173, n173, n164, n173, n173, 
        n173, n173, n173, n172, n173, n173, n159, n158, n155, n153, n94, n149, 
        n146, n145, n142, n140, n70, n68, n135, n133, n131, n130, n126, n124, 
        n123, n92, n93, n118, n91, n115, n113, n111, n110, n108, n105, n102, 
        n99, n212, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n279, n279, n279, n279, n279, 
        n279, n279, n294, n279, n279, n279, n280, n280, n280, n280, n280, n277, 
        n274, n272, n269, n267, n264, n262, n259, n257, n254, n252, n249, n247, 
        n244, n242, n239, n238, n236, n235, n232, n231, n230, n228, n225, A[6], 
        n221, n76, n218, n96, n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .E({n203, n203, n203, n203, n203, n203, n203, n203, n203, n203, n203, 
        n203, n202, n202, n202, n160, n158, n155, n153, n150, n149, n147, n144, 
        n142, n139, n70, n68, n135, n133, n132, n129, n127, n124, n123, n92, 
        n119, n118, n116, n114, n113, n111, n110, n109, n106, n103, n100, n213, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[8][2] , 
        \select_array[8][1] , \select_array[8][0] }), .Y({
        \array_mux_out[8][63] , \array_mux_out[8][62] , \array_mux_out[8][61] , 
        \array_mux_out[8][60] , \array_mux_out[8][59] , \array_mux_out[8][58] , 
        \array_mux_out[8][57] , \array_mux_out[8][56] , \array_mux_out[8][55] , 
        \array_mux_out[8][54] , \array_mux_out[8][53] , \array_mux_out[8][52] , 
        \array_mux_out[8][51] , \array_mux_out[8][50] , \array_mux_out[8][49] , 
        \array_mux_out[8][48] , \array_mux_out[8][47] , \array_mux_out[8][46] , 
        \array_mux_out[8][45] , \array_mux_out[8][44] , \array_mux_out[8][43] , 
        \array_mux_out[8][42] , \array_mux_out[8][41] , \array_mux_out[8][40] , 
        \array_mux_out[8][39] , \array_mux_out[8][38] , \array_mux_out[8][37] , 
        \array_mux_out[8][36] , \array_mux_out[8][35] , \array_mux_out[8][34] , 
        \array_mux_out[8][33] , \array_mux_out[8][32] , \array_mux_out[8][31] , 
        \array_mux_out[8][30] , \array_mux_out[8][29] , \array_mux_out[8][28] , 
        \array_mux_out[8][27] , \array_mux_out[8][26] , \array_mux_out[8][25] , 
        \array_mux_out[8][24] , \array_mux_out[8][23] , \array_mux_out[8][22] , 
        \array_mux_out[8][21] , \array_mux_out[8][20] , \array_mux_out[8][19] , 
        \array_mux_out[8][18] , \array_mux_out[8][17] , \array_mux_out[8][16] , 
        \array_mux_out[8][15] , \array_mux_out[8][14] , \array_mux_out[8][13] , 
        \array_mux_out[8][12] , \array_mux_out[8][11] , \array_mux_out[8][10] , 
        \array_mux_out[8][9] , \array_mux_out[8][8] , \array_mux_out[8][7] , 
        \array_mux_out[8][6] , \array_mux_out[8][5] , \array_mux_out[8][4] , 
        \array_mux_out[8][3] , \array_mux_out[8][2] , \array_mux_out[8][1] , 
        \array_mux_out[8][0] }) );
  P4_ADDER_N64_8 adder_8 ( .A({\array_mux_out[8][63] , \array_mux_out[8][62] , 
        \array_mux_out[8][61] , \array_mux_out[8][60] , \array_mux_out[8][59] , 
        \array_mux_out[8][58] , \array_mux_out[8][57] , \array_mux_out[8][56] , 
        \array_mux_out[8][55] , \array_mux_out[8][54] , \array_mux_out[8][53] , 
        \array_mux_out[8][52] , \array_mux_out[8][51] , \array_mux_out[8][50] , 
        \array_mux_out[8][49] , \array_mux_out[8][48] , \array_mux_out[8][47] , 
        \array_mux_out[8][46] , \array_mux_out[8][45] , \array_mux_out[8][44] , 
        \array_mux_out[8][43] , \array_mux_out[8][42] , \array_mux_out[8][41] , 
        \array_mux_out[8][40] , \array_mux_out[8][39] , \array_mux_out[8][38] , 
        \array_mux_out[8][37] , \array_mux_out[8][36] , \array_mux_out[8][35] , 
        \array_mux_out[8][34] , \array_mux_out[8][33] , \array_mux_out[8][32] , 
        \array_mux_out[8][31] , \array_mux_out[8][30] , \array_mux_out[8][29] , 
        \array_mux_out[8][28] , \array_mux_out[8][27] , \array_mux_out[8][26] , 
        \array_mux_out[8][25] , \array_mux_out[8][24] , \array_mux_out[8][23] , 
        \array_mux_out[8][22] , \array_mux_out[8][21] , \array_mux_out[8][20] , 
        \array_mux_out[8][19] , \array_mux_out[8][18] , \array_mux_out[8][17] , 
        \array_mux_out[8][16] , \array_mux_out[8][15] , \array_mux_out[8][14] , 
        \array_mux_out[8][13] , \array_mux_out[8][12] , \array_mux_out[8][11] , 
        \array_mux_out[8][10] , \array_mux_out[8][9] , \array_mux_out[8][8] , 
        \array_mux_out[8][7] , \array_mux_out[8][6] , \array_mux_out[8][5] , 
        \array_mux_out[8][4] , \array_mux_out[8][3] , \array_mux_out[8][2] , 
        \array_mux_out[8][1] , \array_mux_out[8][0] }), .B({
        \result_array[7][63] , \result_array[7][62] , \result_array[7][61] , 
        \result_array[7][60] , \result_array[7][59] , \result_array[7][58] , 
        \result_array[7][57] , \result_array[7][56] , \result_array[7][55] , 
        \result_array[7][54] , \result_array[7][53] , \result_array[7][52] , 
        \result_array[7][51] , \result_array[7][50] , \result_array[7][49] , 
        \result_array[7][48] , \result_array[7][47] , \result_array[7][46] , 
        \result_array[7][45] , \result_array[7][44] , \result_array[7][43] , 
        \result_array[7][42] , \result_array[7][41] , \result_array[7][40] , 
        \result_array[7][39] , \result_array[7][38] , \result_array[7][37] , 
        \result_array[7][36] , \result_array[7][35] , \result_array[7][34] , 
        \result_array[7][33] , \result_array[7][32] , \result_array[7][31] , 
        \result_array[7][30] , \result_array[7][29] , \result_array[7][28] , 
        \result_array[7][27] , \result_array[7][26] , \result_array[7][25] , 
        \result_array[7][24] , \result_array[7][23] , \result_array[7][22] , 
        \result_array[7][21] , \result_array[7][20] , \result_array[7][19] , 
        \result_array[7][18] , \result_array[7][17] , \result_array[7][16] , 
        \result_array[7][15] , \result_array[7][14] , \result_array[7][13] , 
        \result_array[7][12] , \result_array[7][11] , \result_array[7][10] , 
        \result_array[7][9] , \result_array[7][8] , \result_array[7][7] , 
        \result_array[7][6] , \result_array[7][5] , \result_array[7][4] , 
        \result_array[7][3] , \result_array[7][2] , \result_array[7][1] , 
        \result_array[7][0] }), .Cin(1'b0), .S({\result_array[8][63] , 
        \result_array[8][62] , \result_array[8][61] , \result_array[8][60] , 
        \result_array[8][59] , \result_array[8][58] , \result_array[8][57] , 
        \result_array[8][56] , \result_array[8][55] , \result_array[8][54] , 
        \result_array[8][53] , \result_array[8][52] , \result_array[8][51] , 
        \result_array[8][50] , \result_array[8][49] , \result_array[8][48] , 
        \result_array[8][47] , \result_array[8][46] , \result_array[8][45] , 
        \result_array[8][44] , \result_array[8][43] , \result_array[8][42] , 
        \result_array[8][41] , \result_array[8][40] , \result_array[8][39] , 
        \result_array[8][38] , \result_array[8][37] , \result_array[8][36] , 
        \result_array[8][35] , \result_array[8][34] , \result_array[8][33] , 
        \result_array[8][32] , \result_array[8][31] , \result_array[8][30] , 
        \result_array[8][29] , \result_array[8][28] , \result_array[8][27] , 
        \result_array[8][26] , \result_array[8][25] , \result_array[8][24] , 
        \result_array[8][23] , \result_array[8][22] , \result_array[8][21] , 
        \result_array[8][20] , \result_array[8][19] , \result_array[8][18] , 
        \result_array[8][17] , \result_array[8][16] , \result_array[8][15] , 
        \result_array[8][14] , \result_array[8][13] , \result_array[8][12] , 
        \result_array[8][11] , \result_array[8][10] , \result_array[8][9] , 
        \result_array[8][8] , \result_array[8][7] , \result_array[8][6] , 
        \result_array[8][5] , \result_array[8][4] , \result_array[8][3] , 
        \result_array[8][2] , \result_array[8][1] , \result_array[8][0] }) );
  Booth_Encoder_7 booth_j_9 ( .i(B[19:17]), .o({\select_array[9][2] , 
        \select_array[9][1] , \select_array[9][0] }) );
  MUX_booth_N64_7 mux_j_9 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n315, n315, n314, 
        n314, n314, n314, n314, n314, n314, n314, n314, n312, n312, n312, n312, 
        n277, n275, n272, n270, n267, n265, n262, n260, n257, n255, n252, n250, 
        n247, n245, n242, n240, n238, n236, n235, n233, n72, n230, n228, n226, 
        A[6], n222, n77, n219, n96, n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .C({n171, n171, n172, n172, n172, n172, n172, n173, n173, n173, 
        n173, n173, n173, n173, n159, n157, n155, n153, n94, n149, n146, n145, 
        n142, n139, n138, n68, n135, n133, n131, n130, n126, n124, n123, n120, 
        n93, n118, n91, n114, n113, n111, n110, n108, n105, n102, n99, n212, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n301, n301, n301, n301, n300, 
        n301, n300, n300, n300, n300, n301, n300, n301, n286, n277, n274, n272, 
        n269, n267, n264, n262, n259, n257, n254, n252, n249, n247, n244, n242, 
        n239, n238, n236, n235, n232, n231, n229, n228, n225, A[6], n221, n75, 
        n218, n96, n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .E({n183, n183, n183, n182, n183, n183, n183, n183, n182, n183, n182, 
        n183, n182, n160, n157, n155, n153, n150, n149, n147, n144, n142, n140, 
        n70, n69, n135, n133, n132, n130, n127, n124, n122, n92, n119, n117, 
        n116, n114, n113, n111, n110, n109, n106, n103, n100, n213, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[9][2] , 
        \select_array[9][1] , \select_array[9][0] }), .Y({
        \array_mux_out[9][63] , \array_mux_out[9][62] , \array_mux_out[9][61] , 
        \array_mux_out[9][60] , \array_mux_out[9][59] , \array_mux_out[9][58] , 
        \array_mux_out[9][57] , \array_mux_out[9][56] , \array_mux_out[9][55] , 
        \array_mux_out[9][54] , \array_mux_out[9][53] , \array_mux_out[9][52] , 
        \array_mux_out[9][51] , \array_mux_out[9][50] , \array_mux_out[9][49] , 
        \array_mux_out[9][48] , \array_mux_out[9][47] , \array_mux_out[9][46] , 
        \array_mux_out[9][45] , \array_mux_out[9][44] , \array_mux_out[9][43] , 
        \array_mux_out[9][42] , \array_mux_out[9][41] , \array_mux_out[9][40] , 
        \array_mux_out[9][39] , \array_mux_out[9][38] , \array_mux_out[9][37] , 
        \array_mux_out[9][36] , \array_mux_out[9][35] , \array_mux_out[9][34] , 
        \array_mux_out[9][33] , \array_mux_out[9][32] , \array_mux_out[9][31] , 
        \array_mux_out[9][30] , \array_mux_out[9][29] , \array_mux_out[9][28] , 
        \array_mux_out[9][27] , \array_mux_out[9][26] , \array_mux_out[9][25] , 
        \array_mux_out[9][24] , \array_mux_out[9][23] , \array_mux_out[9][22] , 
        \array_mux_out[9][21] , \array_mux_out[9][20] , \array_mux_out[9][19] , 
        \array_mux_out[9][18] , \array_mux_out[9][17] , \array_mux_out[9][16] , 
        \array_mux_out[9][15] , \array_mux_out[9][14] , \array_mux_out[9][13] , 
        \array_mux_out[9][12] , \array_mux_out[9][11] , \array_mux_out[9][10] , 
        \array_mux_out[9][9] , \array_mux_out[9][8] , \array_mux_out[9][7] , 
        \array_mux_out[9][6] , \array_mux_out[9][5] , \array_mux_out[9][4] , 
        \array_mux_out[9][3] , \array_mux_out[9][2] , \array_mux_out[9][1] , 
        \array_mux_out[9][0] }) );
  P4_ADDER_N64_7 adder_9 ( .A({\array_mux_out[9][63] , \array_mux_out[9][62] , 
        \array_mux_out[9][61] , \array_mux_out[9][60] , \array_mux_out[9][59] , 
        \array_mux_out[9][58] , \array_mux_out[9][57] , \array_mux_out[9][56] , 
        \array_mux_out[9][55] , \array_mux_out[9][54] , \array_mux_out[9][53] , 
        \array_mux_out[9][52] , \array_mux_out[9][51] , \array_mux_out[9][50] , 
        \array_mux_out[9][49] , \array_mux_out[9][48] , \array_mux_out[9][47] , 
        \array_mux_out[9][46] , \array_mux_out[9][45] , \array_mux_out[9][44] , 
        \array_mux_out[9][43] , \array_mux_out[9][42] , \array_mux_out[9][41] , 
        \array_mux_out[9][40] , \array_mux_out[9][39] , \array_mux_out[9][38] , 
        \array_mux_out[9][37] , \array_mux_out[9][36] , \array_mux_out[9][35] , 
        \array_mux_out[9][34] , \array_mux_out[9][33] , \array_mux_out[9][32] , 
        \array_mux_out[9][31] , \array_mux_out[9][30] , \array_mux_out[9][29] , 
        \array_mux_out[9][28] , \array_mux_out[9][27] , \array_mux_out[9][26] , 
        \array_mux_out[9][25] , \array_mux_out[9][24] , \array_mux_out[9][23] , 
        \array_mux_out[9][22] , \array_mux_out[9][21] , \array_mux_out[9][20] , 
        \array_mux_out[9][19] , \array_mux_out[9][18] , \array_mux_out[9][17] , 
        \array_mux_out[9][16] , \array_mux_out[9][15] , \array_mux_out[9][14] , 
        \array_mux_out[9][13] , \array_mux_out[9][12] , \array_mux_out[9][11] , 
        \array_mux_out[9][10] , \array_mux_out[9][9] , \array_mux_out[9][8] , 
        \array_mux_out[9][7] , \array_mux_out[9][6] , \array_mux_out[9][5] , 
        \array_mux_out[9][4] , \array_mux_out[9][3] , \array_mux_out[9][2] , 
        \array_mux_out[9][1] , \array_mux_out[9][0] }), .B({
        \result_array[8][63] , \result_array[8][62] , \result_array[8][61] , 
        \result_array[8][60] , \result_array[8][59] , \result_array[8][58] , 
        \result_array[8][57] , \result_array[8][56] , \result_array[8][55] , 
        \result_array[8][54] , \result_array[8][53] , \result_array[8][52] , 
        \result_array[8][51] , \result_array[8][50] , \result_array[8][49] , 
        \result_array[8][48] , \result_array[8][47] , \result_array[8][46] , 
        \result_array[8][45] , \result_array[8][44] , \result_array[8][43] , 
        \result_array[8][42] , \result_array[8][41] , \result_array[8][40] , 
        \result_array[8][39] , \result_array[8][38] , \result_array[8][37] , 
        \result_array[8][36] , \result_array[8][35] , \result_array[8][34] , 
        \result_array[8][33] , \result_array[8][32] , \result_array[8][31] , 
        \result_array[8][30] , \result_array[8][29] , \result_array[8][28] , 
        \result_array[8][27] , \result_array[8][26] , \result_array[8][25] , 
        \result_array[8][24] , \result_array[8][23] , \result_array[8][22] , 
        \result_array[8][21] , \result_array[8][20] , \result_array[8][19] , 
        \result_array[8][18] , \result_array[8][17] , \result_array[8][16] , 
        \result_array[8][15] , \result_array[8][14] , \result_array[8][13] , 
        \result_array[8][12] , \result_array[8][11] , \result_array[8][10] , 
        \result_array[8][9] , \result_array[8][8] , \result_array[8][7] , 
        \result_array[8][6] , \result_array[8][5] , \result_array[8][4] , 
        \result_array[8][3] , \result_array[8][2] , \result_array[8][1] , 
        \result_array[8][0] }), .Cin(1'b0), .S({\result_array[9][63] , 
        \result_array[9][62] , \result_array[9][61] , \result_array[9][60] , 
        \result_array[9][59] , \result_array[9][58] , \result_array[9][57] , 
        \result_array[9][56] , \result_array[9][55] , \result_array[9][54] , 
        \result_array[9][53] , \result_array[9][52] , \result_array[9][51] , 
        \result_array[9][50] , \result_array[9][49] , \result_array[9][48] , 
        \result_array[9][47] , \result_array[9][46] , \result_array[9][45] , 
        \result_array[9][44] , \result_array[9][43] , \result_array[9][42] , 
        \result_array[9][41] , \result_array[9][40] , \result_array[9][39] , 
        \result_array[9][38] , \result_array[9][37] , \result_array[9][36] , 
        \result_array[9][35] , \result_array[9][34] , \result_array[9][33] , 
        \result_array[9][32] , \result_array[9][31] , \result_array[9][30] , 
        \result_array[9][29] , \result_array[9][28] , \result_array[9][27] , 
        \result_array[9][26] , \result_array[9][25] , \result_array[9][24] , 
        \result_array[9][23] , \result_array[9][22] , \result_array[9][21] , 
        \result_array[9][20] , \result_array[9][19] , \result_array[9][18] , 
        \result_array[9][17] , \result_array[9][16] , \result_array[9][15] , 
        \result_array[9][14] , \result_array[9][13] , \result_array[9][12] , 
        \result_array[9][11] , \result_array[9][10] , \result_array[9][9] , 
        \result_array[9][8] , \result_array[9][7] , \result_array[9][6] , 
        \result_array[9][5] , \result_array[9][4] , \result_array[9][3] , 
        \result_array[9][2] , \result_array[9][1] , \result_array[9][0] }) );
  Booth_Encoder_6 booth_j_10 ( .i(B[21:19]), .o({\select_array[10][2] , 
        \select_array[10][1] , \select_array[10][0] }) );
  MUX_booth_N64_6 mux_j_10 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n317, n317, 
        n317, n317, n317, n317, n317, n317, n317, n317, n316, n316, n316, n277, 
        n275, n272, n270, n267, n265, n262, n260, n257, n255, n252, n250, n247, 
        n245, n242, n240, n238, n236, n235, n233, n72, n229, n228, n226, A[6], 
        n222, n78, n219, n96, n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n168, n168, n168, n168, n168, n168, n170, n170, n170, 
        n171, n171, n171, n159, n158, n156, n153, n150, n149, n146, n144, n142, 
        n140, n70, n68, n135, n133, n131, n130, n126, n124, n123, n120, n93, 
        n118, n91, n114, n113, n111, n110, n108, n105, n102, n99, n212, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n298, n298, n299, n299, 
        n299, n299, n300, n300, n300, n300, n300, n301, n277, n274, n272, n269, 
        n267, n264, n262, n259, n257, n254, n252, n249, n247, n244, n242, n239, 
        n238, n236, n235, n232, n71, n230, n228, n225, A[6], n221, n80, n218, 
        n96, n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n185, n185, n185, n185, n184, n184, n184, n184, n184, n184, n184, n160, 
        n158, n155, n152, n150, n149, n147, n145, n142, n139, n70, n68, n135, 
        n133, n132, n130, n127, n124, n122, n92, n119, n118, n116, n115, n113, 
        n111, n110, n109, n106, n103, n100, n213, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[10][2] , 
        \select_array[10][1] , \select_array[10][0] }), .Y({
        \array_mux_out[10][63] , \array_mux_out[10][62] , 
        \array_mux_out[10][61] , \array_mux_out[10][60] , 
        \array_mux_out[10][59] , \array_mux_out[10][58] , 
        \array_mux_out[10][57] , \array_mux_out[10][56] , 
        \array_mux_out[10][55] , \array_mux_out[10][54] , 
        \array_mux_out[10][53] , \array_mux_out[10][52] , 
        \array_mux_out[10][51] , \array_mux_out[10][50] , 
        \array_mux_out[10][49] , \array_mux_out[10][48] , 
        \array_mux_out[10][47] , \array_mux_out[10][46] , 
        \array_mux_out[10][45] , \array_mux_out[10][44] , 
        \array_mux_out[10][43] , \array_mux_out[10][42] , 
        \array_mux_out[10][41] , \array_mux_out[10][40] , 
        \array_mux_out[10][39] , \array_mux_out[10][38] , 
        \array_mux_out[10][37] , \array_mux_out[10][36] , 
        \array_mux_out[10][35] , \array_mux_out[10][34] , 
        \array_mux_out[10][33] , \array_mux_out[10][32] , 
        \array_mux_out[10][31] , \array_mux_out[10][30] , 
        \array_mux_out[10][29] , \array_mux_out[10][28] , 
        \array_mux_out[10][27] , \array_mux_out[10][26] , 
        \array_mux_out[10][25] , \array_mux_out[10][24] , 
        \array_mux_out[10][23] , \array_mux_out[10][22] , 
        \array_mux_out[10][21] , \array_mux_out[10][20] , 
        \array_mux_out[10][19] , \array_mux_out[10][18] , 
        \array_mux_out[10][17] , \array_mux_out[10][16] , 
        \array_mux_out[10][15] , \array_mux_out[10][14] , 
        \array_mux_out[10][13] , \array_mux_out[10][12] , 
        \array_mux_out[10][11] , \array_mux_out[10][10] , 
        \array_mux_out[10][9] , \array_mux_out[10][8] , \array_mux_out[10][7] , 
        \array_mux_out[10][6] , \array_mux_out[10][5] , \array_mux_out[10][4] , 
        \array_mux_out[10][3] , \array_mux_out[10][2] , \array_mux_out[10][1] , 
        \array_mux_out[10][0] }) );
  P4_ADDER_N64_6 adder_10 ( .A({\array_mux_out[10][63] , 
        \array_mux_out[10][62] , \array_mux_out[10][61] , 
        \array_mux_out[10][60] , \array_mux_out[10][59] , 
        \array_mux_out[10][58] , \array_mux_out[10][57] , 
        \array_mux_out[10][56] , \array_mux_out[10][55] , 
        \array_mux_out[10][54] , \array_mux_out[10][53] , 
        \array_mux_out[10][52] , \array_mux_out[10][51] , 
        \array_mux_out[10][50] , \array_mux_out[10][49] , 
        \array_mux_out[10][48] , \array_mux_out[10][47] , 
        \array_mux_out[10][46] , \array_mux_out[10][45] , 
        \array_mux_out[10][44] , \array_mux_out[10][43] , 
        \array_mux_out[10][42] , \array_mux_out[10][41] , 
        \array_mux_out[10][40] , \array_mux_out[10][39] , 
        \array_mux_out[10][38] , \array_mux_out[10][37] , 
        \array_mux_out[10][36] , \array_mux_out[10][35] , 
        \array_mux_out[10][34] , \array_mux_out[10][33] , 
        \array_mux_out[10][32] , \array_mux_out[10][31] , 
        \array_mux_out[10][30] , \array_mux_out[10][29] , 
        \array_mux_out[10][28] , \array_mux_out[10][27] , 
        \array_mux_out[10][26] , \array_mux_out[10][25] , 
        \array_mux_out[10][24] , \array_mux_out[10][23] , 
        \array_mux_out[10][22] , \array_mux_out[10][21] , 
        \array_mux_out[10][20] , \array_mux_out[10][19] , 
        \array_mux_out[10][18] , \array_mux_out[10][17] , 
        \array_mux_out[10][16] , \array_mux_out[10][15] , 
        \array_mux_out[10][14] , \array_mux_out[10][13] , 
        \array_mux_out[10][12] , \array_mux_out[10][11] , 
        \array_mux_out[10][10] , \array_mux_out[10][9] , 
        \array_mux_out[10][8] , \array_mux_out[10][7] , \array_mux_out[10][6] , 
        \array_mux_out[10][5] , \array_mux_out[10][4] , \array_mux_out[10][3] , 
        \array_mux_out[10][2] , \array_mux_out[10][1] , \array_mux_out[10][0] }), .B({\result_array[9][63] , \result_array[9][62] , \result_array[9][61] , 
        \result_array[9][60] , \result_array[9][59] , \result_array[9][58] , 
        \result_array[9][57] , \result_array[9][56] , \result_array[9][55] , 
        \result_array[9][54] , \result_array[9][53] , \result_array[9][52] , 
        \result_array[9][51] , \result_array[9][50] , \result_array[9][49] , 
        \result_array[9][48] , \result_array[9][47] , \result_array[9][46] , 
        \result_array[9][45] , \result_array[9][44] , \result_array[9][43] , 
        \result_array[9][42] , \result_array[9][41] , \result_array[9][40] , 
        \result_array[9][39] , \result_array[9][38] , \result_array[9][37] , 
        \result_array[9][36] , \result_array[9][35] , \result_array[9][34] , 
        \result_array[9][33] , \result_array[9][32] , \result_array[9][31] , 
        \result_array[9][30] , \result_array[9][29] , \result_array[9][28] , 
        \result_array[9][27] , \result_array[9][26] , \result_array[9][25] , 
        \result_array[9][24] , \result_array[9][23] , \result_array[9][22] , 
        \result_array[9][21] , \result_array[9][20] , \result_array[9][19] , 
        \result_array[9][18] , \result_array[9][17] , \result_array[9][16] , 
        \result_array[9][15] , \result_array[9][14] , \result_array[9][13] , 
        \result_array[9][12] , \result_array[9][11] , \result_array[9][10] , 
        \result_array[9][9] , \result_array[9][8] , \result_array[9][7] , 
        \result_array[9][6] , \result_array[9][5] , \result_array[9][4] , 
        \result_array[9][3] , \result_array[9][2] , \result_array[9][1] , 
        \result_array[9][0] }), .Cin(1'b0), .S({\result_array[10][63] , 
        \result_array[10][62] , \result_array[10][61] , \result_array[10][60] , 
        \result_array[10][59] , \result_array[10][58] , \result_array[10][57] , 
        \result_array[10][56] , \result_array[10][55] , \result_array[10][54] , 
        \result_array[10][53] , \result_array[10][52] , \result_array[10][51] , 
        \result_array[10][50] , \result_array[10][49] , \result_array[10][48] , 
        \result_array[10][47] , \result_array[10][46] , \result_array[10][45] , 
        \result_array[10][44] , \result_array[10][43] , \result_array[10][42] , 
        \result_array[10][41] , \result_array[10][40] , \result_array[10][39] , 
        \result_array[10][38] , \result_array[10][37] , \result_array[10][36] , 
        \result_array[10][35] , \result_array[10][34] , \result_array[10][33] , 
        \result_array[10][32] , \result_array[10][31] , \result_array[10][30] , 
        \result_array[10][29] , \result_array[10][28] , \result_array[10][27] , 
        \result_array[10][26] , \result_array[10][25] , \result_array[10][24] , 
        \result_array[10][23] , \result_array[10][22] , \result_array[10][21] , 
        \result_array[10][20] , \result_array[10][19] , \result_array[10][18] , 
        \result_array[10][17] , \result_array[10][16] , \result_array[10][15] , 
        \result_array[10][14] , \result_array[10][13] , \result_array[10][12] , 
        \result_array[10][11] , \result_array[10][10] , \result_array[10][9] , 
        \result_array[10][8] , \result_array[10][7] , \result_array[10][6] , 
        \result_array[10][5] , \result_array[10][4] , \result_array[10][3] , 
        \result_array[10][2] , \result_array[10][1] , \result_array[10][0] })
         );
  Booth_Encoder_5 booth_j_11 ( .i(B[23:21]), .o({\select_array[11][2] , 
        \select_array[11][1] , \select_array[11][0] }) );
  MUX_booth_N64_5 mux_j_11 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n320, n320, 
        n320, n320, n320, n320, n319, n319, n319, n319, n319, n277, n275, n272, 
        n270, n267, n265, n262, n260, n257, n255, n252, n250, n247, n245, n242, 
        n240, n238, n236, n235, n233, n71, n230, n228, n226, A[6], n222, n81, 
        n219, n96, n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n165, n165, n165, n165, n167, n167, n168, n168, n168, 
        n168, n159, n157, n155, n153, n150, n149, n146, n145, n142, n140, n138, 
        n68, n135, n133, n131, n129, n126, n124, n123, n92, n93, n118, n91, 
        n114, n113, n111, n110, n108, n105, n102, n99, n212, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n296, n296, n296, n296, 
        n296, n297, n297, n297, n297, n297, n277, n274, n272, n270, n267, n264, 
        n262, n260, n257, n254, n252, n250, n247, n244, n242, n240, n238, n237, 
        n235, n233, n72, n229, n228, n226, A[6], n221, n79, n219, n96, n216, 
        n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n187, n187, n187, n187, n187, n187, n186, n186, n186, n160, n157, n155, 
        n153, n94, n149, n147, n144, n142, n139, n70, n69, n135, n133, n132, 
        n130, n127, n124, n123, n92, n119, n117, n116, n114, n113, n111, n110, 
        n109, n106, n103, n100, n213, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[11][2] , 
        \select_array[11][1] , \select_array[11][0] }), .Y({
        \array_mux_out[11][63] , \array_mux_out[11][62] , 
        \array_mux_out[11][61] , \array_mux_out[11][60] , 
        \array_mux_out[11][59] , \array_mux_out[11][58] , 
        \array_mux_out[11][57] , \array_mux_out[11][56] , 
        \array_mux_out[11][55] , \array_mux_out[11][54] , 
        \array_mux_out[11][53] , \array_mux_out[11][52] , 
        \array_mux_out[11][51] , \array_mux_out[11][50] , 
        \array_mux_out[11][49] , \array_mux_out[11][48] , 
        \array_mux_out[11][47] , \array_mux_out[11][46] , 
        \array_mux_out[11][45] , \array_mux_out[11][44] , 
        \array_mux_out[11][43] , \array_mux_out[11][42] , 
        \array_mux_out[11][41] , \array_mux_out[11][40] , 
        \array_mux_out[11][39] , \array_mux_out[11][38] , 
        \array_mux_out[11][37] , \array_mux_out[11][36] , 
        \array_mux_out[11][35] , \array_mux_out[11][34] , 
        \array_mux_out[11][33] , \array_mux_out[11][32] , 
        \array_mux_out[11][31] , \array_mux_out[11][30] , 
        \array_mux_out[11][29] , \array_mux_out[11][28] , 
        \array_mux_out[11][27] , \array_mux_out[11][26] , 
        \array_mux_out[11][25] , \array_mux_out[11][24] , 
        \array_mux_out[11][23] , \array_mux_out[11][22] , 
        \array_mux_out[11][21] , \array_mux_out[11][20] , 
        \array_mux_out[11][19] , \array_mux_out[11][18] , 
        \array_mux_out[11][17] , \array_mux_out[11][16] , 
        \array_mux_out[11][15] , \array_mux_out[11][14] , 
        \array_mux_out[11][13] , \array_mux_out[11][12] , 
        \array_mux_out[11][11] , \array_mux_out[11][10] , 
        \array_mux_out[11][9] , \array_mux_out[11][8] , \array_mux_out[11][7] , 
        \array_mux_out[11][6] , \array_mux_out[11][5] , \array_mux_out[11][4] , 
        \array_mux_out[11][3] , \array_mux_out[11][2] , \array_mux_out[11][1] , 
        \array_mux_out[11][0] }) );
  P4_ADDER_N64_5 adder_11 ( .A({\array_mux_out[11][63] , 
        \array_mux_out[11][62] , \array_mux_out[11][61] , 
        \array_mux_out[11][60] , \array_mux_out[11][59] , 
        \array_mux_out[11][58] , \array_mux_out[11][57] , 
        \array_mux_out[11][56] , \array_mux_out[11][55] , 
        \array_mux_out[11][54] , \array_mux_out[11][53] , 
        \array_mux_out[11][52] , \array_mux_out[11][51] , 
        \array_mux_out[11][50] , \array_mux_out[11][49] , 
        \array_mux_out[11][48] , \array_mux_out[11][47] , 
        \array_mux_out[11][46] , \array_mux_out[11][45] , 
        \array_mux_out[11][44] , \array_mux_out[11][43] , 
        \array_mux_out[11][42] , \array_mux_out[11][41] , 
        \array_mux_out[11][40] , \array_mux_out[11][39] , 
        \array_mux_out[11][38] , \array_mux_out[11][37] , 
        \array_mux_out[11][36] , \array_mux_out[11][35] , 
        \array_mux_out[11][34] , \array_mux_out[11][33] , 
        \array_mux_out[11][32] , \array_mux_out[11][31] , 
        \array_mux_out[11][30] , \array_mux_out[11][29] , 
        \array_mux_out[11][28] , \array_mux_out[11][27] , 
        \array_mux_out[11][26] , \array_mux_out[11][25] , 
        \array_mux_out[11][24] , \array_mux_out[11][23] , 
        \array_mux_out[11][22] , \array_mux_out[11][21] , 
        \array_mux_out[11][20] , \array_mux_out[11][19] , 
        \array_mux_out[11][18] , \array_mux_out[11][17] , 
        \array_mux_out[11][16] , \array_mux_out[11][15] , 
        \array_mux_out[11][14] , \array_mux_out[11][13] , 
        \array_mux_out[11][12] , \array_mux_out[11][11] , 
        \array_mux_out[11][10] , \array_mux_out[11][9] , 
        \array_mux_out[11][8] , \array_mux_out[11][7] , \array_mux_out[11][6] , 
        \array_mux_out[11][5] , \array_mux_out[11][4] , \array_mux_out[11][3] , 
        \array_mux_out[11][2] , \array_mux_out[11][1] , \array_mux_out[11][0] }), .B({\result_array[10][63] , \result_array[10][62] , \result_array[10][61] , 
        \result_array[10][60] , \result_array[10][59] , \result_array[10][58] , 
        \result_array[10][57] , \result_array[10][56] , \result_array[10][55] , 
        \result_array[10][54] , \result_array[10][53] , \result_array[10][52] , 
        \result_array[10][51] , \result_array[10][50] , \result_array[10][49] , 
        \result_array[10][48] , \result_array[10][47] , \result_array[10][46] , 
        \result_array[10][45] , \result_array[10][44] , \result_array[10][43] , 
        \result_array[10][42] , \result_array[10][41] , \result_array[10][40] , 
        \result_array[10][39] , \result_array[10][38] , \result_array[10][37] , 
        \result_array[10][36] , \result_array[10][35] , \result_array[10][34] , 
        \result_array[10][33] , \result_array[10][32] , \result_array[10][31] , 
        \result_array[10][30] , \result_array[10][29] , \result_array[10][28] , 
        \result_array[10][27] , \result_array[10][26] , \result_array[10][25] , 
        \result_array[10][24] , \result_array[10][23] , \result_array[10][22] , 
        \result_array[10][21] , \result_array[10][20] , \result_array[10][19] , 
        \result_array[10][18] , \result_array[10][17] , \result_array[10][16] , 
        \result_array[10][15] , \result_array[10][14] , \result_array[10][13] , 
        \result_array[10][12] , \result_array[10][11] , \result_array[10][10] , 
        \result_array[10][9] , \result_array[10][8] , \result_array[10][7] , 
        \result_array[10][6] , \result_array[10][5] , \result_array[10][4] , 
        \result_array[10][3] , \result_array[10][2] , \result_array[10][1] , 
        \result_array[10][0] }), .Cin(1'b0), .S({\result_array[11][63] , 
        \result_array[11][62] , \result_array[11][61] , \result_array[11][60] , 
        \result_array[11][59] , \result_array[11][58] , \result_array[11][57] , 
        \result_array[11][56] , \result_array[11][55] , \result_array[11][54] , 
        \result_array[11][53] , \result_array[11][52] , \result_array[11][51] , 
        \result_array[11][50] , \result_array[11][49] , \result_array[11][48] , 
        \result_array[11][47] , \result_array[11][46] , \result_array[11][45] , 
        \result_array[11][44] , \result_array[11][43] , \result_array[11][42] , 
        \result_array[11][41] , \result_array[11][40] , \result_array[11][39] , 
        \result_array[11][38] , \result_array[11][37] , \result_array[11][36] , 
        \result_array[11][35] , \result_array[11][34] , \result_array[11][33] , 
        \result_array[11][32] , \result_array[11][31] , \result_array[11][30] , 
        \result_array[11][29] , \result_array[11][28] , \result_array[11][27] , 
        \result_array[11][26] , \result_array[11][25] , \result_array[11][24] , 
        \result_array[11][23] , \result_array[11][22] , \result_array[11][21] , 
        \result_array[11][20] , \result_array[11][19] , \result_array[11][18] , 
        \result_array[11][17] , \result_array[11][16] , \result_array[11][15] , 
        \result_array[11][14] , \result_array[11][13] , \result_array[11][12] , 
        \result_array[11][11] , \result_array[11][10] , \result_array[11][9] , 
        \result_array[11][8] , \result_array[11][7] , \result_array[11][6] , 
        \result_array[11][5] , \result_array[11][4] , \result_array[11][3] , 
        \result_array[11][2] , \result_array[11][1] , \result_array[11][0] })
         );
  Booth_Encoder_4 booth_j_12 ( .i(B[25:23]), .o({\select_array[12][2] , 
        \select_array[12][1] , \select_array[12][0] }) );
  MUX_booth_N64_4 mux_j_12 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n323, n323, 
        n322, n322, n322, n322, n322, n322, n322, n278, n275, n272, n270, n268, 
        n265, n262, n260, n258, n255, n252, n250, n248, n245, n242, n240, n238, 
        n236, n235, n233, n231, n229, n228, n226, n224, n222, n83, n219, n96, 
        n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n164, n164, n165, n165, n165, n165, n165, n165, n159, 
        n158, n155, n153, n94, n149, n146, n144, n142, n140, n138, n68, n135, 
        n133, n131, n129, n126, n124, n123, n120, n93, n118, n91, n115, n113, 
        n111, n110, n108, n105, n102, n99, n212, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n294, n295, n295, n295, 
        n295, n296, n296, n296, n277, n275, n272, n270, n267, n265, n262, n260, 
        n257, n255, n252, n250, n247, n245, n242, n240, n238, n236, n235, n233, 
        n71, n230, n228, n226, A[6], n222, n84, n219, n96, n216, n97, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n189, n188, n188, n188, n188, n188, n188, n161, n158, n156, n153, n150, 
        n149, n147, n145, n142, n139, n70, n137, n135, n133, n62, n130, n128, 
        n124, n123, n92, n93, n117, n91, n114, n113, n65, n110, n109, n107, 
        n104, n101, n214, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[12][2] , 
        \select_array[12][1] , \select_array[12][0] }), .Y({
        \array_mux_out[12][63] , \array_mux_out[12][62] , 
        \array_mux_out[12][61] , \array_mux_out[12][60] , 
        \array_mux_out[12][59] , \array_mux_out[12][58] , 
        \array_mux_out[12][57] , \array_mux_out[12][56] , 
        \array_mux_out[12][55] , \array_mux_out[12][54] , 
        \array_mux_out[12][53] , \array_mux_out[12][52] , 
        \array_mux_out[12][51] , \array_mux_out[12][50] , 
        \array_mux_out[12][49] , \array_mux_out[12][48] , 
        \array_mux_out[12][47] , \array_mux_out[12][46] , 
        \array_mux_out[12][45] , \array_mux_out[12][44] , 
        \array_mux_out[12][43] , \array_mux_out[12][42] , 
        \array_mux_out[12][41] , \array_mux_out[12][40] , 
        \array_mux_out[12][39] , \array_mux_out[12][38] , 
        \array_mux_out[12][37] , \array_mux_out[12][36] , 
        \array_mux_out[12][35] , \array_mux_out[12][34] , 
        \array_mux_out[12][33] , \array_mux_out[12][32] , 
        \array_mux_out[12][31] , \array_mux_out[12][30] , 
        \array_mux_out[12][29] , \array_mux_out[12][28] , 
        \array_mux_out[12][27] , \array_mux_out[12][26] , 
        \array_mux_out[12][25] , \array_mux_out[12][24] , 
        \array_mux_out[12][23] , \array_mux_out[12][22] , 
        \array_mux_out[12][21] , \array_mux_out[12][20] , 
        \array_mux_out[12][19] , \array_mux_out[12][18] , 
        \array_mux_out[12][17] , \array_mux_out[12][16] , 
        \array_mux_out[12][15] , \array_mux_out[12][14] , 
        \array_mux_out[12][13] , \array_mux_out[12][12] , 
        \array_mux_out[12][11] , \array_mux_out[12][10] , 
        \array_mux_out[12][9] , \array_mux_out[12][8] , \array_mux_out[12][7] , 
        \array_mux_out[12][6] , \array_mux_out[12][5] , \array_mux_out[12][4] , 
        \array_mux_out[12][3] , \array_mux_out[12][2] , \array_mux_out[12][1] , 
        \array_mux_out[12][0] }) );
  P4_ADDER_N64_4 adder_12 ( .A({\array_mux_out[12][63] , 
        \array_mux_out[12][62] , \array_mux_out[12][61] , 
        \array_mux_out[12][60] , \array_mux_out[12][59] , 
        \array_mux_out[12][58] , \array_mux_out[12][57] , 
        \array_mux_out[12][56] , \array_mux_out[12][55] , 
        \array_mux_out[12][54] , \array_mux_out[12][53] , 
        \array_mux_out[12][52] , \array_mux_out[12][51] , 
        \array_mux_out[12][50] , \array_mux_out[12][49] , 
        \array_mux_out[12][48] , \array_mux_out[12][47] , 
        \array_mux_out[12][46] , \array_mux_out[12][45] , 
        \array_mux_out[12][44] , \array_mux_out[12][43] , 
        \array_mux_out[12][42] , \array_mux_out[12][41] , 
        \array_mux_out[12][40] , \array_mux_out[12][39] , 
        \array_mux_out[12][38] , \array_mux_out[12][37] , 
        \array_mux_out[12][36] , \array_mux_out[12][35] , 
        \array_mux_out[12][34] , \array_mux_out[12][33] , 
        \array_mux_out[12][32] , \array_mux_out[12][31] , 
        \array_mux_out[12][30] , \array_mux_out[12][29] , 
        \array_mux_out[12][28] , \array_mux_out[12][27] , 
        \array_mux_out[12][26] , \array_mux_out[12][25] , 
        \array_mux_out[12][24] , \array_mux_out[12][23] , 
        \array_mux_out[12][22] , \array_mux_out[12][21] , 
        \array_mux_out[12][20] , \array_mux_out[12][19] , 
        \array_mux_out[12][18] , \array_mux_out[12][17] , 
        \array_mux_out[12][16] , \array_mux_out[12][15] , 
        \array_mux_out[12][14] , \array_mux_out[12][13] , 
        \array_mux_out[12][12] , \array_mux_out[12][11] , 
        \array_mux_out[12][10] , \array_mux_out[12][9] , 
        \array_mux_out[12][8] , \array_mux_out[12][7] , \array_mux_out[12][6] , 
        \array_mux_out[12][5] , \array_mux_out[12][4] , \array_mux_out[12][3] , 
        \array_mux_out[12][2] , \array_mux_out[12][1] , \array_mux_out[12][0] }), .B({\result_array[11][63] , \result_array[11][62] , \result_array[11][61] , 
        \result_array[11][60] , \result_array[11][59] , \result_array[11][58] , 
        \result_array[11][57] , \result_array[11][56] , \result_array[11][55] , 
        \result_array[11][54] , \result_array[11][53] , \result_array[11][52] , 
        \result_array[11][51] , \result_array[11][50] , \result_array[11][49] , 
        \result_array[11][48] , \result_array[11][47] , \result_array[11][46] , 
        \result_array[11][45] , \result_array[11][44] , \result_array[11][43] , 
        \result_array[11][42] , \result_array[11][41] , \result_array[11][40] , 
        \result_array[11][39] , \result_array[11][38] , \result_array[11][37] , 
        \result_array[11][36] , \result_array[11][35] , \result_array[11][34] , 
        \result_array[11][33] , \result_array[11][32] , \result_array[11][31] , 
        \result_array[11][30] , \result_array[11][29] , \result_array[11][28] , 
        \result_array[11][27] , \result_array[11][26] , \result_array[11][25] , 
        \result_array[11][24] , \result_array[11][23] , \result_array[11][22] , 
        \result_array[11][21] , \result_array[11][20] , \result_array[11][19] , 
        \result_array[11][18] , \result_array[11][17] , \result_array[11][16] , 
        \result_array[11][15] , \result_array[11][14] , \result_array[11][13] , 
        \result_array[11][12] , \result_array[11][11] , \result_array[11][10] , 
        \result_array[11][9] , \result_array[11][8] , \result_array[11][7] , 
        \result_array[11][6] , \result_array[11][5] , \result_array[11][4] , 
        \result_array[11][3] , \result_array[11][2] , \result_array[11][1] , 
        \result_array[11][0] }), .Cin(1'b0), .S({\result_array[12][63] , 
        \result_array[12][62] , \result_array[12][61] , \result_array[12][60] , 
        \result_array[12][59] , \result_array[12][58] , \result_array[12][57] , 
        \result_array[12][56] , \result_array[12][55] , \result_array[12][54] , 
        \result_array[12][53] , \result_array[12][52] , \result_array[12][51] , 
        \result_array[12][50] , \result_array[12][49] , \result_array[12][48] , 
        \result_array[12][47] , \result_array[12][46] , \result_array[12][45] , 
        \result_array[12][44] , \result_array[12][43] , \result_array[12][42] , 
        \result_array[12][41] , \result_array[12][40] , \result_array[12][39] , 
        \result_array[12][38] , \result_array[12][37] , \result_array[12][36] , 
        \result_array[12][35] , \result_array[12][34] , \result_array[12][33] , 
        \result_array[12][32] , \result_array[12][31] , \result_array[12][30] , 
        \result_array[12][29] , \result_array[12][28] , \result_array[12][27] , 
        \result_array[12][26] , \result_array[12][25] , \result_array[12][24] , 
        \result_array[12][23] , \result_array[12][22] , \result_array[12][21] , 
        \result_array[12][20] , \result_array[12][19] , \result_array[12][18] , 
        \result_array[12][17] , \result_array[12][16] , \result_array[12][15] , 
        \result_array[12][14] , \result_array[12][13] , \result_array[12][12] , 
        \result_array[12][11] , \result_array[12][10] , \result_array[12][9] , 
        \result_array[12][8] , \result_array[12][7] , \result_array[12][6] , 
        \result_array[12][5] , \result_array[12][4] , \result_array[12][3] , 
        \result_array[12][2] , \result_array[12][1] , \result_array[12][0] })
         );
  Booth_Encoder_3 booth_j_13 ( .i(B[27:25]), .o({\select_array[13][2] , 
        \select_array[13][1] , \select_array[13][0] }) );
  MUX_booth_N64_3 mux_j_13 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n303, n305, 
        n303, n323, n323, n323, n323, n278, n276, n272, n271, n268, n266, n262, 
        n261, n258, n256, n252, n251, n248, n246, n242, n241, n238, n237, n235, 
        n234, n71, n230, n228, n227, n224, n223, n85, n220, n96, n216, n97, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n180, n180, n180, n179, n180, n181, n159, n157, n155, 
        n153, n150, n149, n146, n145, n142, n139, n70, n68, n135, n133, n131, 
        n129, n126, n124, n122, n92, n93, n118, n91, n114, n113, n111, n110, 
        n108, n105, n102, n99, n212, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n294, n294, n294, n294, 
        n294, n294, n277, n275, n272, n270, n267, n265, n262, n260, n257, n255, 
        n252, n250, n247, n245, n242, n240, n238, n236, n235, n233, n231, n229, 
        n228, n226, A[6], n222, n82, n219, n96, n216, n97, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n189, n183, n189, n189, n189, n161, n158, n155, n152, n150, n66, n147, 
        n144, n142, n139, n138, n137, n135, n133, n62, n130, n128, n124, n122, 
        n120, n93, n117, n91, n114, n113, n65, n110, n109, n107, n104, n101, 
        n214, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[13][2] , 
        \select_array[13][1] , \select_array[13][0] }), .Y({
        \array_mux_out[13][63] , \array_mux_out[13][62] , 
        \array_mux_out[13][61] , \array_mux_out[13][60] , 
        \array_mux_out[13][59] , \array_mux_out[13][58] , 
        \array_mux_out[13][57] , \array_mux_out[13][56] , 
        \array_mux_out[13][55] , \array_mux_out[13][54] , 
        \array_mux_out[13][53] , \array_mux_out[13][52] , 
        \array_mux_out[13][51] , \array_mux_out[13][50] , 
        \array_mux_out[13][49] , \array_mux_out[13][48] , 
        \array_mux_out[13][47] , \array_mux_out[13][46] , 
        \array_mux_out[13][45] , \array_mux_out[13][44] , 
        \array_mux_out[13][43] , \array_mux_out[13][42] , 
        \array_mux_out[13][41] , \array_mux_out[13][40] , 
        \array_mux_out[13][39] , \array_mux_out[13][38] , 
        \array_mux_out[13][37] , \array_mux_out[13][36] , 
        \array_mux_out[13][35] , \array_mux_out[13][34] , 
        \array_mux_out[13][33] , \array_mux_out[13][32] , 
        \array_mux_out[13][31] , \array_mux_out[13][30] , 
        \array_mux_out[13][29] , \array_mux_out[13][28] , 
        \array_mux_out[13][27] , \array_mux_out[13][26] , 
        \array_mux_out[13][25] , \array_mux_out[13][24] , 
        \array_mux_out[13][23] , \array_mux_out[13][22] , 
        \array_mux_out[13][21] , \array_mux_out[13][20] , 
        \array_mux_out[13][19] , \array_mux_out[13][18] , 
        \array_mux_out[13][17] , \array_mux_out[13][16] , 
        \array_mux_out[13][15] , \array_mux_out[13][14] , 
        \array_mux_out[13][13] , \array_mux_out[13][12] , 
        \array_mux_out[13][11] , \array_mux_out[13][10] , 
        \array_mux_out[13][9] , \array_mux_out[13][8] , \array_mux_out[13][7] , 
        \array_mux_out[13][6] , \array_mux_out[13][5] , \array_mux_out[13][4] , 
        \array_mux_out[13][3] , \array_mux_out[13][2] , \array_mux_out[13][1] , 
        \array_mux_out[13][0] }) );
  P4_ADDER_N64_3 adder_13 ( .A({\array_mux_out[13][63] , 
        \array_mux_out[13][62] , \array_mux_out[13][61] , 
        \array_mux_out[13][60] , \array_mux_out[13][59] , 
        \array_mux_out[13][58] , \array_mux_out[13][57] , 
        \array_mux_out[13][56] , \array_mux_out[13][55] , 
        \array_mux_out[13][54] , \array_mux_out[13][53] , 
        \array_mux_out[13][52] , \array_mux_out[13][51] , 
        \array_mux_out[13][50] , \array_mux_out[13][49] , 
        \array_mux_out[13][48] , \array_mux_out[13][47] , 
        \array_mux_out[13][46] , \array_mux_out[13][45] , 
        \array_mux_out[13][44] , \array_mux_out[13][43] , 
        \array_mux_out[13][42] , \array_mux_out[13][41] , 
        \array_mux_out[13][40] , \array_mux_out[13][39] , 
        \array_mux_out[13][38] , \array_mux_out[13][37] , 
        \array_mux_out[13][36] , \array_mux_out[13][35] , 
        \array_mux_out[13][34] , \array_mux_out[13][33] , 
        \array_mux_out[13][32] , \array_mux_out[13][31] , 
        \array_mux_out[13][30] , \array_mux_out[13][29] , 
        \array_mux_out[13][28] , \array_mux_out[13][27] , 
        \array_mux_out[13][26] , \array_mux_out[13][25] , 
        \array_mux_out[13][24] , \array_mux_out[13][23] , 
        \array_mux_out[13][22] , \array_mux_out[13][21] , 
        \array_mux_out[13][20] , \array_mux_out[13][19] , 
        \array_mux_out[13][18] , \array_mux_out[13][17] , 
        \array_mux_out[13][16] , \array_mux_out[13][15] , 
        \array_mux_out[13][14] , \array_mux_out[13][13] , 
        \array_mux_out[13][12] , \array_mux_out[13][11] , 
        \array_mux_out[13][10] , \array_mux_out[13][9] , 
        \array_mux_out[13][8] , \array_mux_out[13][7] , \array_mux_out[13][6] , 
        \array_mux_out[13][5] , \array_mux_out[13][4] , \array_mux_out[13][3] , 
        \array_mux_out[13][2] , \array_mux_out[13][1] , \array_mux_out[13][0] }), .B({\result_array[12][63] , \result_array[12][62] , \result_array[12][61] , 
        \result_array[12][60] , \result_array[12][59] , \result_array[12][58] , 
        \result_array[12][57] , \result_array[12][56] , \result_array[12][55] , 
        \result_array[12][54] , \result_array[12][53] , \result_array[12][52] , 
        \result_array[12][51] , \result_array[12][50] , \result_array[12][49] , 
        \result_array[12][48] , \result_array[12][47] , \result_array[12][46] , 
        \result_array[12][45] , \result_array[12][44] , \result_array[12][43] , 
        \result_array[12][42] , \result_array[12][41] , \result_array[12][40] , 
        \result_array[12][39] , \result_array[12][38] , \result_array[12][37] , 
        \result_array[12][36] , \result_array[12][35] , \result_array[12][34] , 
        \result_array[12][33] , \result_array[12][32] , \result_array[12][31] , 
        \result_array[12][30] , \result_array[12][29] , \result_array[12][28] , 
        \result_array[12][27] , \result_array[12][26] , \result_array[12][25] , 
        \result_array[12][24] , \result_array[12][23] , \result_array[12][22] , 
        \result_array[12][21] , \result_array[12][20] , \result_array[12][19] , 
        \result_array[12][18] , \result_array[12][17] , \result_array[12][16] , 
        \result_array[12][15] , \result_array[12][14] , \result_array[12][13] , 
        \result_array[12][12] , \result_array[12][11] , \result_array[12][10] , 
        \result_array[12][9] , \result_array[12][8] , \result_array[12][7] , 
        \result_array[12][6] , \result_array[12][5] , \result_array[12][4] , 
        \result_array[12][3] , \result_array[12][2] , \result_array[12][1] , 
        \result_array[12][0] }), .Cin(1'b0), .S({\result_array[13][63] , 
        \result_array[13][62] , \result_array[13][61] , \result_array[13][60] , 
        \result_array[13][59] , \result_array[13][58] , \result_array[13][57] , 
        \result_array[13][56] , \result_array[13][55] , \result_array[13][54] , 
        \result_array[13][53] , \result_array[13][52] , \result_array[13][51] , 
        \result_array[13][50] , \result_array[13][49] , \result_array[13][48] , 
        \result_array[13][47] , \result_array[13][46] , \result_array[13][45] , 
        \result_array[13][44] , \result_array[13][43] , \result_array[13][42] , 
        \result_array[13][41] , \result_array[13][40] , \result_array[13][39] , 
        \result_array[13][38] , \result_array[13][37] , \result_array[13][36] , 
        \result_array[13][35] , \result_array[13][34] , \result_array[13][33] , 
        \result_array[13][32] , \result_array[13][31] , \result_array[13][30] , 
        \result_array[13][29] , \result_array[13][28] , \result_array[13][27] , 
        \result_array[13][26] , \result_array[13][25] , \result_array[13][24] , 
        \result_array[13][23] , \result_array[13][22] , \result_array[13][21] , 
        \result_array[13][20] , \result_array[13][19] , \result_array[13][18] , 
        \result_array[13][17] , \result_array[13][16] , \result_array[13][15] , 
        \result_array[13][14] , \result_array[13][13] , \result_array[13][12] , 
        \result_array[13][11] , \result_array[13][10] , \result_array[13][9] , 
        \result_array[13][8] , \result_array[13][7] , \result_array[13][6] , 
        \result_array[13][5] , \result_array[13][4] , \result_array[13][3] , 
        \result_array[13][2] , \result_array[13][1] , \result_array[13][0] })
         );
  Booth_Encoder_2 booth_j_14 ( .i(B[29:27]), .o({\select_array[14][2] , 
        \select_array[14][1] , \select_array[14][0] }) );
  MUX_booth_N64_2 mux_j_14 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n304, n304, 
        n304, n304, n305, n278, n276, n273, n271, n268, n266, n263, n261, n258, 
        n256, n253, n251, n248, n246, n243, n241, n238, n237, n235, n234, n231, 
        n229, n228, n227, n224, n223, n87, n220, n96, n216, n97, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n179, n179, n179, n179, n159, n157, n155, n153, n94, 
        n149, n146, n144, n142, n140, n138, n68, n135, n133, n131, n129, n126, 
        n124, n122, n120, n93, n117, n91, n114, n113, n111, n110, n108, n105, 
        n102, n99, n212, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n295, n295, n295, n295, 
        n277, n275, n272, n270, n267, n265, n262, n260, n257, n255, n252, n250, 
        n247, n245, n242, n240, n238, n236, n235, n233, n72, n230, n228, n226, 
        A[6], n222, n86, n219, n96, n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n188, n188, n188, n161, n158, n156, n152, n150, n149, n147, n145, n142, 
        n139, n70, n137, n135, n133, n62, n130, n128, n124, n123, n92, n93, 
        n118, n91, n115, n113, n65, n110, n109, n107, n104, n101, n214, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[14][2] , 
        \select_array[14][1] , \select_array[14][0] }), .Y({
        \array_mux_out[14][63] , \array_mux_out[14][62] , 
        \array_mux_out[14][61] , \array_mux_out[14][60] , 
        \array_mux_out[14][59] , \array_mux_out[14][58] , 
        \array_mux_out[14][57] , \array_mux_out[14][56] , 
        \array_mux_out[14][55] , \array_mux_out[14][54] , 
        \array_mux_out[14][53] , \array_mux_out[14][52] , 
        \array_mux_out[14][51] , \array_mux_out[14][50] , 
        \array_mux_out[14][49] , \array_mux_out[14][48] , 
        \array_mux_out[14][47] , \array_mux_out[14][46] , 
        \array_mux_out[14][45] , \array_mux_out[14][44] , 
        \array_mux_out[14][43] , \array_mux_out[14][42] , 
        \array_mux_out[14][41] , \array_mux_out[14][40] , 
        \array_mux_out[14][39] , \array_mux_out[14][38] , 
        \array_mux_out[14][37] , \array_mux_out[14][36] , 
        \array_mux_out[14][35] , \array_mux_out[14][34] , 
        \array_mux_out[14][33] , \array_mux_out[14][32] , 
        \array_mux_out[14][31] , \array_mux_out[14][30] , 
        \array_mux_out[14][29] , \array_mux_out[14][28] , 
        \array_mux_out[14][27] , \array_mux_out[14][26] , 
        \array_mux_out[14][25] , \array_mux_out[14][24] , 
        \array_mux_out[14][23] , \array_mux_out[14][22] , 
        \array_mux_out[14][21] , \array_mux_out[14][20] , 
        \array_mux_out[14][19] , \array_mux_out[14][18] , 
        \array_mux_out[14][17] , \array_mux_out[14][16] , 
        \array_mux_out[14][15] , \array_mux_out[14][14] , 
        \array_mux_out[14][13] , \array_mux_out[14][12] , 
        \array_mux_out[14][11] , \array_mux_out[14][10] , 
        \array_mux_out[14][9] , \array_mux_out[14][8] , \array_mux_out[14][7] , 
        \array_mux_out[14][6] , \array_mux_out[14][5] , \array_mux_out[14][4] , 
        \array_mux_out[14][3] , \array_mux_out[14][2] , \array_mux_out[14][1] , 
        \array_mux_out[14][0] }) );
  P4_ADDER_N64_2 adder_14 ( .A({\array_mux_out[14][63] , 
        \array_mux_out[14][62] , \array_mux_out[14][61] , 
        \array_mux_out[14][60] , \array_mux_out[14][59] , 
        \array_mux_out[14][58] , \array_mux_out[14][57] , 
        \array_mux_out[14][56] , \array_mux_out[14][55] , 
        \array_mux_out[14][54] , \array_mux_out[14][53] , 
        \array_mux_out[14][52] , \array_mux_out[14][51] , 
        \array_mux_out[14][50] , \array_mux_out[14][49] , 
        \array_mux_out[14][48] , \array_mux_out[14][47] , 
        \array_mux_out[14][46] , \array_mux_out[14][45] , 
        \array_mux_out[14][44] , \array_mux_out[14][43] , 
        \array_mux_out[14][42] , \array_mux_out[14][41] , 
        \array_mux_out[14][40] , \array_mux_out[14][39] , 
        \array_mux_out[14][38] , \array_mux_out[14][37] , 
        \array_mux_out[14][36] , \array_mux_out[14][35] , 
        \array_mux_out[14][34] , \array_mux_out[14][33] , 
        \array_mux_out[14][32] , \array_mux_out[14][31] , 
        \array_mux_out[14][30] , \array_mux_out[14][29] , 
        \array_mux_out[14][28] , \array_mux_out[14][27] , 
        \array_mux_out[14][26] , \array_mux_out[14][25] , 
        \array_mux_out[14][24] , \array_mux_out[14][23] , 
        \array_mux_out[14][22] , \array_mux_out[14][21] , 
        \array_mux_out[14][20] , \array_mux_out[14][19] , 
        \array_mux_out[14][18] , \array_mux_out[14][17] , 
        \array_mux_out[14][16] , \array_mux_out[14][15] , 
        \array_mux_out[14][14] , \array_mux_out[14][13] , 
        \array_mux_out[14][12] , \array_mux_out[14][11] , 
        \array_mux_out[14][10] , \array_mux_out[14][9] , 
        \array_mux_out[14][8] , \array_mux_out[14][7] , \array_mux_out[14][6] , 
        \array_mux_out[14][5] , \array_mux_out[14][4] , \array_mux_out[14][3] , 
        \array_mux_out[14][2] , \array_mux_out[14][1] , \array_mux_out[14][0] }), .B({\result_array[13][63] , \result_array[13][62] , \result_array[13][61] , 
        \result_array[13][60] , \result_array[13][59] , \result_array[13][58] , 
        \result_array[13][57] , \result_array[13][56] , \result_array[13][55] , 
        \result_array[13][54] , \result_array[13][53] , \result_array[13][52] , 
        \result_array[13][51] , \result_array[13][50] , \result_array[13][49] , 
        \result_array[13][48] , \result_array[13][47] , \result_array[13][46] , 
        \result_array[13][45] , \result_array[13][44] , \result_array[13][43] , 
        \result_array[13][42] , \result_array[13][41] , \result_array[13][40] , 
        \result_array[13][39] , \result_array[13][38] , \result_array[13][37] , 
        \result_array[13][36] , \result_array[13][35] , \result_array[13][34] , 
        \result_array[13][33] , \result_array[13][32] , \result_array[13][31] , 
        \result_array[13][30] , \result_array[13][29] , \result_array[13][28] , 
        \result_array[13][27] , \result_array[13][26] , \result_array[13][25] , 
        \result_array[13][24] , \result_array[13][23] , \result_array[13][22] , 
        \result_array[13][21] , \result_array[13][20] , \result_array[13][19] , 
        \result_array[13][18] , \result_array[13][17] , \result_array[13][16] , 
        \result_array[13][15] , \result_array[13][14] , \result_array[13][13] , 
        \result_array[13][12] , \result_array[13][11] , \result_array[13][10] , 
        \result_array[13][9] , \result_array[13][8] , \result_array[13][7] , 
        \result_array[13][6] , \result_array[13][5] , \result_array[13][4] , 
        \result_array[13][3] , \result_array[13][2] , \result_array[13][1] , 
        \result_array[13][0] }), .Cin(1'b0), .S({\result_array[14][63] , 
        \result_array[14][62] , \result_array[14][61] , \result_array[14][60] , 
        \result_array[14][59] , \result_array[14][58] , \result_array[14][57] , 
        \result_array[14][56] , \result_array[14][55] , \result_array[14][54] , 
        \result_array[14][53] , \result_array[14][52] , \result_array[14][51] , 
        \result_array[14][50] , \result_array[14][49] , \result_array[14][48] , 
        \result_array[14][47] , \result_array[14][46] , \result_array[14][45] , 
        \result_array[14][44] , \result_array[14][43] , \result_array[14][42] , 
        \result_array[14][41] , \result_array[14][40] , \result_array[14][39] , 
        \result_array[14][38] , \result_array[14][37] , \result_array[14][36] , 
        \result_array[14][35] , \result_array[14][34] , \result_array[14][33] , 
        \result_array[14][32] , \result_array[14][31] , \result_array[14][30] , 
        \result_array[14][29] , \result_array[14][28] , \result_array[14][27] , 
        \result_array[14][26] , \result_array[14][25] , \result_array[14][24] , 
        \result_array[14][23] , \result_array[14][22] , \result_array[14][21] , 
        \result_array[14][20] , \result_array[14][19] , \result_array[14][18] , 
        \result_array[14][17] , \result_array[14][16] , \result_array[14][15] , 
        \result_array[14][14] , \result_array[14][13] , \result_array[14][12] , 
        \result_array[14][11] , \result_array[14][10] , \result_array[14][9] , 
        \result_array[14][8] , \result_array[14][7] , \result_array[14][6] , 
        \result_array[14][5] , \result_array[14][4] , \result_array[14][3] , 
        \result_array[14][2] , \result_array[14][1] , \result_array[14][0] })
         );
  Booth_Encoder_1 booth_j_15 ( .i(B[31:29]), .o({\select_array[15][2] , 
        \select_array[15][1] , \select_array[15][0] }) );
  MUX_booth_N64_1 mux_j_15 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n304, n305, 
        n304, n278, n276, n273, n271, n268, n266, n263, n261, n258, n256, n253, 
        n251, n248, n246, n243, n241, n238, n237, n235, n234, n231, n230, n228, 
        n227, n224, n223, n89, n220, n96, n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n179, n179, n159, n158, n156, n152, n94, n149, n146, 
        n145, n142, n139, n70, n68, n135, n133, n131, n130, n126, n124, n123, 
        n120, n93, n117, n91, n115, n113, n111, n110, n108, n105, n102, n99, 
        n212, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n295, n295, n277, n275, 
        n272, n270, n267, n265, n262, n260, n257, n255, n252, n250, n247, n245, 
        n242, n240, n238, n236, n235, n233, n231, n229, n228, n226, n224, n222, 
        n88, n219, n96, n216, n97, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n188, n161, n157, n155, n153, n150, n66, n147, n144, n142, n140, n138, 
        n137, n135, n133, n62, n130, n128, n124, n122, n92, n93, n118, n91, 
        n114, n113, n65, n110, n109, n107, n104, n101, n214, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .sel({\select_array[15][2] , 
        \select_array[15][1] , \select_array[15][0] }), .Y({
        \array_mux_out[15][63] , \array_mux_out[15][62] , 
        \array_mux_out[15][61] , \array_mux_out[15][60] , 
        \array_mux_out[15][59] , \array_mux_out[15][58] , 
        \array_mux_out[15][57] , \array_mux_out[15][56] , 
        \array_mux_out[15][55] , \array_mux_out[15][54] , 
        \array_mux_out[15][53] , \array_mux_out[15][52] , 
        \array_mux_out[15][51] , \array_mux_out[15][50] , 
        \array_mux_out[15][49] , \array_mux_out[15][48] , 
        \array_mux_out[15][47] , \array_mux_out[15][46] , 
        \array_mux_out[15][45] , \array_mux_out[15][44] , 
        \array_mux_out[15][43] , \array_mux_out[15][42] , 
        \array_mux_out[15][41] , \array_mux_out[15][40] , 
        \array_mux_out[15][39] , \array_mux_out[15][38] , 
        \array_mux_out[15][37] , \array_mux_out[15][36] , 
        \array_mux_out[15][35] , \array_mux_out[15][34] , 
        \array_mux_out[15][33] , \array_mux_out[15][32] , 
        \array_mux_out[15][31] , \array_mux_out[15][30] , 
        \array_mux_out[15][29] , \array_mux_out[15][28] , 
        \array_mux_out[15][27] , \array_mux_out[15][26] , 
        \array_mux_out[15][25] , \array_mux_out[15][24] , 
        \array_mux_out[15][23] , \array_mux_out[15][22] , 
        \array_mux_out[15][21] , \array_mux_out[15][20] , 
        \array_mux_out[15][19] , \array_mux_out[15][18] , 
        \array_mux_out[15][17] , \array_mux_out[15][16] , 
        \array_mux_out[15][15] , \array_mux_out[15][14] , 
        \array_mux_out[15][13] , \array_mux_out[15][12] , 
        \array_mux_out[15][11] , \array_mux_out[15][10] , 
        \array_mux_out[15][9] , \array_mux_out[15][8] , \array_mux_out[15][7] , 
        \array_mux_out[15][6] , \array_mux_out[15][5] , \array_mux_out[15][4] , 
        \array_mux_out[15][3] , \array_mux_out[15][2] , \array_mux_out[15][1] , 
        \array_mux_out[15][0] }) );
  P4_ADDER_N64_1 adder_15 ( .A({\array_mux_out[15][63] , 
        \array_mux_out[15][62] , \array_mux_out[15][61] , 
        \array_mux_out[15][60] , \array_mux_out[15][59] , 
        \array_mux_out[15][58] , \array_mux_out[15][57] , 
        \array_mux_out[15][56] , \array_mux_out[15][55] , 
        \array_mux_out[15][54] , \array_mux_out[15][53] , 
        \array_mux_out[15][52] , \array_mux_out[15][51] , 
        \array_mux_out[15][50] , \array_mux_out[15][49] , 
        \array_mux_out[15][48] , \array_mux_out[15][47] , 
        \array_mux_out[15][46] , \array_mux_out[15][45] , 
        \array_mux_out[15][44] , \array_mux_out[15][43] , 
        \array_mux_out[15][42] , \array_mux_out[15][41] , 
        \array_mux_out[15][40] , \array_mux_out[15][39] , 
        \array_mux_out[15][38] , \array_mux_out[15][37] , 
        \array_mux_out[15][36] , \array_mux_out[15][35] , 
        \array_mux_out[15][34] , \array_mux_out[15][33] , 
        \array_mux_out[15][32] , \array_mux_out[15][31] , 
        \array_mux_out[15][30] , \array_mux_out[15][29] , 
        \array_mux_out[15][28] , \array_mux_out[15][27] , 
        \array_mux_out[15][26] , \array_mux_out[15][25] , 
        \array_mux_out[15][24] , \array_mux_out[15][23] , 
        \array_mux_out[15][22] , \array_mux_out[15][21] , 
        \array_mux_out[15][20] , \array_mux_out[15][19] , 
        \array_mux_out[15][18] , \array_mux_out[15][17] , 
        \array_mux_out[15][16] , \array_mux_out[15][15] , 
        \array_mux_out[15][14] , \array_mux_out[15][13] , 
        \array_mux_out[15][12] , \array_mux_out[15][11] , 
        \array_mux_out[15][10] , \array_mux_out[15][9] , 
        \array_mux_out[15][8] , \array_mux_out[15][7] , \array_mux_out[15][6] , 
        \array_mux_out[15][5] , \array_mux_out[15][4] , \array_mux_out[15][3] , 
        \array_mux_out[15][2] , \array_mux_out[15][1] , \array_mux_out[15][0] }), .B({\result_array[14][63] , \result_array[14][62] , \result_array[14][61] , 
        \result_array[14][60] , \result_array[14][59] , \result_array[14][58] , 
        \result_array[14][57] , \result_array[14][56] , \result_array[14][55] , 
        \result_array[14][54] , \result_array[14][53] , \result_array[14][52] , 
        \result_array[14][51] , \result_array[14][50] , \result_array[14][49] , 
        \result_array[14][48] , \result_array[14][47] , \result_array[14][46] , 
        \result_array[14][45] , \result_array[14][44] , \result_array[14][43] , 
        \result_array[14][42] , \result_array[14][41] , \result_array[14][40] , 
        \result_array[14][39] , \result_array[14][38] , \result_array[14][37] , 
        \result_array[14][36] , \result_array[14][35] , \result_array[14][34] , 
        \result_array[14][33] , \result_array[14][32] , \result_array[14][31] , 
        \result_array[14][30] , \result_array[14][29] , \result_array[14][28] , 
        \result_array[14][27] , \result_array[14][26] , \result_array[14][25] , 
        \result_array[14][24] , \result_array[14][23] , \result_array[14][22] , 
        \result_array[14][21] , \result_array[14][20] , \result_array[14][19] , 
        \result_array[14][18] , \result_array[14][17] , \result_array[14][16] , 
        \result_array[14][15] , \result_array[14][14] , \result_array[14][13] , 
        \result_array[14][12] , \result_array[14][11] , \result_array[14][10] , 
        \result_array[14][9] , \result_array[14][8] , \result_array[14][7] , 
        \result_array[14][6] , \result_array[14][5] , \result_array[14][4] , 
        \result_array[14][3] , \result_array[14][2] , \result_array[14][1] , 
        \result_array[14][0] }), .Cin(1'b0), .S(S) );
  booth_mul_N32_DW01_sub_0 sub_57 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({n323, n323, n277, n274, n272, n269, n267, n264, 
        n262, n259, n257, n254, n252, n249, n247, n244, n242, n239, A[14:5], 
        n75, n218, A[2:0]}), .CI(1'b0), .DIFF({minus_A_63, minus_A}) );
  CLKBUF_X1 U7 ( .A(minus_A[7]), .Z(n61) );
  CLKBUF_X1 U8 ( .A(minus_A[18]), .Z(n58) );
  CLKBUF_X2 U9 ( .A(minus_A[19]), .Z(n135) );
  BUF_X1 U10 ( .A(A[27]), .Z(n269) );
  BUF_X2 U11 ( .A(A[21]), .Z(n254) );
  BUF_X1 U12 ( .A(A[25]), .Z(n264) );
  BUF_X1 U13 ( .A(A[10]), .Z(n71) );
  BUF_X1 U14 ( .A(A[11]), .Z(n233) );
  BUF_X2 U15 ( .A(n63), .Z(n113) );
  BUF_X1 U16 ( .A(minus_A[6]), .Z(n112) );
  BUF_X2 U17 ( .A(A[3]), .Z(n218) );
  BUF_X1 U18 ( .A(A[19]), .Z(n249) );
  BUF_X1 U19 ( .A(A[23]), .Z(n259) );
  BUF_X1 U20 ( .A(A[29]), .Z(n274) );
  BUF_X1 U21 ( .A(n334), .Z(n324) );
  BUF_X1 U22 ( .A(minus_A[1]), .Z(n101) );
  BUF_X1 U23 ( .A(A[18]), .Z(n248) );
  BUF_X1 U24 ( .A(A[30]), .Z(n278) );
  BUF_X1 U25 ( .A(n326), .Z(n310) );
  BUF_X1 U26 ( .A(A[17]), .Z(n245) );
  BUF_X1 U27 ( .A(A[29]), .Z(n275) );
  BUF_X1 U28 ( .A(A[3]), .Z(n219) );
  BUF_X1 U29 ( .A(A[3]), .Z(n220) );
  BUF_X1 U30 ( .A(A[19]), .Z(n251) );
  BUF_X1 U31 ( .A(minus_A[16]), .Z(n130) );
  BUF_X1 U32 ( .A(minus_A[21]), .Z(n70) );
  CLKBUF_X1 U33 ( .A(minus_A[11]), .Z(n59) );
  BUF_X2 U34 ( .A(minus_A[4]), .Z(n108) );
  CLKBUF_X3 U35 ( .A(minus_A[15]), .Z(n126) );
  BUF_X1 U36 ( .A(minus_A[14]), .Z(n125) );
  CLKBUF_X2 U37 ( .A(minus_A[5]), .Z(n110) );
  BUF_X2 U38 ( .A(minus_A[4]), .Z(n109) );
  CLKBUF_X1 U39 ( .A(n58), .Z(n60) );
  BUF_X1 U40 ( .A(minus_A[13]), .Z(n64) );
  CLKBUF_X1 U41 ( .A(minus_A[7]), .Z(n63) );
  BUF_X1 U42 ( .A(minus_A[0]), .Z(n213) );
  BUF_X1 U43 ( .A(minus_A[0]), .Z(n214) );
  BUF_X2 U44 ( .A(minus_A[9]), .Z(n116) );
  CLKBUF_X1 U45 ( .A(minus_A[8]), .Z(n114) );
  BUF_X1 U46 ( .A(n211), .Z(n209) );
  BUF_X4 U47 ( .A(n125), .Z(n124) );
  BUF_X4 U48 ( .A(n60), .Z(n133) );
  BUF_X1 U49 ( .A(A[10]), .Z(n72) );
  CLKBUF_X1 U50 ( .A(minus_A[28]), .Z(n153) );
  CLKBUF_X1 U51 ( .A(minus_A[17]), .Z(n62) );
  BUF_X1 U52 ( .A(A[5]), .Z(n223) );
  BUF_X1 U53 ( .A(A[5]), .Z(n221) );
  CLKBUF_X1 U54 ( .A(n111), .Z(n65) );
  CLKBUF_X1 U55 ( .A(minus_A[26]), .Z(n66) );
  BUF_X1 U56 ( .A(A[0]), .Z(n67) );
  BUF_X4 U57 ( .A(A[13]), .Z(n236) );
  BUF_X1 U58 ( .A(A[7]), .Z(n225) );
  BUF_X2 U59 ( .A(minus_A[8]), .Z(n115) );
  CLKBUF_X1 U60 ( .A(minus_A[10]), .Z(n117) );
  CLKBUF_X1 U61 ( .A(n136), .Z(n137) );
  BUF_X1 U62 ( .A(A[11]), .Z(n232) );
  BUF_X2 U63 ( .A(minus_A[11]), .Z(n119) );
  CLKBUF_X1 U64 ( .A(n64), .Z(n123) );
  BUF_X4 U65 ( .A(A[14]), .Z(n238) );
  CLKBUF_X1 U66 ( .A(n205), .Z(n180) );
  CLKBUF_X1 U67 ( .A(n137), .Z(n68) );
  CLKBUF_X1 U68 ( .A(n137), .Z(n69) );
  CLKBUF_X1 U69 ( .A(minus_A[20]), .Z(n136) );
  CLKBUF_X1 U70 ( .A(minus_A[12]), .Z(n120) );
  CLKBUF_X1 U71 ( .A(minus_A[21]), .Z(n138) );
  BUF_X2 U72 ( .A(A[9]), .Z(n229) );
  BUF_X2 U73 ( .A(A[9]), .Z(n230) );
  CLKBUF_X1 U74 ( .A(minus_A[22]), .Z(n139) );
  CLKBUF_X1 U75 ( .A(minus_A[22]), .Z(n140) );
  BUF_X1 U76 ( .A(minus_A[26]), .Z(n148) );
  BUF_X1 U77 ( .A(A[4]), .Z(n73) );
  BUF_X1 U78 ( .A(A[4]), .Z(n74) );
  BUF_X1 U79 ( .A(A[4]), .Z(n75) );
  BUF_X1 U80 ( .A(A[4]), .Z(n76) );
  BUF_X1 U81 ( .A(A[4]), .Z(n77) );
  BUF_X1 U82 ( .A(A[4]), .Z(n78) );
  BUF_X1 U83 ( .A(A[4]), .Z(n79) );
  BUF_X1 U84 ( .A(A[4]), .Z(n80) );
  BUF_X1 U85 ( .A(n73), .Z(n81) );
  BUF_X1 U86 ( .A(n73), .Z(n82) );
  BUF_X1 U87 ( .A(n73), .Z(n83) );
  BUF_X1 U88 ( .A(n73), .Z(n84) );
  BUF_X1 U89 ( .A(n73), .Z(n85) );
  BUF_X1 U90 ( .A(n73), .Z(n86) );
  BUF_X1 U91 ( .A(n74), .Z(n87) );
  BUF_X1 U92 ( .A(n74), .Z(n88) );
  BUF_X1 U93 ( .A(n74), .Z(n89) );
  BUF_X1 U94 ( .A(n74), .Z(n90) );
  BUF_X1 U95 ( .A(minus_A[24]), .Z(n143) );
  CLKBUF_X3 U96 ( .A(minus_A[10]), .Z(n118) );
  BUF_X2 U97 ( .A(minus_A[15]), .Z(n128) );
  BUF_X1 U98 ( .A(minus_A[17]), .Z(n132) );
  BUF_X1 U99 ( .A(minus_A[17]), .Z(n131) );
  CLKBUF_X1 U100 ( .A(minus_A[23]), .Z(n141) );
  BUF_X4 U101 ( .A(minus_A[23]), .Z(n142) );
  CLKBUF_X1 U102 ( .A(n116), .Z(n91) );
  CLKBUF_X1 U103 ( .A(n121), .Z(n92) );
  BUF_X1 U104 ( .A(minus_A[12]), .Z(n121) );
  BUF_X2 U105 ( .A(minus_A[31]), .Z(n160) );
  CLKBUF_X1 U106 ( .A(n162), .Z(n211) );
  BUF_X2 U107 ( .A(n162), .Z(n206) );
  BUF_X1 U108 ( .A(n328), .Z(n295) );
  BUF_X1 U109 ( .A(minus_A_63), .Z(n163) );
  BUF_X4 U110 ( .A(A[8]), .Z(n228) );
  BUF_X2 U111 ( .A(n206), .Z(n187) );
  BUF_X2 U112 ( .A(minus_A[25]), .Z(n146) );
  BUF_X2 U113 ( .A(n207), .Z(n183) );
  BUF_X4 U114 ( .A(n66), .Z(n149) );
  BUF_X1 U115 ( .A(minus_A_63), .Z(n162) );
  BUF_X2 U116 ( .A(minus_A[30]), .Z(n158) );
  BUF_X2 U117 ( .A(minus_A[30]), .Z(n157) );
  BUF_X2 U118 ( .A(n206), .Z(n189) );
  BUF_X1 U119 ( .A(minus_A[19]), .Z(n134) );
  CLKBUF_X1 U120 ( .A(n119), .Z(n93) );
  BUF_X1 U121 ( .A(n163), .Z(n207) );
  BUF_X1 U122 ( .A(n162), .Z(n208) );
  BUF_X2 U123 ( .A(minus_A[31]), .Z(n161) );
  BUF_X2 U124 ( .A(minus_A[27]), .Z(n94) );
  BUF_X2 U125 ( .A(minus_A[29]), .Z(n155) );
  CLKBUF_X1 U126 ( .A(n327), .Z(n303) );
  CLKBUF_X1 U127 ( .A(n327), .Z(n304) );
  CLKBUF_X1 U128 ( .A(n328), .Z(n299) );
  BUF_X1 U129 ( .A(A[27]), .Z(n270) );
  BUF_X1 U130 ( .A(A[28]), .Z(n273) );
  CLKBUF_X1 U131 ( .A(n210), .Z(n184) );
  CLKBUF_X1 U132 ( .A(n160), .Z(n159) );
  BUF_X2 U133 ( .A(n209), .Z(n173) );
  BUF_X2 U134 ( .A(n206), .Z(n188) );
  CLKBUF_X1 U135 ( .A(n211), .Z(n164) );
  CLKBUF_X1 U136 ( .A(n209), .Z(n172) );
  CLKBUF_X1 U137 ( .A(n163), .Z(n205) );
  CLKBUF_X1 U138 ( .A(n163), .Z(n210) );
  BUF_X2 U139 ( .A(minus_A[3]), .Z(n105) );
  BUF_X2 U140 ( .A(minus_A[6]), .Z(n111) );
  BUF_X2 U141 ( .A(minus_A[3]), .Z(n106) );
  BUF_X2 U142 ( .A(minus_A[25]), .Z(n147) );
  BUF_X2 U143 ( .A(minus_A[3]), .Z(n107) );
  CLKBUF_X1 U144 ( .A(n326), .Z(n307) );
  CLKBUF_X1 U145 ( .A(n326), .Z(n308) );
  CLKBUF_X1 U146 ( .A(n326), .Z(n306) );
  CLKBUF_X1 U147 ( .A(n326), .Z(n309) );
  CLKBUF_X1 U148 ( .A(n326), .Z(n311) );
  CLKBUF_X1 U149 ( .A(n331), .Z(n281) );
  CLKBUF_X1 U150 ( .A(n331), .Z(n280) );
  CLKBUF_X1 U151 ( .A(n333), .Z(n328) );
  CLKBUF_X1 U152 ( .A(n332), .Z(n329) );
  CLKBUF_X1 U153 ( .A(n333), .Z(n327) );
  CLKBUF_X1 U154 ( .A(n332), .Z(n330) );
  CLKBUF_X1 U155 ( .A(n334), .Z(n325) );
  BUF_X4 U156 ( .A(A[20]), .Z(n252) );
  BUF_X1 U157 ( .A(A[6]), .Z(n224) );
  BUF_X1 U158 ( .A(n207), .Z(n196) );
  BUF_X1 U159 ( .A(n208), .Z(n175) );
  BUF_X1 U160 ( .A(n208), .Z(n176) );
  BUF_X1 U161 ( .A(n208), .Z(n177) );
  BUF_X1 U162 ( .A(n208), .Z(n174) );
  BUF_X1 U163 ( .A(n208), .Z(n178) );
  CLKBUF_X1 U164 ( .A(n206), .Z(n191) );
  CLKBUF_X1 U165 ( .A(n206), .Z(n186) );
  CLKBUF_X1 U166 ( .A(n206), .Z(n190) );
  BUF_X1 U167 ( .A(n210), .Z(n192) );
  BUF_X1 U168 ( .A(n210), .Z(n181) );
  BUF_X1 U169 ( .A(n205), .Z(n166) );
  BUF_X1 U170 ( .A(n205), .Z(n168) );
  BUF_X1 U171 ( .A(n208), .Z(n179) );
  BUF_X1 U172 ( .A(n210), .Z(n171) );
  BUF_X1 U173 ( .A(n205), .Z(n167) );
  BUF_X1 U174 ( .A(n205), .Z(n169) );
  BUF_X1 U175 ( .A(n205), .Z(n170) );
  BUF_X1 U176 ( .A(n211), .Z(n165) );
  BUF_X1 U177 ( .A(n205), .Z(n182) );
  BUF_X1 U178 ( .A(n210), .Z(n194) );
  BUF_X1 U179 ( .A(n204), .Z(n198) );
  BUF_X1 U180 ( .A(n205), .Z(n193) );
  BUF_X1 U181 ( .A(n210), .Z(n185) );
  BUF_X1 U182 ( .A(n210), .Z(n195) );
  BUF_X1 U183 ( .A(n210), .Z(n197) );
  BUF_X1 U184 ( .A(n204), .Z(n199) );
  BUF_X1 U185 ( .A(n204), .Z(n200) );
  BUF_X1 U186 ( .A(n204), .Z(n201) );
  BUF_X1 U187 ( .A(n204), .Z(n202) );
  BUF_X1 U188 ( .A(n204), .Z(n203) );
  CLKBUF_X1 U189 ( .A(n162), .Z(n204) );
  BUF_X1 U190 ( .A(minus_A[29]), .Z(n154) );
  BUF_X1 U191 ( .A(n64), .Z(n122) );
  CLKBUF_X1 U192 ( .A(n94), .Z(n150) );
  CLKBUF_X1 U193 ( .A(minus_A[15]), .Z(n127) );
  BUF_X1 U194 ( .A(minus_A[28]), .Z(n151) );
  BUF_X1 U195 ( .A(minus_A[16]), .Z(n129) );
  CLKBUF_X1 U196 ( .A(minus_A[28]), .Z(n152) );
  BUF_X1 U197 ( .A(minus_A[24]), .Z(n144) );
  CLKBUF_X1 U198 ( .A(minus_A[29]), .Z(n156) );
  BUF_X1 U199 ( .A(minus_A[24]), .Z(n145) );
  BUF_X1 U200 ( .A(n327), .Z(n302) );
  BUF_X1 U201 ( .A(n327), .Z(n305) );
  BUF_X1 U202 ( .A(n324), .Z(n322) );
  BUF_X1 U203 ( .A(n329), .Z(n291) );
  BUF_X1 U204 ( .A(n328), .Z(n297) );
  BUF_X1 U205 ( .A(n329), .Z(n293) );
  BUF_X1 U206 ( .A(n327), .Z(n300) );
  BUF_X1 U207 ( .A(n329), .Z(n289) );
  BUF_X1 U208 ( .A(n329), .Z(n288) );
  BUF_X1 U209 ( .A(n328), .Z(n298) );
  BUF_X1 U210 ( .A(n331), .Z(n279) );
  BUF_X1 U211 ( .A(n328), .Z(n296) );
  BUF_X1 U212 ( .A(n328), .Z(n294) );
  BUF_X1 U213 ( .A(n324), .Z(n323) );
  BUF_X1 U214 ( .A(n324), .Z(n321) );
  BUF_X1 U215 ( .A(n325), .Z(n316) );
  BUF_X1 U216 ( .A(n324), .Z(n319) );
  BUF_X1 U217 ( .A(n329), .Z(n292) );
  BUF_X1 U218 ( .A(n329), .Z(n290) );
  BUF_X1 U219 ( .A(n330), .Z(n285) );
  BUF_X1 U220 ( .A(n330), .Z(n287) );
  BUF_X1 U221 ( .A(n330), .Z(n286) );
  BUF_X1 U222 ( .A(n330), .Z(n284) );
  BUF_X1 U223 ( .A(n327), .Z(n301) );
  BUF_X1 U224 ( .A(n324), .Z(n318) );
  BUF_X1 U225 ( .A(n325), .Z(n315) );
  BUF_X1 U226 ( .A(n325), .Z(n313) );
  BUF_X1 U227 ( .A(n325), .Z(n314) );
  BUF_X1 U228 ( .A(n325), .Z(n312) );
  BUF_X1 U229 ( .A(n330), .Z(n283) );
  BUF_X1 U230 ( .A(n330), .Z(n282) );
  BUF_X1 U231 ( .A(n324), .Z(n320) );
  BUF_X1 U232 ( .A(n325), .Z(n317) );
  BUF_X1 U233 ( .A(minus_A[2]), .Z(n102) );
  CLKBUF_X1 U234 ( .A(minus_A[2]), .Z(n103) );
  BUF_X2 U235 ( .A(minus_A[2]), .Z(n104) );
  BUF_X1 U236 ( .A(n95), .Z(n97) );
  BUF_X1 U237 ( .A(n333), .Z(n326) );
  BUF_X1 U238 ( .A(n332), .Z(n331) );
  BUF_X4 U239 ( .A(A[12]), .Z(n235) );
  BUF_X4 U240 ( .A(A[16]), .Z(n242) );
  BUF_X4 U241 ( .A(A[24]), .Z(n262) );
  BUF_X1 U242 ( .A(A[10]), .Z(n231) );
  BUF_X2 U243 ( .A(A[17]), .Z(n244) );
  BUF_X1 U244 ( .A(A[7]), .Z(n226) );
  BUF_X1 U245 ( .A(A[15]), .Z(n240) );
  BUF_X1 U246 ( .A(A[19]), .Z(n250) );
  BUF_X2 U247 ( .A(A[15]), .Z(n239) );
  BUF_X2 U248 ( .A(A[18]), .Z(n247) );
  BUF_X1 U249 ( .A(A[7]), .Z(n227) );
  BUF_X1 U250 ( .A(A[11]), .Z(n234) );
  BUF_X1 U251 ( .A(A[15]), .Z(n241) );
  BUF_X1 U252 ( .A(A[13]), .Z(n237) );
  BUF_X1 U253 ( .A(A[17]), .Z(n246) );
  BUF_X1 U254 ( .A(A[5]), .Z(n222) );
  BUF_X2 U255 ( .A(A[22]), .Z(n257) );
  BUF_X1 U256 ( .A(A[16]), .Z(n243) );
  BUF_X1 U257 ( .A(A[20]), .Z(n253) );
  BUF_X2 U258 ( .A(A[1]), .Z(n216) );
  BUF_X1 U259 ( .A(A[22]), .Z(n258) );
  BUF_X1 U260 ( .A(A[26]), .Z(n268) );
  BUF_X4 U261 ( .A(A[28]), .Z(n272) );
  BUF_X1 U262 ( .A(A[21]), .Z(n255) );
  BUF_X1 U263 ( .A(A[25]), .Z(n265) );
  BUF_X1 U264 ( .A(A[21]), .Z(n256) );
  BUF_X1 U265 ( .A(A[29]), .Z(n276) );
  BUF_X1 U266 ( .A(A[25]), .Z(n266) );
  BUF_X4 U267 ( .A(A[26]), .Z(n267) );
  BUF_X4 U268 ( .A(A[30]), .Z(n277) );
  BUF_X1 U269 ( .A(A[23]), .Z(n260) );
  BUF_X1 U270 ( .A(A[27]), .Z(n271) );
  BUF_X1 U271 ( .A(A[23]), .Z(n261) );
  BUF_X1 U272 ( .A(A[24]), .Z(n263) );
  BUF_X1 U273 ( .A(n67), .Z(n95) );
  BUF_X1 U274 ( .A(A[31]), .Z(n333) );
  BUF_X1 U275 ( .A(A[31]), .Z(n332) );
  BUF_X1 U276 ( .A(A[31]), .Z(n334) );
  BUF_X1 U277 ( .A(minus_A[1]), .Z(n99) );
  BUF_X1 U278 ( .A(minus_A[1]), .Z(n100) );
  BUF_X4 U279 ( .A(A[2]), .Z(n96) );
  BUF_X1 U280 ( .A(A[1]), .Z(n98) );
  BUF_X1 U281 ( .A(A[1]), .Z(n217) );
  BUF_X1 U282 ( .A(A[1]), .Z(n215) );
  BUF_X1 U283 ( .A(minus_A[0]), .Z(n212) );
endmodule

