
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity address_conversion_M8_N4_N_bit64_F3_DW01_add_2 is

   port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (4 downto 0);  CO : out std_logic);

end address_conversion_M8_N4_N_bit64_F3_DW01_add_2;

architecture SYN_rpl of address_conversion_M8_N4_N_bit64_F3_DW01_add_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, n4, n5, n6, n10, n11, n12, n_1005 : 
      std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           n_1005, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1 : INV_X1 port map( A => A(2), ZN => n12);
   U2 : OAI21_X1 port map( B1 => A(2), B2 => n10, A => B(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => A(1), B2 => B(1), A => n11, ZN => n4);
   U4 : INV_X1 port map( A => n6, ZN => n11);
   U5 : OAI211_X1 port map( C1 => A(1), C2 => B(1), A => A(0), B => B(0), ZN =>
                           n6);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n12, A => n5, ZN => carry_3_port);
   U7 : INV_X1 port map( A => n4, ZN => n10);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity address_conversion_M8_N4_N_bit64_F3_DW01_add_1 is

   port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (4 downto 0);  CO : out std_logic);

end address_conversion_M8_N4_N_bit64_F3_DW01_add_1;

architecture SYN_rpl of address_conversion_M8_N4_N_bit64_F3_DW01_add_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, n4, n5, n6, n10, n11, n12, n_1011 : 
      std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           n_1011, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1 : INV_X1 port map( A => n6, ZN => n11);
   U2 : INV_X1 port map( A => A(2), ZN => n12);
   U3 : OAI21_X1 port map( B1 => A(2), B2 => n10, A => B(2), ZN => n5);
   U4 : AOI21_X1 port map( B1 => A(1), B2 => B(1), A => n11, ZN => n4);
   U5 : OAI211_X1 port map( C1 => A(1), C2 => B(1), A => A(0), B => B(0), ZN =>
                           n6);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n12, A => n5, ZN => carry_3_port);
   U7 : INV_X1 port map( A => n4, ZN => n10);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity address_conversion_M8_N4_N_bit64_F3_DW01_add_0 is

   port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (4 downto 0);  CO : out std_logic);

end address_conversion_M8_N4_N_bit64_F3_DW01_add_0;

architecture SYN_rpl of address_conversion_M8_N4_N_bit64_F3_DW01_add_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, n4, n5, n6, n10, n11, n12, n_1017 : 
      std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           n_1017, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1 : AOI21_X1 port map( B1 => A(1), B2 => B(1), A => n11, ZN => n4);
   U2 : INV_X1 port map( A => n6, ZN => n11);
   U3 : OAI211_X1 port map( C1 => A(1), C2 => B(1), A => A(0), B => B(0), ZN =>
                           n6);
   U4 : OAI21_X1 port map( B1 => n4, B2 => n12, A => n5, ZN => carry_3_port);
   U5 : OAI21_X1 port map( B1 => A(2), B2 => n10, A => B(2), ZN => n5);
   U6 : INV_X1 port map( A => n4, ZN => n10);
   U7 : INV_X1 port map( A => A(2), ZN => n12);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity address_conversion_M8_N4_N_bit64_F3_DW01_addsub_2 is

   port( A, B : in std_logic_vector (4 downto 0);  CI, ADD_SUB : in std_logic; 
         SUM : out std_logic_vector (4 downto 0);  CO : out std_logic);

end address_conversion_M8_N4_N_bit64_F3_DW01_addsub_2;

architecture SYN_rpl of address_conversion_M8_N4_N_bit64_F3_DW01_addsub_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, carry_1_port, B_AS_4_port, 
      B_AS_3_port, B_AS_2_port, B_AS_1_port, B_AS_0_port, n_1020 : std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B_AS_4_port, CI => carry_4_port, CO 
                           => n_1020, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B_AS_3_port, CI => carry_3_port, CO 
                           => carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B_AS_2_port, CI => carry_2_port, CO 
                           => carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B_AS_1_port, CI => carry_1_port, CO 
                           => carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B_AS_0_port, CI => ADD_SUB, CO => 
                           carry_1_port, S => SUM(0));
   U1 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_AS_4_port);
   U2 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_AS_3_port);
   U3 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_AS_2_port);
   U4 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_AS_1_port);
   U5 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_AS_0_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity address_conversion_M8_N4_N_bit64_F3_DW01_addsub_1 is

   port( A, B : in std_logic_vector (4 downto 0);  CI, ADD_SUB : in std_logic; 
         SUM : out std_logic_vector (4 downto 0);  CO : out std_logic);

end address_conversion_M8_N4_N_bit64_F3_DW01_addsub_1;

architecture SYN_rpl of address_conversion_M8_N4_N_bit64_F3_DW01_addsub_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, carry_1_port, B_AS_4_port, 
      B_AS_3_port, B_AS_2_port, B_AS_1_port, B_AS_0_port, n_1023 : std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B_AS_4_port, CI => carry_4_port, CO 
                           => n_1023, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B_AS_3_port, CI => carry_3_port, CO 
                           => carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B_AS_2_port, CI => carry_2_port, CO 
                           => carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B_AS_1_port, CI => carry_1_port, CO 
                           => carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B_AS_0_port, CI => ADD_SUB, CO => 
                           carry_1_port, S => SUM(0));
   U1 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_AS_4_port);
   U2 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_AS_3_port);
   U3 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_AS_2_port);
   U4 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_AS_1_port);
   U5 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_AS_0_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity address_conversion_M8_N4_N_bit64_F3_DW01_addsub_0 is

   port( A, B : in std_logic_vector (4 downto 0);  CI, ADD_SUB : in std_logic; 
         SUM : out std_logic_vector (4 downto 0);  CO : out std_logic);

end address_conversion_M8_N4_N_bit64_F3_DW01_addsub_0;

architecture SYN_rpl of address_conversion_M8_N4_N_bit64_F3_DW01_addsub_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, carry_1_port, B_AS_4_port, 
      B_AS_3_port, B_AS_2_port, B_AS_1_port, B_AS_0_port, n_1026 : std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B_AS_4_port, CI => carry_4_port, CO 
                           => n_1026, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B_AS_3_port, CI => carry_3_port, CO 
                           => carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B_AS_2_port, CI => carry_2_port, CO 
                           => carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B_AS_1_port, CI => carry_1_port, CO 
                           => carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B_AS_0_port, CI => ADD_SUB, CO => 
                           carry_1_port, S => SUM(0));
   U1 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_AS_4_port);
   U2 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_AS_3_port);
   U3 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_AS_2_port);
   U4 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_AS_1_port);
   U5 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_AS_0_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity MUX21_generic_N5 is

   port( A, B : in std_logic_vector (4 downto 0);  sel : in std_logic;  Y : out
         std_logic_vector (4 downto 0));

end MUX21_generic_N5;

architecture SYN_BEHAVIORAL of MUX21_generic_N5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8, n9, n10, n11, n22 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n11, ZN => Y(0));
   U2 : AOI22_X1 port map( A1 => A(0), A2 => sel, B1 => B(0), B2 => n22, ZN => 
                           n11);
   U3 : INV_X1 port map( A => n9, ZN => Y(2));
   U4 : AOI22_X1 port map( A1 => A(2), A2 => sel, B1 => B(2), B2 => n22, ZN => 
                           n9);
   U5 : INV_X1 port map( A => n10, ZN => Y(1));
   U6 : AOI22_X1 port map( A1 => A(1), A2 => sel, B1 => B(1), B2 => n22, ZN => 
                           n10);
   U7 : INV_X1 port map( A => n8, ZN => Y(3));
   U8 : AOI22_X1 port map( A1 => A(3), A2 => sel, B1 => B(3), B2 => n22, ZN => 
                           n8);
   U9 : INV_X1 port map( A => sel, ZN => n22);
   U10 : INV_X1 port map( A => n7, ZN => Y(4));
   U11 : AOI22_X1 port map( A1 => sel, A2 => A(4), B1 => B(4), B2 => n22, ZN =>
                           n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_3 is

   port( A : in std_logic_vector (31 downto 0);  INC_DEC : in std_logic;  SUM :
         out std_logic_vector (31 downto 0));

end windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_3;

architecture SYN_cla of windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_3 
   is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n36, n37, n38, n39
      , n40, n41, n42, n43, n46, n47, n48, n49, n50, n51, n52, n53, n55, n56, 
      n59, n60, n61, n62, n65, n66, n68, n69, n70, n71, n72, n74, n75, n76, n77
      , n78, n79, n80, n81, n82, n83, n84, n85, n86, n88, n90, n92, n93, n94, 
      n95, n96, n98, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109
      , n110, n111, n112, n114, n116, n118, n119, n120, n121, n122, n124, n125,
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n138, 
      n139, n140, n143, n145, n146, n147, n149, n150, n151, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n174, n175, n176, n177, n179, n182, n184, 
      n185, n186, n188, n190, n191, n192, n193, n195, n196, n198, n199, n200, 
      n201, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269 : std_logic;

begin
   
   U183 : XOR2_X1 port map( A => INC_DEC, B => A(31), Z => n6);
   U225 : NAND3_X1 port map( A1 => n83, A2 => n84, A3 => n85, ZN => n75);
   U227 : NAND3_X1 port map( A1 => n109, A2 => n110, A3 => n111, ZN => n101);
   U230 : NAND3_X1 port map( A1 => n134, A2 => n135, A3 => n136, ZN => n126);
   U244 : NAND3_X1 port map( A1 => n46, A2 => n65, A3 => n50, ZN => n157);
   U1 : INV_X1 port map( A => n19, ZN => n226);
   U2 : BUF_X1 port map( A => n221, Z => n216);
   U3 : BUF_X1 port map( A => n221, Z => n215);
   U4 : BUF_X1 port map( A => n221, Z => n217);
   U5 : BUF_X1 port map( A => n221, Z => n218);
   U6 : BUF_X1 port map( A => n221, Z => n220);
   U7 : BUF_X1 port map( A => n221, Z => n219);
   U8 : NAND2_X1 port map( A1 => n154, A2 => n155, ZN => n150);
   U9 : NOR2_X1 port map( A1 => n156, A2 => n157, ZN => n155);
   U10 : AOI21_X1 port map( B1 => n158, B2 => n159, A => n160, ZN => n154);
   U11 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n156);
   U12 : OAI21_X1 port map( B1 => n227, B2 => n165, A => n1, ZN => n19);
   U13 : INV_X1 port map( A => n39, ZN => n227);
   U14 : OAI21_X1 port map( B1 => n226, B2 => n167, A => n2, ZN => n186);
   U15 : INV_X1 port map( A => INC_DEC, ZN => n221);
   U16 : OAI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n121);
   U17 : NOR2_X1 port map( A1 => n128, A2 => n129, ZN => n127);
   U18 : NAND2_X1 port map( A1 => n132, A2 => n133, ZN => n128);
   U19 : OAI21_X1 port map( B1 => n265, B2 => n59, A => n60, ZN => n52);
   U20 : INV_X1 port map( A => n61, ZN => n265);
   U21 : OAI21_X1 port map( B1 => n100, B2 => n101, A => n102, ZN => n95);
   U22 : NOR2_X1 port map( A1 => n103, A2 => n104, ZN => n102);
   U23 : NAND2_X1 port map( A1 => n107, A2 => n108, ZN => n103);
   U24 : OAI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n70);
   U25 : NOR2_X1 port map( A1 => n77, A2 => n78, ZN => n76);
   U26 : NAND2_X1 port map( A1 => n81, A2 => n82, ZN => n77);
   U27 : AOI21_X1 port map( B1 => n52, B2 => n53, A => n269, ZN => n51);
   U28 : INV_X1 port map( A => n55, ZN => n269);
   U29 : AOI21_X1 port map( B1 => n83, B2 => n88, A => n241, ZN => n86);
   U30 : INV_X1 port map( A => n80, ZN => n241);
   U31 : NAND4_X1 port map( A1 => n192, A2 => n193, A3 => n17, A4 => n21, ZN =>
                           n167);
   U32 : NAND4_X1 port map( A1 => n40, A2 => n36, A3 => n26, A4 => n29, ZN => 
                           n165);
   U33 : NOR2_X1 port map( A1 => n165, A2 => n166, ZN => n159);
   U34 : NOR2_X1 port map( A1 => n167, A2 => n168, ZN => n158);
   U35 : NAND4_X1 port map( A1 => n169, A2 => n170, A3 => n171, A4 => n172, ZN 
                           => n168);
   U36 : NAND4_X1 port map( A1 => n161, A2 => n162, A3 => n163, A4 => n164, ZN 
                           => n160);
   U37 : NAND2_X1 port map( A1 => n74, A2 => n82, ZN => n93);
   U38 : NAND2_X1 port map( A1 => n92, A2 => n81, ZN => n88);
   U39 : NAND2_X1 port map( A1 => n85, A2 => n93, ZN => n92);
   U40 : NAND2_X1 port map( A1 => n121, A2 => n122, ZN => n100);
   U41 : NAND2_X1 port map( A1 => n150, A2 => n151, ZN => n125);
   U42 : NAND2_X1 port map( A1 => n95, A2 => n96, ZN => n74);
   U43 : AND2_X1 port map( A1 => n68, A2 => n69, ZN => n59);
   U44 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => n68);
   U45 : AND4_X1 port map( A1 => n28, A2 => n24, A3 => n33, A4 => n38, ZN => n1
                           );
   U46 : AND4_X1 port map( A1 => n190, A2 => n16, A3 => n20, A4 => n191, ZN => 
                           n2);
   U47 : OAI21_X1 port map( B1 => n225, B2 => n256, A => n163, ZN => n177);
   U48 : INV_X1 port map( A => n170, ZN => n256);
   U49 : INV_X1 port map( A => n182, ZN => n225);
   U50 : OAI21_X1 port map( B1 => n31, B2 => n232, A => n33, ZN => n27);
   U51 : OAI21_X1 port map( B1 => n262, B2 => n226, A => n20, ZN => n14);
   U52 : INV_X1 port map( A => n21, ZN => n262);
   U53 : AOI21_X1 port map( B1 => n109, B2 => n114, A => n246, ZN => n112);
   U54 : INV_X1 port map( A => n106, ZN => n246);
   U55 : OAI21_X1 port map( B1 => n224, B2 => n250, A => n131, ZN => n140);
   U56 : INV_X1 port map( A => n134, ZN => n250);
   U57 : INV_X1 port map( A => n143, ZN => n224);
   U58 : OAI21_X1 port map( B1 => n222, B2 => n237, A => n46, ZN => n43);
   U59 : INV_X1 port map( A => n47, ZN => n237);
   U60 : INV_X1 port map( A => n48, ZN => n222);
   U61 : NAND2_X1 port map( A1 => n229, A2 => n166, ZN => n39);
   U62 : INV_X1 port map( A => n157, ZN => n229);
   U63 : NAND2_X1 port map( A1 => n125, A2 => n133, ZN => n147);
   U64 : NAND2_X1 port map( A1 => n100, A2 => n108, ZN => n119);
   U65 : NAND2_X1 port map( A1 => n201, A2 => n16, ZN => n199);
   U66 : NAND2_X1 port map( A1 => n14, A2 => n17, ZN => n201);
   U67 : NAND2_X1 port map( A1 => n185, A2 => n164, ZN => n182);
   U68 : NAND2_X1 port map( A1 => n186, A2 => n169, ZN => n185);
   U69 : NAND2_X1 port map( A1 => n146, A2 => n132, ZN => n143);
   U70 : NAND2_X1 port map( A1 => n136, A2 => n147, ZN => n146);
   U71 : NAND2_X1 port map( A1 => n118, A2 => n107, ZN => n114);
   U72 : NAND2_X1 port map( A1 => n111, A2 => n119, ZN => n118);
   U73 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => n23);
   U74 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => n25);
   U75 : NAND2_X1 port map( A1 => n162, A2 => n176, ZN => n175);
   U76 : NAND2_X1 port map( A1 => n171, A2 => n177, ZN => n176);
   U77 : INV_X1 port map( A => n36, ZN => n232);
   U78 : NAND2_X1 port map( A1 => n191, A2 => n198, ZN => n195);
   U79 : NAND2_X1 port map( A1 => n199, A2 => n193, ZN => n198);
   U80 : NAND2_X1 port map( A1 => n105, A2 => n106, ZN => n104);
   U81 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => n78);
   U82 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => n129);
   U83 : INV_X1 port map( A => n33, ZN => n234);
   U84 : AND2_X1 port map( A1 => n37, A2 => n38, ZN => n31);
   U85 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => n37);
   U86 : XNOR2_X1 port map( A => n51, B => n6, ZN => SUM(31));
   U87 : XNOR2_X1 port map( A => n86, B => n4, ZN => SUM(27));
   U88 : AND2_X1 port map( A1 => n79, A2 => n84, ZN => n4);
   U89 : NAND4_X1 port map( A1 => A(0), A2 => n66, A3 => n47, A4 => n49, ZN => 
                           n166);
   U90 : NAND2_X1 port map( A1 => INC_DEC, A2 => A(8), ZN => n20);
   U91 : NAND2_X1 port map( A1 => A(5), A2 => INC_DEC, ZN => n33);
   U92 : NAND2_X1 port map( A1 => A(10), A2 => INC_DEC, ZN => n191);
   U93 : NAND2_X1 port map( A1 => A(9), A2 => INC_DEC, ZN => n16);
   U94 : NAND2_X1 port map( A1 => A(6), A2 => INC_DEC, ZN => n24);
   U95 : XNOR2_X1 port map( A => n52, B => n56, ZN => SUM(30));
   U96 : NAND2_X1 port map( A1 => n55, A2 => n53, ZN => n56);
   U97 : NAND2_X1 port map( A1 => A(4), A2 => INC_DEC, ZN => n38);
   U98 : NAND2_X1 port map( A1 => n219, A2 => n263, ZN => n21);
   U99 : INV_X1 port map( A => A(8), ZN => n263);
   U100 : NAND2_X1 port map( A1 => A(12), A2 => INC_DEC, ZN => n164);
   U101 : NAND2_X1 port map( A1 => n220, A2 => n261, ZN => n17);
   U102 : INV_X1 port map( A => A(9), ZN => n261);
   U103 : NAND2_X1 port map( A1 => n220, A2 => n260, ZN => n193);
   U104 : INV_X1 port map( A => A(10), ZN => n260);
   U105 : NAND2_X1 port map( A1 => n220, A2 => n255, ZN => n171);
   U106 : INV_X1 port map( A => A(14), ZN => n255);
   U107 : NAND2_X1 port map( A1 => n220, A2 => n258, ZN => n169);
   U108 : INV_X1 port map( A => A(12), ZN => n258);
   U109 : NAND2_X1 port map( A1 => n220, A2 => n235, ZN => n40);
   U110 : INV_X1 port map( A => A(4), ZN => n235);
   U111 : NAND2_X1 port map( A1 => n219, A2 => n238, ZN => n47);
   U112 : INV_X1 port map( A => A(2), ZN => n238);
   U113 : NAND2_X1 port map( A1 => n219, A2 => n231, ZN => n26);
   U114 : INV_X1 port map( A => A(6), ZN => n231);
   U115 : NAND2_X1 port map( A1 => n219, A2 => n228, ZN => n66);
   U116 : INV_X1 port map( A => A(1), ZN => n228);
   U117 : NAND2_X1 port map( A1 => n219, A2 => n264, ZN => n29);
   U118 : INV_X1 port map( A => A(7), ZN => n264);
   U119 : NAND2_X1 port map( A1 => n218, A2 => n254, ZN => n172);
   U120 : INV_X1 port map( A => A(15), ZN => n254);
   U121 : NAND2_X1 port map( A1 => n218, A2 => n236, ZN => n49);
   U122 : INV_X1 port map( A => A(3), ZN => n236);
   U123 : NAND2_X1 port map( A1 => n218, A2 => n233, ZN => n36);
   U124 : INV_X1 port map( A => A(5), ZN => n233);
   U125 : NAND2_X1 port map( A1 => n218, A2 => n259, ZN => n192);
   U126 : INV_X1 port map( A => A(11), ZN => n259);
   U127 : NAND2_X1 port map( A1 => A(7), A2 => INC_DEC, ZN => n28);
   U128 : NAND2_X1 port map( A1 => A(11), A2 => INC_DEC, ZN => n190);
   U129 : NAND2_X1 port map( A1 => n218, A2 => n257, ZN => n170);
   U130 : INV_X1 port map( A => A(13), ZN => n257);
   U131 : OAI21_X1 port map( B1 => n230, B2 => n223, A => n65, ZN => n48);
   U132 : INV_X1 port map( A => A(0), ZN => n230);
   U133 : INV_X1 port map( A => n66, ZN => n223);
   U134 : XNOR2_X1 port map( A => n62, B => n48, ZN => SUM(2));
   U135 : NAND2_X1 port map( A1 => n47, A2 => n46, ZN => n62);
   U136 : XNOR2_X1 port map( A => n42, B => n43, ZN => SUM(3));
   U137 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => n42);
   U138 : XNOR2_X1 port map( A => n41, B => n39, ZN => SUM(4));
   U139 : NAND2_X1 port map( A1 => n38, A2 => n40, ZN => n41);
   U140 : XNOR2_X1 port map( A => n31, B => n34, ZN => SUM(5));
   U141 : NOR2_X1 port map( A1 => n234, A2 => n232, ZN => n34);
   U142 : XNOR2_X1 port map( A => n30, B => n27, ZN => SUM(6));
   U143 : NAND2_X1 port map( A1 => n26, A2 => n24, ZN => n30);
   U144 : XNOR2_X1 port map( A => n22, B => n23, ZN => SUM(7));
   U145 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => n22);
   U146 : XNOR2_X1 port map( A => n18, B => n19, ZN => SUM(8));
   U147 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => n18);
   U148 : XNOR2_X1 port map( A => n14, B => n15, ZN => SUM(9));
   U149 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => n15);
   U150 : XNOR2_X1 port map( A => n188, B => n186, ZN => SUM(12));
   U151 : NAND2_X1 port map( A1 => n164, A2 => n169, ZN => n188);
   U152 : XNOR2_X1 port map( A => n153, B => n150, ZN => SUM(16));
   U153 : NAND2_X1 port map( A1 => n133, A2 => n151, ZN => n153);
   U154 : XNOR2_X1 port map( A => n149, B => n147, ZN => SUM(17));
   U155 : NAND2_X1 port map( A1 => n132, A2 => n136, ZN => n149);
   U156 : XNOR2_X1 port map( A => n139, B => n140, ZN => SUM(19));
   U157 : NAND2_X1 port map( A1 => n130, A2 => n135, ZN => n139);
   U158 : XNOR2_X1 port map( A => n124, B => n121, ZN => SUM(20));
   U159 : NAND2_X1 port map( A1 => n108, A2 => n122, ZN => n124);
   U160 : XNOR2_X1 port map( A => n120, B => n119, ZN => SUM(21));
   U161 : NAND2_X1 port map( A1 => n107, A2 => n111, ZN => n120);
   U162 : XNOR2_X1 port map( A => n112, B => n5, ZN => SUM(23));
   U163 : AND2_X1 port map( A1 => n105, A2 => n110, ZN => n5);
   U164 : XNOR2_X1 port map( A => A(0), B => n138, ZN => SUM(1));
   U165 : NAND2_X1 port map( A1 => n66, A2 => n65, ZN => n138);
   U166 : XNOR2_X1 port map( A => n174, B => n175, ZN => SUM(15));
   U167 : NAND2_X1 port map( A1 => n161, A2 => n172, ZN => n174);
   U168 : XNOR2_X1 port map( A => n195, B => n196, ZN => SUM(11));
   U169 : NAND2_X1 port map( A1 => n190, A2 => n192, ZN => n196);
   U170 : XNOR2_X1 port map( A => n114, B => n116, ZN => SUM(22));
   U171 : NAND2_X1 port map( A1 => n109, A2 => n106, ZN => n116);
   U172 : XNOR2_X1 port map( A => n95, B => n98, ZN => SUM(24));
   U173 : NAND2_X1 port map( A1 => n82, A2 => n96, ZN => n98);
   U174 : XNOR2_X1 port map( A => n70, B => n72, ZN => SUM(28));
   U175 : NAND2_X1 port map( A1 => n69, A2 => n71, ZN => n72);
   U176 : NAND2_X1 port map( A1 => A(22), A2 => INC_DEC, ZN => n106);
   U177 : NAND2_X1 port map( A1 => A(26), A2 => INC_DEC, ZN => n80);
   U178 : NAND2_X1 port map( A1 => A(16), A2 => INC_DEC, ZN => n133);
   U179 : NAND2_X1 port map( A1 => A(20), A2 => INC_DEC, ZN => n108);
   U180 : NAND2_X1 port map( A1 => A(24), A2 => INC_DEC, ZN => n82);
   U181 : NAND2_X1 port map( A1 => A(13), A2 => INC_DEC, ZN => n163);
   U182 : NAND2_X1 port map( A1 => A(18), A2 => INC_DEC, ZN => n131);
   U184 : NAND2_X1 port map( A1 => A(17), A2 => INC_DEC, ZN => n132);
   U185 : NAND2_X1 port map( A1 => A(21), A2 => INC_DEC, ZN => n107);
   U186 : NAND2_X1 port map( A1 => A(25), A2 => INC_DEC, ZN => n81);
   U187 : NAND2_X1 port map( A1 => A(14), A2 => INC_DEC, ZN => n162);
   U188 : NAND2_X1 port map( A1 => A(1), A2 => INC_DEC, ZN => n65);
   U189 : NAND2_X1 port map( A1 => A(2), A2 => INC_DEC, ZN => n46);
   U190 : NAND2_X1 port map( A1 => n217, A2 => n245, ZN => n109);
   U191 : INV_X1 port map( A => A(22), ZN => n245);
   U192 : NAND2_X1 port map( A1 => n217, A2 => n240, ZN => n83);
   U193 : INV_X1 port map( A => A(26), ZN => n240);
   U194 : NAND2_X1 port map( A1 => n216, A2 => n268, ZN => n53);
   U195 : INV_X1 port map( A => A(30), ZN => n268);
   U196 : NAND2_X1 port map( A1 => n216, A2 => n253, ZN => n151);
   U197 : INV_X1 port map( A => A(16), ZN => n253);
   U198 : NAND2_X1 port map( A1 => n217, A2 => n248, ZN => n122);
   U199 : INV_X1 port map( A => A(20), ZN => n248);
   U200 : NAND2_X1 port map( A1 => n217, A2 => n243, ZN => n96);
   U201 : INV_X1 port map( A => A(24), ZN => n243);
   U202 : NAND2_X1 port map( A1 => n217, A2 => n239, ZN => n71);
   U203 : INV_X1 port map( A => A(28), ZN => n239);
   U204 : NAND2_X1 port map( A1 => A(30), A2 => INC_DEC, ZN => n55);
   U205 : NAND2_X1 port map( A1 => A(19), A2 => INC_DEC, ZN => n130);
   U206 : NAND2_X1 port map( A1 => A(15), A2 => INC_DEC, ZN => n161);
   U207 : NAND2_X1 port map( A1 => A(3), A2 => INC_DEC, ZN => n50);
   U208 : NAND2_X1 port map( A1 => A(29), A2 => INC_DEC, ZN => n60);
   U209 : NAND2_X1 port map( A1 => A(28), A2 => INC_DEC, ZN => n69);
   U210 : NAND2_X1 port map( A1 => A(27), A2 => INC_DEC, ZN => n79);
   U211 : NAND2_X1 port map( A1 => A(23), A2 => INC_DEC, ZN => n105);
   U212 : NAND2_X1 port map( A1 => n215, A2 => n249, ZN => n135);
   U213 : INV_X1 port map( A => A(19), ZN => n249);
   U214 : NAND2_X1 port map( A1 => n216, A2 => n266, ZN => n61);
   U215 : INV_X1 port map( A => A(29), ZN => n266);
   U216 : NAND2_X1 port map( A1 => n216, A2 => n267, ZN => n84);
   U217 : INV_X1 port map( A => A(27), ZN => n267);
   U218 : NAND2_X1 port map( A1 => n216, A2 => n244, ZN => n110);
   U219 : INV_X1 port map( A => A(23), ZN => n244);
   U220 : XNOR2_X1 port map( A => n179, B => n177, ZN => SUM(14));
   U221 : NAND2_X1 port map( A1 => n162, A2 => n171, ZN => n179);
   U222 : NAND2_X1 port map( A1 => n215, A2 => n252, ZN => n136);
   U223 : INV_X1 port map( A => A(17), ZN => n252);
   U224 : NAND2_X1 port map( A1 => n215, A2 => n251, ZN => n134);
   U226 : INV_X1 port map( A => A(18), ZN => n251);
   U228 : NAND2_X1 port map( A1 => n215, A2 => n247, ZN => n111);
   U229 : INV_X1 port map( A => A(21), ZN => n247);
   U231 : NAND2_X1 port map( A1 => n215, A2 => n242, ZN => n85);
   U232 : INV_X1 port map( A => A(25), ZN => n242);
   U233 : XNOR2_X1 port map( A => n94, B => n93, ZN => SUM(25));
   U234 : NAND2_X1 port map( A1 => n81, A2 => n85, ZN => n94);
   U235 : XNOR2_X1 port map( A => n200, B => n199, ZN => SUM(10));
   U236 : NAND2_X1 port map( A1 => n191, A2 => n193, ZN => n200);
   U237 : XNOR2_X1 port map( A => n184, B => n182, ZN => SUM(13));
   U238 : NAND2_X1 port map( A1 => n163, A2 => n170, ZN => n184);
   U239 : XNOR2_X1 port map( A => n145, B => n143, ZN => SUM(18));
   U240 : NAND2_X1 port map( A1 => n131, A2 => n134, ZN => n145);
   U241 : XNOR2_X1 port map( A => n88, B => n90, ZN => SUM(26));
   U242 : NAND2_X1 port map( A1 => n83, A2 => n80, ZN => n90);
   U243 : XNOR2_X1 port map( A => n59, B => n3, ZN => SUM(29));
   U245 : AND2_X1 port map( A1 => n60, A2 => n61, ZN => n3);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_2 is

   port( A : in std_logic_vector (31 downto 0);  INC_DEC : in std_logic;  SUM :
         out std_logic_vector (31 downto 0));

end windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_2;

architecture SYN_cla of windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_2 
   is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, 
      n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, 
      n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, 
      n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, 
      n357, n358, n359, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, SUM_0_port, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n360, n361 : 
      std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port, SUM_0_port );
   
   U128 : XOR2_X1 port map( A => n241, B => INC_DEC, Z => n247);
   U129 : XOR2_X1 port map( A => n249, B => n227, Z => SUM_8_port);
   U130 : XOR2_X1 port map( A => n239, B => INC_DEC, Z => n249);
   U131 : XOR2_X1 port map( A => n250, B => n251, Z => SUM_7_port);
   U132 : XOR2_X1 port map( A => INC_DEC, B => A(7), Z => n251);
   U133 : XOR2_X1 port map( A => n255, B => n252, Z => SUM_6_port);
   U134 : XOR2_X1 port map( A => n256, B => n258, Z => SUM_5_port);
   U135 : XOR2_X1 port map( A => n261, B => n262, Z => SUM_4_port);
   U136 : XOR2_X1 port map( A => INC_DEC, B => A(4), Z => n262);
   U137 : XOR2_X1 port map( A => n263, B => n264, Z => SUM_3_port);
   U138 : XOR2_X1 port map( A => INC_DEC, B => A(3), Z => n264);
   U139 : XOR2_X1 port map( A => n268, B => n269, Z => SUM_31_port);
   U140 : XOR2_X1 port map( A => INC_DEC, B => A(31), Z => n269);
   U141 : XOR2_X1 port map( A => INC_DEC, B => A(30), Z => n272);
   U142 : XOR2_X1 port map( A => n274, B => n265, Z => SUM_2_port);
   U143 : XOR2_X1 port map( A => n222, B => n276, Z => SUM_29_port);
   U144 : XOR2_X1 port map( A => INC_DEC, B => A(29), Z => n276);
   U145 : XOR2_X1 port map( A => n278, B => n280, Z => SUM_28_port);
   U146 : XOR2_X1 port map( A => INC_DEC, B => A(28), Z => n280);
   U147 : XOR2_X1 port map( A => n287, B => n288, Z => SUM_27_port);
   U148 : XOR2_X1 port map( A => n217, B => A(27), Z => n288);
   U149 : XOR2_X1 port map( A => n286, B => n295, Z => SUM_24_port);
   U150 : XOR2_X1 port map( A => INC_DEC, B => A(24), Z => n295);
   U151 : XOR2_X1 port map( A => n302, B => n303, Z => SUM_23_port);
   U152 : XOR2_X1 port map( A => A(23), B => n219, Z => n302);
   U153 : XOR2_X1 port map( A => n304, B => n306, Z => SUM_22_port);
   U154 : XOR2_X1 port map( A => n309, B => n307, Z => SUM_21_port);
   U155 : XOR2_X1 port map( A => A(20), B => n219, Z => n310);
   U156 : XOR2_X1 port map( A => A(0), B => n316, Z => SUM_1_port);
   U157 : XOR2_X1 port map( A => INC_DEC, B => A(1), Z => n316);
   U158 : XOR2_X1 port map( A => INC_DEC, B => A(19), Z => n318);
   U159 : XOR2_X1 port map( A => n319, B => n321, Z => SUM_18_port);
   U160 : XOR2_X1 port map( A => n217, B => A(18), Z => n321);
   U161 : XOR2_X1 port map( A => n217, B => A(17), Z => n324);
   U162 : XOR2_X1 port map( A => n313, B => n325, Z => SUM_16_port);
   U163 : XOR2_X1 port map( A => n217, B => A(16), Z => n325);
   U164 : XOR2_X1 port map( A => n336, B => n337, Z => SUM_15_port);
   U165 : XOR2_X1 port map( A => n217, B => A(15), Z => n337);
   U166 : XOR2_X1 port map( A => n217, B => A(14), Z => n340);
   U167 : XOR2_X1 port map( A => n217, B => A(13), Z => n343);
   U168 : XOR2_X1 port map( A => n344, B => n346, Z => SUM_12_port);
   U169 : XOR2_X1 port map( A => n217, B => A(12), Z => n346);
   U170 : XOR2_X1 port map( A => n349, B => n350, Z => SUM_11_port);
   U171 : XOR2_X1 port map( A => n246, B => INC_DEC, Z => n349);
   U172 : XOR2_X1 port map( A => n353, B => n352, Z => SUM_10_port);
   U173 : NAND3_X1 port map( A1 => n333, A2 => n267, A3 => n358, ZN => n261);
   U174 : XOR2_X1 port map( A => n245, B => INC_DEC, Z => n353);
   U1 : INV_X1 port map( A => INC_DEC, ZN => n219);
   U2 : OAI21_X1 port map( B1 => n227, B2 => n347, A => n329, ZN => n344);
   U3 : NOR2_X1 port map( A1 => n330, A2 => n217, ZN => n347);
   U4 : INV_X1 port map( A => n356, ZN => n227);
   U5 : NOR4_X1 port map( A1 => n246, A2 => n245, A3 => n241, A4 => n239, ZN =>
                           n330);
   U6 : NOR4_X1 port map( A1 => n332, A2 => n242, A3 => n244, A4 => n360, ZN =>
                           n331);
   U7 : NAND4_X1 port map( A1 => n245, A2 => n246, A3 => n239, A4 => n241, ZN 
                           => n348);
   U8 : OAI21_X1 port map( B1 => n332, B2 => n230, A => n326, ZN => n356);
   U9 : AOI21_X1 port map( B1 => n235, B2 => n256, A => n231, ZN => n252);
   U10 : INV_X1 port map( A => n257, ZN => n235);
   U11 : AOI21_X1 port map( B1 => n304, B2 => n232, A => n233, ZN => n303);
   U12 : INV_X1 port map( A => n305, ZN => n232);
   U13 : OAI21_X1 port map( B1 => n289, B2 => n290, A => n282, ZN => n287);
   U14 : NAND4_X1 port map( A1 => SUM_0_port, A2 => n242, A3 => n244, A4 => 
                           n360, ZN => n335);
   U15 : INV_X1 port map( A => n261, ZN => n230);
   U16 : INV_X1 port map( A => n297, ZN => n233);
   U17 : INV_X1 port map( A => n259, ZN => n231);
   U18 : INV_X1 port map( A => n339, ZN => n225);
   U19 : INV_X1 port map( A => n282, ZN => n234);
   U20 : OAI22_X1 port map( A1 => n227, A2 => n239, B1 => n355, B2 => n219, ZN 
                           => n248);
   U21 : NOR2_X1 port map( A1 => A(8), A2 => n356, ZN => n355);
   U22 : AOI22_X1 port map( A1 => n344, A2 => A(12), B1 => n345, B2 => n218, ZN
                           => n341);
   U23 : OR2_X1 port map( A1 => A(12), A2 => n344, ZN => n345);
   U24 : AOI22_X1 port map( A1 => n313, A2 => A(16), B1 => n315, B2 => n218, ZN
                           => n322);
   U25 : INV_X1 port map( A => n299, ZN => n220);
   U26 : AOI22_X1 port map( A1 => n248, A2 => A(9), B1 => n354, B2 => n218, ZN 
                           => n352);
   U27 : OR2_X1 port map( A1 => A(9), A2 => n248, ZN => n354);
   U28 : OAI21_X1 port map( B1 => n322, B2 => n240, A => n323, ZN => n319);
   U29 : INV_X1 port map( A => A(17), ZN => n240);
   U30 : OAI21_X1 port map( B1 => A(17), B2 => n229, A => n218, ZN => n323);
   U31 : INV_X1 port map( A => n322, ZN => n229);
   U32 : AOI22_X1 port map( A1 => n222, A2 => A(29), B1 => n273, B2 => n218, ZN
                           => n271);
   U33 : OR2_X1 port map( A1 => n222, A2 => A(29), ZN => n273);
   U34 : NAND4_X1 port map( A1 => n326, A2 => n327, A3 => n328, A4 => n329, ZN 
                           => n313);
   U35 : NAND4_X1 port map( A1 => n237, A2 => A(15), A3 => n330, A4 => n331, ZN
                           => n328);
   U36 : OAI21_X1 port map( B1 => n334, B2 => n335, A => n218, ZN => n327);
   U37 : INV_X1 port map( A => n333, ZN => n237);
   U38 : OAI21_X1 port map( B1 => A(3), B2 => n275, A => n217, ZN => n358);
   U39 : OAI21_X1 port map( B1 => n311, B2 => n219, A => n312, ZN => n301);
   U40 : NAND4_X1 port map( A1 => A(16), A2 => n313, A3 => A(17), A4 => n314, 
                           ZN => n312);
   U41 : NOR4_X1 port map( A1 => A(19), A2 => A(18), A3 => A(17), A4 => n315, 
                           ZN => n311);
   U42 : AND2_X1 port map( A1 => A(18), A2 => A(19), ZN => n314);
   U43 : NOR2_X1 port map( A1 => n257, A2 => n231, ZN => n258);
   U44 : NOR2_X1 port map( A1 => n217, A2 => A(5), ZN => n257);
   U45 : OAI21_X1 port map( B1 => n221, B2 => n243, A => n284, ZN => n293);
   U46 : INV_X1 port map( A => A(24), ZN => n243);
   U47 : AOI21_X1 port map( B1 => n238, B2 => n230, A => n260, ZN => n256);
   U48 : INV_X1 port map( A => A(4), ZN => n238);
   U49 : AOI21_X1 port map( B1 => n261, B2 => A(4), A => n218, ZN => n260);
   U50 : OAI21_X1 port map( B1 => n341, B2 => n244, A => n342, ZN => n339);
   U51 : OAI21_X1 port map( B1 => A(13), B2 => n226, A => n218, ZN => n342);
   U52 : INV_X1 port map( A => n341, ZN => n226);
   U53 : AOI22_X1 port map( A1 => n218, A2 => n351, B1 => A(10), B2 => n224, ZN
                           => n350);
   U54 : NAND2_X1 port map( A1 => n352, A2 => n245, ZN => n351);
   U55 : INV_X1 port map( A => n352, ZN => n224);
   U56 : INV_X1 port map( A => A(30), ZN => n361);
   U57 : NAND4_X1 port map( A1 => n281, A2 => n282, A3 => n283, A4 => n284, ZN 
                           => n278);
   U58 : OAI21_X1 port map( B1 => n285, B2 => n217, A => A(27), ZN => n281);
   U59 : NAND2_X1 port map( A1 => A(21), A2 => n217, ZN => n298);
   U60 : NAND2_X1 port map( A1 => A(26), A2 => n217, ZN => n282);
   U61 : NAND4_X1 port map( A1 => n296, A2 => n297, A3 => n298, A4 => n299, ZN 
                           => n286);
   U62 : OAI21_X1 port map( B1 => n300, B2 => n217, A => A(23), ZN => n296);
   U63 : OAI21_X1 port map( B1 => n307, B2 => n308, A => n298, ZN => n304);
   U64 : NOR2_X1 port map( A1 => A(21), A2 => n217, ZN => n308);
   U65 : NAND2_X1 port map( A1 => A(25), A2 => n218, ZN => n283);
   U66 : NAND2_X1 port map( A1 => A(2), A2 => n217, ZN => n267);
   U67 : AOI21_X1 port map( B1 => n319, B2 => A(18), A => n228, ZN => n317);
   U68 : INV_X1 port map( A => n320, ZN => n228);
   U69 : OAI21_X1 port map( B1 => A(18), B2 => n319, A => n218, ZN => n320);
   U70 : NOR2_X1 port map( A1 => A(6), A2 => n218, ZN => n253);
   U71 : NAND2_X1 port map( A1 => A(22), A2 => n217, ZN => n297);
   U72 : NAND4_X1 port map( A1 => A(3), A2 => A(1), A3 => A(2), A4 => A(0), ZN 
                           => n333);
   U73 : OAI21_X1 port map( B1 => n225, B2 => n360, A => n338, ZN => n336);
   U74 : OAI21_X1 port map( B1 => A(14), B2 => n339, A => n217, ZN => n338);
   U75 : NAND2_X1 port map( A1 => A(5), A2 => n218, ZN => n259);
   U76 : INV_X1 port map( A => A(8), ZN => n239);
   U77 : INV_X1 port map( A => A(10), ZN => n245);
   U78 : OR4_X1 port map( A1 => A(15), A2 => A(1), A3 => A(2), A4 => A(3), ZN 
                           => n334);
   U79 : INV_X1 port map( A => A(14), ZN => n360);
   U80 : XNOR2_X1 port map( A => n225, B => n340, ZN => SUM_14_port);
   U81 : XNOR2_X1 port map( A => n341, B => n343, ZN => SUM_13_port);
   U82 : INV_X1 port map( A => A(13), ZN => n244);
   U83 : XNOR2_X1 port map( A => n290, B => n291, ZN => SUM_26_port);
   U84 : NOR2_X1 port map( A1 => n289, A2 => n234, ZN => n291);
   U85 : XNOR2_X1 port map( A => n293, B => n294, ZN => SUM_25_port);
   U86 : OAI21_X1 port map( B1 => A(25), B2 => n217, A => n283, ZN => n294);
   U87 : NOR2_X1 port map( A1 => n305, A2 => n233, ZN => n306);
   U88 : XNOR2_X1 port map( A => n317, B => n318, ZN => SUM_19_port);
   U89 : OAI21_X1 port map( B1 => n218, B2 => A(21), A => n298, ZN => n309);
   U90 : XNOR2_X1 port map( A => n247, B => n248, ZN => SUM_9_port);
   U91 : XNOR2_X1 port map( A => n322, B => n324, ZN => SUM_17_port);
   U92 : INV_X1 port map( A => A(9), ZN => n241);
   U93 : INV_X1 port map( A => A(11), ZN => n246);
   U94 : AND3_X1 port map( A1 => n259, A2 => n254, A3 => n357, ZN => n326);
   U95 : OAI21_X1 port map( B1 => A(4), B2 => A(7), A => n218, ZN => n357);
   U96 : AND2_X1 port map( A1 => n283, A2 => n292, ZN => n290);
   U97 : OAI21_X1 port map( B1 => A(25), B2 => n217, A => n293, ZN => n292);
   U98 : AND2_X1 port map( A1 => n359, A2 => n219, ZN => n332);
   U99 : NAND4_X1 port map( A1 => A(7), A2 => A(4), A3 => A(5), A4 => A(6), ZN 
                           => n359);
   U100 : INV_X1 port map( A => n277, ZN => n222);
   U101 : OAI21_X1 port map( B1 => A(28), B2 => n278, A => n223, ZN => n277);
   U102 : INV_X1 port map( A => n279, ZN => n223);
   U103 : AOI21_X1 port map( B1 => n278, B2 => A(28), A => n218, ZN => n279);
   U104 : INV_X1 port map( A => A(0), ZN => SUM_0_port);
   U105 : INV_X1 port map( A => A(12), ZN => n242);
   U106 : OR2_X1 port map( A1 => n313, A2 => A(16), ZN => n315);
   U107 : OR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n275);
   U108 : AOI22_X1 port map( A1 => A(0), A2 => A(1), B1 => n275, B2 => n218, ZN
                           => n265);
   U109 : NOR2_X1 port map( A1 => n217, A2 => A(22), ZN => n305);
   U110 : NOR2_X1 port map( A1 => n217, A2 => A(26), ZN => n289);
   U111 : OAI21_X1 port map( B1 => n265, B2 => n266, A => n267, ZN => n263);
   U112 : NOR2_X1 port map( A1 => A(2), A2 => n217, ZN => n266);
   U113 : OAI21_X1 port map( B1 => n218, B2 => A(2), A => n267, ZN => n274);
   U114 : XNOR2_X1 port map( A => n310, B => n301, ZN => SUM_20_port);
   U115 : XNOR2_X1 port map( A => n271, B => n272, ZN => SUM_30_port);
   U116 : OAI21_X1 port map( B1 => n252, B2 => n253, A => n254, ZN => n250);
   U117 : OAI21_X1 port map( B1 => n218, B2 => A(6), A => n254, ZN => n255);
   U118 : AOI22_X1 port map( A1 => n270, A2 => n219, B1 => n271, B2 => n361, ZN
                           => n268);
   U119 : OR2_X1 port map( A1 => n361, A2 => n271, ZN => n270);
   U120 : AOI21_X1 port map( B1 => n301, B2 => A(20), A => n220, ZN => n307);
   U121 : INV_X1 port map( A => n286, ZN => n221);
   U122 : OAI21_X1 port map( B1 => A(24), B2 => n286, A => n218, ZN => n284);
   U123 : AND4_X1 port map( A1 => n286, A2 => A(25), A3 => A(26), A4 => A(24), 
                           ZN => n285);
   U124 : OAI21_X1 port map( B1 => A(20), B2 => n301, A => n218, ZN => n299);
   U125 : AND4_X1 port map( A1 => n301, A2 => A(21), A3 => A(22), A4 => A(20), 
                           ZN => n300);
   U126 : NAND2_X1 port map( A1 => n218, A2 => n348, ZN => n329);
   U127 : NAND2_X1 port map( A1 => INC_DEC, A2 => A(6), ZN => n254);
   U175 : INV_X1 port map( A => n219, ZN => n217);
   U176 : INV_X1 port map( A => n219, ZN => n218);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity MUX21_generic_N64 is

   port( A, B : in std_logic_vector (63 downto 0);  sel : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_generic_N64;

architecture SYN_BEHAVIORAL of MUX21_generic_N64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n243, ZN => n221);
   U2 : INV_X1 port map( A => n243, ZN => n222);
   U3 : INV_X1 port map( A => n243, ZN => n223);
   U4 : INV_X1 port map( A => n243, ZN => n224);
   U5 : INV_X1 port map( A => n243, ZN => n225);
   U6 : BUF_X1 port map( A => n244, Z => n243);
   U7 : BUF_X1 port map( A => n245, Z => n234);
   U8 : BUF_X1 port map( A => n245, Z => n233);
   U9 : BUF_X1 port map( A => n245, Z => n232);
   U10 : BUF_X1 port map( A => n246, Z => n242);
   U11 : BUF_X1 port map( A => n245, Z => n241);
   U12 : BUF_X1 port map( A => n245, Z => n240);
   U13 : BUF_X1 port map( A => n244, Z => n239);
   U14 : BUF_X1 port map( A => n245, Z => n238);
   U15 : BUF_X1 port map( A => n244, Z => n237);
   U16 : BUF_X1 port map( A => n244, Z => n236);
   U17 : BUF_X1 port map( A => n244, Z => n235);
   U18 : BUF_X1 port map( A => n246, Z => n231);
   U19 : BUF_X1 port map( A => n246, Z => n230);
   U20 : BUF_X1 port map( A => n246, Z => n229);
   U21 : BUF_X1 port map( A => n246, Z => n228);
   U22 : BUF_X1 port map( A => n246, Z => n227);
   U23 : INV_X1 port map( A => n220, ZN => n245);
   U24 : INV_X1 port map( A => n220, ZN => n244);
   U25 : INV_X1 port map( A => n220, ZN => n246);
   U26 : BUF_X1 port map( A => sel, Z => n220);
   U27 : INV_X1 port map( A => n66, ZN => Y(63));
   U28 : AOI22_X1 port map( A1 => n226, A2 => A(63), B1 => B(63), B2 => n227, 
                           ZN => n66);
   U29 : INV_X1 port map( A => n100, ZN => Y(29));
   U30 : AOI22_X1 port map( A1 => A(29), A2 => n223, B1 => B(29), B2 => n235, 
                           ZN => n100);
   U31 : INV_X1 port map( A => n99, ZN => Y(30));
   U32 : AOI22_X1 port map( A1 => A(30), A2 => n223, B1 => B(30), B2 => n235, 
                           ZN => n99);
   U33 : INV_X1 port map( A => n98, ZN => Y(31));
   U34 : AOI22_X1 port map( A1 => A(31), A2 => n223, B1 => B(31), B2 => n235, 
                           ZN => n98);
   U35 : INV_X1 port map( A => n97, ZN => Y(32));
   U36 : AOI22_X1 port map( A1 => A(32), A2 => n223, B1 => B(32), B2 => n234, 
                           ZN => n97);
   U37 : INV_X1 port map( A => n96, ZN => Y(33));
   U38 : AOI22_X1 port map( A1 => A(33), A2 => n223, B1 => B(33), B2 => n234, 
                           ZN => n96);
   U39 : INV_X1 port map( A => n95, ZN => Y(34));
   U40 : AOI22_X1 port map( A1 => A(34), A2 => n223, B1 => B(34), B2 => n234, 
                           ZN => n95);
   U41 : INV_X1 port map( A => n94, ZN => Y(35));
   U42 : AOI22_X1 port map( A1 => A(35), A2 => n223, B1 => B(35), B2 => n234, 
                           ZN => n94);
   U43 : INV_X1 port map( A => n93, ZN => Y(36));
   U44 : AOI22_X1 port map( A1 => A(36), A2 => n224, B1 => B(36), B2 => n233, 
                           ZN => n93);
   U45 : INV_X1 port map( A => n92, ZN => Y(37));
   U46 : AOI22_X1 port map( A1 => A(37), A2 => n224, B1 => B(37), B2 => n233, 
                           ZN => n92);
   U47 : INV_X1 port map( A => n91, ZN => Y(38));
   U48 : AOI22_X1 port map( A1 => A(38), A2 => n224, B1 => B(38), B2 => n233, 
                           ZN => n91);
   U49 : INV_X1 port map( A => n90, ZN => Y(39));
   U50 : AOI22_X1 port map( A1 => A(39), A2 => n224, B1 => B(39), B2 => n233, 
                           ZN => n90);
   U51 : INV_X1 port map( A => n89, ZN => Y(40));
   U52 : AOI22_X1 port map( A1 => A(40), A2 => n224, B1 => B(40), B2 => n232, 
                           ZN => n89);
   U53 : INV_X1 port map( A => n88, ZN => Y(41));
   U54 : AOI22_X1 port map( A1 => A(41), A2 => n224, B1 => B(41), B2 => n232, 
                           ZN => n88);
   U55 : INV_X1 port map( A => n87, ZN => Y(42));
   U56 : AOI22_X1 port map( A1 => A(42), A2 => n224, B1 => B(42), B2 => n232, 
                           ZN => n87);
   U57 : INV_X1 port map( A => n86, ZN => Y(43));
   U58 : AOI22_X1 port map( A1 => A(43), A2 => n224, B1 => B(43), B2 => n232, 
                           ZN => n86);
   U59 : INV_X1 port map( A => n85, ZN => Y(44));
   U60 : AOI22_X1 port map( A1 => A(44), A2 => n224, B1 => B(44), B2 => n231, 
                           ZN => n85);
   U61 : INV_X1 port map( A => n84, ZN => Y(45));
   U62 : AOI22_X1 port map( A1 => A(45), A2 => n224, B1 => B(45), B2 => n231, 
                           ZN => n84);
   U63 : INV_X1 port map( A => n74, ZN => Y(55));
   U64 : AOI22_X1 port map( A1 => A(55), A2 => n225, B1 => B(55), B2 => n229, 
                           ZN => n74);
   U65 : INV_X1 port map( A => n73, ZN => Y(56));
   U66 : AOI22_X1 port map( A1 => A(56), A2 => n225, B1 => B(56), B2 => n228, 
                           ZN => n73);
   U67 : INV_X1 port map( A => n72, ZN => Y(57));
   U68 : AOI22_X1 port map( A1 => A(57), A2 => n225, B1 => B(57), B2 => n228, 
                           ZN => n72);
   U69 : INV_X1 port map( A => n71, ZN => Y(58));
   U70 : AOI22_X1 port map( A1 => A(58), A2 => n225, B1 => B(58), B2 => n228, 
                           ZN => n71);
   U71 : INV_X1 port map( A => n70, ZN => Y(59));
   U72 : AOI22_X1 port map( A1 => A(59), A2 => n225, B1 => B(59), B2 => n228, 
                           ZN => n70);
   U73 : INV_X1 port map( A => n129, ZN => Y(0));
   U74 : AOI22_X1 port map( A1 => A(0), A2 => n221, B1 => B(0), B2 => n242, ZN 
                           => n129);
   U75 : INV_X1 port map( A => n128, ZN => Y(1));
   U76 : AOI22_X1 port map( A1 => A(1), A2 => n221, B1 => B(1), B2 => n242, ZN 
                           => n128);
   U77 : INV_X1 port map( A => n127, ZN => Y(2));
   U78 : AOI22_X1 port map( A1 => A(2), A2 => n221, B1 => B(2), B2 => n242, ZN 
                           => n127);
   U79 : INV_X1 port map( A => n126, ZN => Y(3));
   U80 : AOI22_X1 port map( A1 => A(3), A2 => n221, B1 => B(3), B2 => n242, ZN 
                           => n126);
   U81 : INV_X1 port map( A => n125, ZN => Y(4));
   U82 : AOI22_X1 port map( A1 => A(4), A2 => n221, B1 => B(4), B2 => n241, ZN 
                           => n125);
   U83 : INV_X1 port map( A => n124, ZN => Y(5));
   U84 : AOI22_X1 port map( A1 => A(5), A2 => n221, B1 => B(5), B2 => n241, ZN 
                           => n124);
   U85 : INV_X1 port map( A => n123, ZN => Y(6));
   U86 : AOI22_X1 port map( A1 => A(6), A2 => n221, B1 => B(6), B2 => n241, ZN 
                           => n123);
   U87 : INV_X1 port map( A => n122, ZN => Y(7));
   U88 : AOI22_X1 port map( A1 => A(7), A2 => n221, B1 => B(7), B2 => n241, ZN 
                           => n122);
   U89 : INV_X1 port map( A => n121, ZN => Y(8));
   U90 : AOI22_X1 port map( A1 => A(8), A2 => n221, B1 => B(8), B2 => n240, ZN 
                           => n121);
   U91 : INV_X1 port map( A => n120, ZN => Y(9));
   U92 : AOI22_X1 port map( A1 => A(9), A2 => n221, B1 => B(9), B2 => n240, ZN 
                           => n120);
   U93 : INV_X1 port map( A => n119, ZN => Y(10));
   U94 : AOI22_X1 port map( A1 => A(10), A2 => n221, B1 => B(10), B2 => n240, 
                           ZN => n119);
   U95 : INV_X1 port map( A => n118, ZN => Y(11));
   U96 : AOI22_X1 port map( A1 => A(11), A2 => n221, B1 => B(11), B2 => n240, 
                           ZN => n118);
   U97 : INV_X1 port map( A => n117, ZN => Y(12));
   U98 : AOI22_X1 port map( A1 => A(12), A2 => n222, B1 => B(12), B2 => n239, 
                           ZN => n117);
   U99 : INV_X1 port map( A => n116, ZN => Y(13));
   U100 : AOI22_X1 port map( A1 => A(13), A2 => n222, B1 => B(13), B2 => n239, 
                           ZN => n116);
   U101 : INV_X1 port map( A => n115, ZN => Y(14));
   U102 : AOI22_X1 port map( A1 => A(14), A2 => n222, B1 => B(14), B2 => n239, 
                           ZN => n115);
   U103 : INV_X1 port map( A => n114, ZN => Y(15));
   U104 : AOI22_X1 port map( A1 => A(15), A2 => n222, B1 => B(15), B2 => n239, 
                           ZN => n114);
   U105 : INV_X1 port map( A => n113, ZN => Y(16));
   U106 : AOI22_X1 port map( A1 => A(16), A2 => n222, B1 => B(16), B2 => n238, 
                           ZN => n113);
   U107 : INV_X1 port map( A => n112, ZN => Y(17));
   U108 : AOI22_X1 port map( A1 => A(17), A2 => n222, B1 => B(17), B2 => n238, 
                           ZN => n112);
   U109 : INV_X1 port map( A => n111, ZN => Y(18));
   U110 : AOI22_X1 port map( A1 => A(18), A2 => n222, B1 => B(18), B2 => n238, 
                           ZN => n111);
   U111 : INV_X1 port map( A => n110, ZN => Y(19));
   U112 : AOI22_X1 port map( A1 => A(19), A2 => n222, B1 => B(19), B2 => n238, 
                           ZN => n110);
   U113 : INV_X1 port map( A => n109, ZN => Y(20));
   U114 : AOI22_X1 port map( A1 => A(20), A2 => n222, B1 => B(20), B2 => n237, 
                           ZN => n109);
   U115 : INV_X1 port map( A => n108, ZN => Y(21));
   U116 : AOI22_X1 port map( A1 => A(21), A2 => n222, B1 => B(21), B2 => n237, 
                           ZN => n108);
   U117 : INV_X1 port map( A => n107, ZN => Y(22));
   U118 : AOI22_X1 port map( A1 => A(22), A2 => n222, B1 => B(22), B2 => n237, 
                           ZN => n107);
   U119 : INV_X1 port map( A => n106, ZN => Y(23));
   U120 : AOI22_X1 port map( A1 => A(23), A2 => n222, B1 => B(23), B2 => n237, 
                           ZN => n106);
   U121 : INV_X1 port map( A => n105, ZN => Y(24));
   U122 : AOI22_X1 port map( A1 => A(24), A2 => n223, B1 => B(24), B2 => n236, 
                           ZN => n105);
   U123 : INV_X1 port map( A => n104, ZN => Y(25));
   U124 : AOI22_X1 port map( A1 => A(25), A2 => n223, B1 => B(25), B2 => n236, 
                           ZN => n104);
   U125 : INV_X1 port map( A => n103, ZN => Y(26));
   U126 : AOI22_X1 port map( A1 => A(26), A2 => n223, B1 => B(26), B2 => n236, 
                           ZN => n103);
   U127 : INV_X1 port map( A => n102, ZN => Y(27));
   U128 : AOI22_X1 port map( A1 => A(27), A2 => n223, B1 => B(27), B2 => n236, 
                           ZN => n102);
   U129 : INV_X1 port map( A => n101, ZN => Y(28));
   U130 : AOI22_X1 port map( A1 => A(28), A2 => n223, B1 => B(28), B2 => n235, 
                           ZN => n101);
   U131 : INV_X1 port map( A => n83, ZN => Y(46));
   U132 : AOI22_X1 port map( A1 => A(46), A2 => n224, B1 => B(46), B2 => n231, 
                           ZN => n83);
   U133 : INV_X1 port map( A => n82, ZN => Y(47));
   U134 : AOI22_X1 port map( A1 => A(47), A2 => n224, B1 => B(47), B2 => n231, 
                           ZN => n82);
   U135 : INV_X1 port map( A => n81, ZN => Y(48));
   U136 : AOI22_X1 port map( A1 => A(48), A2 => n225, B1 => B(48), B2 => n230, 
                           ZN => n81);
   U137 : INV_X1 port map( A => n80, ZN => Y(49));
   U138 : AOI22_X1 port map( A1 => A(49), A2 => n225, B1 => B(49), B2 => n230, 
                           ZN => n80);
   U139 : INV_X1 port map( A => n79, ZN => Y(50));
   U140 : AOI22_X1 port map( A1 => A(50), A2 => n225, B1 => B(50), B2 => n230, 
                           ZN => n79);
   U141 : INV_X1 port map( A => n78, ZN => Y(51));
   U142 : AOI22_X1 port map( A1 => A(51), A2 => n225, B1 => B(51), B2 => n230, 
                           ZN => n78);
   U143 : INV_X1 port map( A => n77, ZN => Y(52));
   U144 : AOI22_X1 port map( A1 => A(52), A2 => n225, B1 => B(52), B2 => n229, 
                           ZN => n77);
   U145 : INV_X1 port map( A => n76, ZN => Y(53));
   U146 : AOI22_X1 port map( A1 => A(53), A2 => n225, B1 => B(53), B2 => n229, 
                           ZN => n76);
   U147 : INV_X1 port map( A => n75, ZN => Y(54));
   U148 : AOI22_X1 port map( A1 => A(54), A2 => n225, B1 => B(54), B2 => n229, 
                           ZN => n75);
   U149 : INV_X1 port map( A => n69, ZN => Y(60));
   U150 : AOI22_X1 port map( A1 => A(60), A2 => n226, B1 => B(60), B2 => n227, 
                           ZN => n69);
   U151 : INV_X1 port map( A => n68, ZN => Y(61));
   U152 : AOI22_X1 port map( A1 => A(61), A2 => n226, B1 => B(61), B2 => n227, 
                           ZN => n68);
   U153 : INV_X1 port map( A => n67, ZN => Y(62));
   U154 : AOI22_X1 port map( A1 => A(62), A2 => n226, B1 => B(62), B2 => n227, 
                           ZN => n67);
   U155 : INV_X1 port map( A => n243, ZN => n226);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity address_conversion_M8_N4_N_bit64_F3 is

   port( spill_fill_count : in std_logic;  wait_count, start_write : out 
         std_logic;  clck : in std_logic;  address_input_1, address_input_3 : 
         in std_logic_vector (4 downto 0);  address_output_1, address_output_2,
         address_output_3 : out std_logic_vector (4 downto 0);  swp, cwp : in 
         std_logic_vector (4 downto 0));

end address_conversion_M8_N4_N_bit64_F3;

architecture SYN_behavioral of address_conversion_M8_N4_N_bit64_F3 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFRS_X1
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component address_conversion_M8_N4_N_bit64_F3_DW01_add_2
      port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (4 downto 0);  CO : out std_logic);
   end component;
   
   component address_conversion_M8_N4_N_bit64_F3_DW01_add_1
      port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (4 downto 0);  CO : out std_logic);
   end component;
   
   component address_conversion_M8_N4_N_bit64_F3_DW01_add_0
      port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (4 downto 0);  CO : out std_logic);
   end component;
   
   component address_conversion_M8_N4_N_bit64_F3_DW01_addsub_2
      port( A, B : in std_logic_vector (4 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (4 downto 0);  CO : out 
            std_logic);
   end component;
   
   component address_conversion_M8_N4_N_bit64_F3_DW01_addsub_1
      port( A, B : in std_logic_vector (4 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (4 downto 0);  CO : out 
            std_logic);
   end component;
   
   component address_conversion_M8_N4_N_bit64_F3_DW01_addsub_0
      port( A, B : in std_logic_vector (4 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (4 downto 0);  CO : out 
            std_logic);
   end component;
   
   component MUX21_generic_N5
      port( A, B : in std_logic_vector (4 downto 0);  sel : in std_logic;  Y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, wait_count_port, 
      address_output_2_4_port, address_output_2_3_port, address_output_2_2_port
      , address_output_2_1_port, address_output_2_0_port, N15, N16, N45, N46, 
      ADDRESS_WRITE_cpu_4_port, ADDRESS_WRITE_cpu_3_port, 
      ADDRESS_WRITE_cpu_2_port, ADDRESS_WRITE_cpu_1_port, 
      ADDRESS_WRITE_cpu_0_port, i_4_port, i_3_port, i_2_port, i_1_port, 
      i_0_port, N77, N78, N91, N92, N93, N94, N95, N97, N98, N99, U3_U1_Z_0, 
      U3_U1_Z_1, U3_U1_Z_2, U3_U1_Z_3, U3_U1_Z_4, U3_U2_Z_0, U3_U3_Z_0, 
      U3_U3_Z_1, U3_U3_Z_2, U3_U3_Z_3, U3_U3_Z_4, U3_U4_Z_0, U3_U5_Z_0, 
      U3_U5_Z_1, U3_U5_Z_2, U3_U5_Z_3, U3_U5_Z_4, n76, add_101_carry_2_port, 
      add_101_carry_3_port, add_101_carry_4_port, n2, n20, n21, n22, n23, n24, 
      n25, n27, n28, n30, n31, n33, n34, n35, n36, n1, n9, n10, n11, n12, n13, 
      n42, n43, n44, n45_port, n46_port, n47, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033
      , n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042,
      n_1043, n_1044, n_1045 : std_logic;

begin
   wait_count <= wait_count_port;
   address_output_2 <= ( address_output_2_4_port, address_output_2_3_port, 
      address_output_2_2_port, address_output_2_1_port, address_output_2_0_port
      );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   wait_s_reg : DFFR_X1 port map( D => X_Logic1_port, CK => spill_fill_count, 
                           RN => n36, Q => wait_count_port, QN => n_1028);
   ADDRESS_COUNT_reg_4_inst : DLL_X1 port map( D => N95, GN => n55, Q => 
                           address_output_2_4_port);
   ADDRESS_COUNT_reg_3_inst : DLL_X1 port map( D => N94, GN => n55, Q => 
                           address_output_2_3_port);
   ADDRESS_COUNT_reg_2_inst : DLL_X1 port map( D => N93, GN => n55, Q => 
                           address_output_2_2_port);
   ADDRESS_COUNT_reg_1_inst : DLL_X1 port map( D => N92, GN => n55, Q => 
                           address_output_2_1_port);
   ADDRESS_COUNT_reg_0_inst : DLL_X1 port map( D => N91, GN => n55, Q => 
                           address_output_2_0_port);
   start_reg : DLL_X1 port map( D => n56, GN => n76, Q => start_write);
   add_101_U1_1_1 : HA_X1 port map( A => i_1_port, B => i_0_port, CO => 
                           add_101_carry_2_port, S => N97);
   add_101_U1_1_2 : HA_X1 port map( A => i_2_port, B => add_101_carry_2_port, 
                           CO => add_101_carry_3_port, S => N98);
   add_101_U1_1_3 : HA_X1 port map( A => i_3_port, B => add_101_carry_3_port, 
                           CO => add_101_carry_4_port, S => N99);
   n1 <= '0';
   n9 <= '0';
   n10 <= '0';
   n11 <= '0';
   n12 <= '0';
   n13 <= '0';
   ADDRESS_multiplexer_write : MUX21_generic_N5 port map( A(4) => 
                           address_output_2_4_port, A(3) => 
                           address_output_2_3_port, A(2) => 
                           address_output_2_2_port, A(1) => 
                           address_output_2_1_port, A(0) => 
                           address_output_2_0_port, B(4) => 
                           ADDRESS_WRITE_cpu_4_port, B(3) => 
                           ADDRESS_WRITE_cpu_3_port, B(2) => 
                           ADDRESS_WRITE_cpu_2_port, B(1) => 
                           ADDRESS_WRITE_cpu_1_port, B(0) => 
                           ADDRESS_WRITE_cpu_0_port, sel => wait_count_port, 
                           Y(4) => address_output_3(4), Y(3) => 
                           address_output_3(3), Y(2) => address_output_3(2), 
                           Y(1) => address_output_3(1), Y(0) => 
                           address_output_3(0));
   r150 : address_conversion_M8_N4_N_bit64_F3_DW01_addsub_0 port map( A(4) => 
                           address_input_1(4), A(3) => address_input_1(3), A(2)
                           => address_input_1(2), A(1) => address_input_1(1), 
                           A(0) => address_input_1(0), B(4) => U3_U1_Z_4, B(3) 
                           => U3_U1_Z_3, B(2) => U3_U1_Z_2, B(1) => U3_U1_Z_1, 
                           B(0) => U3_U1_Z_0, CI => n1, ADD_SUB => U3_U2_Z_0, 
                           SUM(4) => address_output_1(4), SUM(3) => 
                           address_output_1(3), SUM(2) => address_output_1(2), 
                           SUM(1) => address_output_1(1), SUM(0) => 
                           address_output_1(0), CO => n_1029);
   r160 : address_conversion_M8_N4_N_bit64_F3_DW01_addsub_1 port map( A(4) => 
                           address_input_3(4), A(3) => address_input_3(3), A(2)
                           => address_input_3(2), A(1) => address_input_3(1), 
                           A(0) => address_input_3(0), B(4) => U3_U3_Z_4, B(3) 
                           => U3_U3_Z_3, B(2) => U3_U3_Z_2, B(1) => U3_U3_Z_1, 
                           B(0) => U3_U3_Z_0, CI => n9, ADD_SUB => U3_U4_Z_0, 
                           SUM(4) => ADDRESS_WRITE_cpu_4_port, SUM(3) => 
                           ADDRESS_WRITE_cpu_3_port, SUM(2) => 
                           ADDRESS_WRITE_cpu_2_port, SUM(1) => 
                           ADDRESS_WRITE_cpu_1_port, SUM(0) => 
                           ADDRESS_WRITE_cpu_0_port, CO => n_1030);
   r174 : address_conversion_M8_N4_N_bit64_F3_DW01_addsub_2 port map( A(4) => 
                           i_4_port, A(3) => i_3_port, A(2) => i_2_port, A(1) 
                           => i_1_port, A(0) => i_0_port, B(4) => U3_U5_Z_4, 
                           B(3) => U3_U5_Z_3, B(2) => U3_U5_Z_2, B(1) => 
                           U3_U5_Z_1, B(0) => U3_U5_Z_0, CI => n10, ADD_SUB => 
                           n57, SUM(4) => N95, SUM(3) => N94, SUM(2) => N93, 
                           SUM(1) => N92, SUM(0) => N91, CO => n_1031);
   add_96 : address_conversion_M8_N4_N_bit64_F3_DW01_add_0 port map( A(4) => 
                           swp(4), A(3) => swp(3), A(2) => swp(2), A(1) => 
                           swp(1), A(0) => swp(0), B(4) => i_4_port, B(3) => 
                           i_3_port, B(2) => i_2_port, B(1) => i_1_port, B(0) 
                           => i_0_port, CI => n11, SUM(4) => N78, SUM(3) => N77
                           , SUM(2) => n_1032, SUM(1) => n_1033, SUM(0) => 
                           n_1034, CO => n_1035);
   add_52 : address_conversion_M8_N4_N_bit64_F3_DW01_add_1 port map( A(4) => 
                           address_input_1(4), A(3) => address_input_1(3), A(2)
                           => address_input_1(2), A(1) => address_input_1(1), 
                           A(0) => address_input_1(0), B(4) => cwp(4), B(3) => 
                           cwp(3), B(2) => cwp(2), B(1) => cwp(1), B(0) => 
                           cwp(0), CI => n12, SUM(4) => N16, SUM(3) => N15, 
                           SUM(2) => n_1036, SUM(1) => n_1037, SUM(0) => n_1038
                           , CO => n_1039);
   add_61 : address_conversion_M8_N4_N_bit64_F3_DW01_add_2 port map( A(4) => 
                           address_input_3(4), A(3) => address_input_3(3), A(2)
                           => address_input_3(2), A(1) => address_input_3(1), 
                           A(0) => address_input_3(0), B(4) => cwp(4), B(3) => 
                           cwp(3), B(2) => cwp(2), B(1) => cwp(1), B(0) => 
                           cwp(0), CI => n13, SUM(4) => N46, SUM(3) => N45, 
                           SUM(2) => n_1040, SUM(1) => n_1041, SUM(0) => n_1042
                           , CO => n_1043);
   i_reg_4_inst : DFFRS_X1 port map( D => X_Logic0_port, CK => spill_fill_count
                           , RN => n25, SN => n27, Q => i_4_port, QN => n22);
   i_reg_2_inst : DFFRS_X1 port map( D => X_Logic0_port, CK => spill_fill_count
                           , RN => n31, SN => n33, Q => i_2_port, QN => n_1044)
                           ;
   i_reg_0_inst : DFFRS_X1 port map( D => X_Logic0_port, CK => spill_fill_count
                           , RN => n23, SN => n24, Q => i_0_port, QN => n21);
   i_reg_3_inst : DFFRS_X1 port map( D => X_Logic0_port, CK => spill_fill_count
                           , RN => n28, SN => n30, Q => i_3_port, QN => n20);
   i_reg_1_inst : DFFRS_X1 port map( D => X_Logic0_port, CK => spill_fill_count
                           , RN => n34, SN => n35, Q => i_1_port, QN => n_1045)
                           ;
   U3 : OR2_X1 port map( A1 => n55, A2 => n21, ZN => n23);
   U4 : NAND2_X1 port map( A1 => n21, A2 => n2, ZN => n24);
   U18 : OR2_X1 port map( A1 => n56, A2 => n76, ZN => n36);
   U12 : OR2_X1 port map( A1 => n55, A2 => N98, ZN => n31);
   U8 : OR2_X1 port map( A1 => n55, A2 => N99, ZN => n28);
   U15 : OR2_X1 port map( A1 => n55, A2 => N97, ZN => n34);
   U5 : OR2_X1 port map( A1 => add_101_carry_4_port, A2 => n55, ZN => n25);
   U6 : NAND2_X1 port map( A1 => add_101_carry_4_port, A2 => n2, ZN => n27);
   U13 : NAND2_X1 port map( A1 => N98, A2 => n2, ZN => n33);
   U10 : NAND2_X1 port map( A1 => N99, A2 => n2, ZN => n30);
   U16 : NAND2_X1 port map( A1 => N97, A2 => n2, ZN => n35);
   U19 : INV_X1 port map( A => n47, ZN => n59);
   U21 : INV_X1 port map( A => n2, ZN => n55);
   U22 : INV_X1 port map( A => n44, ZN => n65);
   U23 : AOI21_X1 port map( B1 => N15, B2 => N16, A => n66, ZN => n47);
   U24 : INV_X1 port map( A => n46_port, ZN => n66);
   U25 : AND3_X1 port map( A1 => N16, A2 => n46_port, A3 => N15, ZN => 
                           U3_U2_Z_0);
   U26 : NOR2_X1 port map( A1 => n42, A2 => n76, ZN => n2);
   U27 : INV_X1 port map( A => n43, ZN => n57);
   U28 : INV_X1 port map( A => n42, ZN => n56);
   U29 : OAI21_X1 port map( B1 => n64, B2 => n59, A => n46_port, ZN => 
                           U3_U1_Z_4);
   U30 : NOR2_X1 port map( A1 => n61, A2 => n59, ZN => U3_U1_Z_2);
   U31 : NOR2_X1 port map( A1 => n62, A2 => n59, ZN => U3_U1_Z_1);
   U32 : NOR2_X1 port map( A1 => n63, A2 => n59, ZN => U3_U1_Z_0);
   U33 : INV_X1 port map( A => cwp(2), ZN => n61);
   U34 : INV_X1 port map( A => cwp(4), ZN => n64);
   U35 : INV_X1 port map( A => cwp(0), ZN => n63);
   U36 : INV_X1 port map( A => cwp(3), ZN => n60);
   U37 : AOI21_X1 port map( B1 => address_input_1(3), B2 => address_input_1(2),
                           A => address_input_1(4), ZN => n46_port);
   U38 : AOI21_X1 port map( B1 => address_input_3(3), B2 => address_input_3(2),
                           A => address_input_3(4), ZN => n44);
   U39 : NAND2_X1 port map( A1 => N78, A2 => N77, ZN => n43);
   U40 : AND2_X1 port map( A1 => swp(0), A2 => n43, ZN => U3_U5_Z_0);
   U41 : AND2_X1 port map( A1 => swp(1), A2 => n43, ZN => U3_U5_Z_1);
   U42 : AND2_X1 port map( A1 => swp(2), A2 => n43, ZN => U3_U5_Z_2);
   U43 : OR2_X1 port map( A1 => n57, A2 => swp(3), ZN => U3_U5_Z_3);
   U44 : NAND2_X1 port map( A1 => n22, A2 => n20, ZN => n42);
   U45 : NAND2_X1 port map( A1 => wait_count_port, A2 => clck, ZN => n76);
   U46 : AND2_X1 port map( A1 => swp(4), A2 => n43, ZN => U3_U5_Z_4);
   U47 : INV_X1 port map( A => cwp(1), ZN => n62);
   U48 : AND3_X1 port map( A1 => N46, A2 => n44, A3 => N45, ZN => U3_U4_Z_0);
   U49 : NAND2_X1 port map( A1 => n47, A2 => n60, ZN => U3_U1_Z_3);
   U50 : AOI21_X1 port map( B1 => N45, B2 => N46, A => n65, ZN => n45_port);
   U51 : OAI21_X1 port map( B1 => n58, B2 => n64, A => n44, ZN => U3_U3_Z_4);
   U52 : NAND2_X1 port map( A1 => n45_port, A2 => n60, ZN => U3_U3_Z_3);
   U53 : NOR2_X1 port map( A1 => n58, A2 => n61, ZN => U3_U3_Z_2);
   U54 : NOR2_X1 port map( A1 => n58, A2 => n62, ZN => U3_U3_Z_1);
   U55 : INV_X1 port map( A => n45_port, ZN => n58);
   U56 : NOR2_X1 port map( A1 => n58, A2 => n63, ZN => U3_U3_Z_0);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity register_file_NBIT64_NREG32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_NBIT64_NREG32;

architecture SYN_A of register_file_NBIT64_NREG32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
      n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, 
      n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, 
      n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, 
      n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, 
      n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, 
      n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, 
      n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, 
      n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, 
      n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, 
      n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, 
      n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, 
      n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, 
      n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, 
      n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, 
      n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, 
      n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, 
      n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, 
      n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, 
      n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, 
      n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, 
      n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, 
      n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, 
      n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, 
      n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, 
      n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, 
      n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, 
      n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, 
      n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, 
      n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, 
      n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, 
      n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, 
      n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, 
      n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, 
      n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, 
      n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, 
      n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, 
      n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, 
      n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, 
      n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, 
      n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, 
      n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, 
      n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, 
      n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, 
      n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, 
      n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, 
      n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, 
      n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, 
      n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, 
      n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, 
      n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, 
      n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, 
      n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, 
      n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, 
      n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, 
      n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, 
      n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, 
      n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, 
      n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, 
      n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, 
      n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, 
      n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, 
      n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, 
      n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, 
      n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, 
      n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, 
      n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, 
      n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, 
      n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, 
      n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, 
      n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, 
      n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, 
      n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, 
      n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, 
      n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, 
      n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, 
      n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, 
      n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, 
      n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, 
      n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, 
      n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, 
      n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, 
      n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, 
      n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, 
      n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, 
      n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, 
      n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, 
      n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, 
      n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, 
      n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, 
      n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, 
      n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, 
      n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, 
      n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, 
      n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, 
      n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, 
      n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, 
      n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, 
      n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, 
      n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, 
      n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, 
      n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, 
      n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, 
      n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, 
      n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, 
      n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, 
      n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, 
      n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, 
      n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, 
      n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, 
      n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, 
      n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, 
      n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, 
      n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, 
      n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, 
      n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, 
      n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, 
      n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, 
      n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, 
      n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, 
      n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, 
      n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, 
      n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, 
      n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, 
      n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, 
      n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, 
      n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, 
      n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, 
      n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, 
      n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, 
      n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, 
      n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, 
      n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, 
      n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, 
      n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, 
      n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, 
      n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, 
      n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, 
      n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, 
      n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, 
      n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, 
      n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, 
      n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, 
      n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, 
      n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, 
      n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, 
      n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, 
      n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, 
      n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, 
      n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, 
      n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, 
      n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, 
      n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, 
      n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, 
      n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, 
      n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, 
      n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, 
      n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, 
      n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, 
      n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, 
      n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, 
      n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, 
      n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, 
      n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, 
      n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, 
      n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, 
      n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, 
      n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, 
      n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, 
      n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, 
      n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, 
      n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, 
      n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, 
      n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, 
      n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, 
      n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, 
      n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, 
      n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, 
      n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, 
      n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, 
      n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, 
      n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, 
      n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, 
      n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, 
      n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, 
      n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, 
      n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, 
      n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, 
      n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, 
      n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, 
      n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, 
      n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, 
      n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, 
      n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, 
      n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, 
      n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, 
      n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, 
      n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, 
      n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, 
      n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, 
      n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, 
      n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, 
      n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, 
      n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, 
      n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, 
      n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, 
      n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, 
      n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, 
      n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, 
      n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, 
      n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, 
      n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, 
      n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, 
      n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, 
      n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, 
      n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, 
      n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, 
      n7032, n7033, n7034, n7035, n7036, n7037, n4765, n4766, n4767, n4768, 
      n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, 
      n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, 
      n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4803, 
      n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, 
      n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, 
      n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, 
      n4834, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, 
      n4846, n4847, n4848, n4849, n4850, n4851, n4854, n4855, n4856, n4857, 
      n4858, n4859, n4860, n4861, n7106, n7107, n7108, n7109, n7110, n7111, 
      n7112, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, 
      n7124, n7125, n7126, n7127, n7128, n7129, n7132, n7133, n7134, n7135, 
      n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, 
      n7146, n7149, n7150, n7151, n7152, n7153, n7234, n7235, n7236, n7237, 
      n7238, n7239, n7240, n7241, n7242, n7243, n7246, n7247, n7248, n7249, 
      n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, 
      n7260, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, 
      n7272, n7273, n7274, n7275, n7276, n7277, n7362, n7363, n7364, n7365, 
      n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, 
      n7376, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, 
      n7388, n7389, n7390, n7391, n7392, n7393, n7396, n7397, n7398, n7399, 
      n7400, n7401, n7402, n7403, n7404, n7490, n7491, n7492, n7493, n7494, 
      n7495, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, 
      n7507, n7508, n7509, n7510, n7511, n7512, n7515, n7516, n7517, n7518, 
      n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, 
      n7529, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, 
      n7628, n7629, n7630, n7631, n7632, n7633, n7636, n7637, n7638, n7639, 
      n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, 
      n7650, n7653, n7654, n7655, n7656, n7742, n7743, n7744, n7745, n7746, 
      n7747, n7748, n7749, n7750, n7751, n7752, n7755, n7756, n7757, n7758, 
      n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, 
      n7769, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, 
      n7781, n7782, n7783, n7784, n7785, n7786, n7789, n7790, n7791, n7792, 
      n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, 
      n7803, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, 
      n7815, n7816, n7817, n7818, n7819, n7820, n7823, n7824, n7825, n7826, 
      n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, 
      n7837, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, 
      n7849, n7850, n7851, n7852, n7853, n7854, n7857, n7858, n7859, n7860, 
      n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, 
      n7871, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, 
      n7883, n7884, n7885, n7886, n7887, n7888, n7891, n7892, n7893, n7894, 
      n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, 
      n7905, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, 
      n7917, n7918, n7919, n7920, n7921, n7922, n7925, n7926, n7927, n7928, 
      n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, 
      n7939, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, 
      n7951, n7952, n7953, n7954, n7955, n7956, n7959, n7960, n7961, n7962, 
      n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, 
      n7973, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, 
      n7985, n7986, n7987, n7988, n7989, n7990, n7993, n7994, n7995, n7996, 
      n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, 
      n8007, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, 
      n8019, n8020, n8021, n8022, n8023, n8024, n8027, n8028, n8029, n8030, 
      n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, 
      n8041, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, 
      n8053, n8054, n8055, n8056, n8057, n8058, n8061, n8062, n8063, n8064, 
      n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, 
      n8075, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, 
      n8087, n8088, n8089, n8090, n8091, n8092, n8095, n8096, n8097, n8098, 
      n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, 
      n8109, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, 
      n8121, n8122, n8123, n8124, n8125, n8126, n8129, n8130, n8131, n8132, 
      n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, 
      n8143, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, 
      n8155, n8156, n8157, n8158, n8159, n8160, n8163, n8164, n8165, n8166, 
      n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, 
      n8177, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, 
      n8189, n8190, n8191, n8192, n8193, n8194, n8197, n8198, n8199, n8200, 
      n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, 
      n8211, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, 
      n8223, n8224, n8225, n8226, n8227, n8228, n8231, n8232, n8233, n8234, 
      n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, 
      n8245, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, 
      n8257, n8258, n8259, n8260, n8261, n8262, n8265, n8266, n8267, n8268, 
      n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, 
      n8279, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, 
      n8291, n8292, n8293, n8294, n8295, n8296, n8299, n8300, n8301, n8302, 
      n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, 
      n8313, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, 
      n8325, n8326, n8327, n8328, n8329, n8330, n8333, n8334, n8335, n8336, 
      n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, 
      n8347, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, 
      n8359, n8360, n8361, n8362, n8363, n8364, n8366, n8367, n8368, n8369, 
      n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, 
      n8380, n8381, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, 
      n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8400, n8401, 
      n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, 
      n8412, n8413, n8414, n8415, n8417, n8418, n8419, n8420, n8421, n8422, 
      n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, 
      n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, 
      n8444, n8445, n8446, n8447, n8448, n8449, n8451, n8452, n8453, n8454, 
      n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, 
      n8465, n8466, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, 
      n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8485, n8486, 
      n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, 
      n8497, n8498, n8499, n8500, n8502, n8503, n8504, n8505, n8506, n8507, 
      n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, 
      n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, 
      n8529, n8530, n8531, n8532, n8533, n8534, n8536, n8537, n8538, n8539, 
      n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, 
      n8550, n8551, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, 
      n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8570, n8571, 
      n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, 
      n8582, n8583, n8584, n9885, n9886, n9887, n9888, n9889, n9890, n9891, 
      n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, 
      n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, 
      n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, 
      n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, 
      n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, 
      n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, 
      n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, 
      n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, 
      n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, 
      n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, 
      n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
      n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
      n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
      n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
      n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
      n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
      n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
      n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
      n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
      n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
      n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
      n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
      n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
      n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
      n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
      n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
      n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
      n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
      n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
      n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
      n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
      n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
      n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
      n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
      n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
      n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
      n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, 
      n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, 
      n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, 
      n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, 
      n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, 
      n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, 
      n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, 
      n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, 
      n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, 
      n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, 
      n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, 
      n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
      n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, 
      n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, 
      n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, 
      n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, 
      n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, 
      n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, 
      n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
      n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
      n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, 
      n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, 
      n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, 
      n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, 
      n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, 
      n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, 
      n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, 
      n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, 
      n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, 
      n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, 
      n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, 
      n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, 
      n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, 
      n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, 
      n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, 
      n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, 
      n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, 
      n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, 
      n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, 
      n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, 
      n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, 
      n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, 
      n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, 
      n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, 
      n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, 
      n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, 
      n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, 
      n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, 
      n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, 
      n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, 
      n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, 
      n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, 
      n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, 
      n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, 
      n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, 
      n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, 
      n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, 
      n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
      n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
      n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
      n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, 
      n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, 
      n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, 
      n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, 
      n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
      n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
      n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, 
      n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
      n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
      n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
      n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
      n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, 
      n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, 
      n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, 
      n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
      n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
      n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, 
      n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
      n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
      n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
      n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, 
      n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, 
      n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, 
      n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, 
      n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
      n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
      n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, 
      n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, 
      n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, 
      n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, 
      n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, 
      n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, 
      n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, 
      n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, 
      n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, 
      n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, 
      n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, 
      n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
      n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, 
      n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, 
      n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, 
      n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, 
      n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, 
      n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, 
      n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, 
      n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
      n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
      n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, 
      n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
      n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
      n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, 
      n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, 
      n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
      n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, 
      n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
      n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, 
      n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
      n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, 
      n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, 
      n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, 
      n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
      n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, 
      n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, 
      n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, 
      n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, 
      n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, 
      n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
      n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, 
      n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, 
      n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, 
      n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, 
      n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, 
      n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, 
      n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, 
      n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, 
      n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, 
      n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, 
      n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, 
      n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, 
      n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, 
      n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, 
      n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, 
      n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, 
      n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, 
      n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, 
      n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, 
      n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, 
      n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, 
      n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, 
      n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, 
      n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, 
      n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, 
      n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
      n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
      n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, 
      n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, 
      n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, 
      n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, 
      n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, 
      n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, 
      n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
      n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, 
      n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, 
      n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, 
      n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, 
      n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, 
      n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, 
      n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, 
      n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, 
      n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, 
      n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, 
      n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, 
      n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, 
      n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, 
      n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, 
      n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, 
      n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, 
      n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, 
      n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, 
      n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, 
      n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, 
      n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, 
      n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, 
      n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, 
      n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, 
      n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, 
      n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, 
      n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, 
      n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, 
      n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, 
      n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
      n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, 
      n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, 
      n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, 
      n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, 
      n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, 
      n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, 
      n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, 
      n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, 
      n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, 
      n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, 
      n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, 
      n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, 
      n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, 
      n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, 
      n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4642, 
      n4643, n4646, n4647, n4648, n4649, n4652, n4653, n4654, n4655, n4656, 
      n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, 
      n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, 
      n4677, n4678, n4679, n4682, n4683, n4684, n4685, n7080, n7081, n7084, 
      n7085, n7088, n7089, n7092, n7093, n7096, n7097, n7100, n7101, n7104, 
      n7105, n7130, n7131, n7154, n7155, n7158, n7159, n7162, n7163, n7166, 
      n7167, n7170, n7171, n7174, n7175, n7178, n7179, n7182, n7183, n7186, 
      n7187, n7190, n7191, n7194, n7195, n7198, n7199, n7202, n7205, n7208, 
      n7211, n7214, n7217, n7220, n7223, n7226, n7229, n7232, n7245, n7278, 
      n7279, n7282, n7283, n7286, n7287, n7290, n7291, n7294, n7295, n7298, 
      n7299, n7302, n7303, n7306, n7307, n7310, n7311, n7314, n7315, n7318, 
      n7319, n7322, n7323, n8599, n8600, n8603, n8604, n8605, n8606, n8611, 
      n8612, n8613, n8614, n8617, n8618, n8619, n8620, n8621, n8622, n8623, 
      n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, 
      n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, 
      n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, 
      n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, 
      n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, 
      n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, 
      n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, 
      n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, 
      n8704, n8705, n8706, n8707, n8708, n11406, n11407, n11408, n11409, n11410
      , n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
      n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, 
      n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, 
      n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, 
      n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, 
      n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, 
      n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, 
      n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, 
      n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, 
      n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, 
      n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, 
      n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, 
      n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, 
      n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, 
      n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, 
      n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, 
      n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, 
      n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, 
      n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, 
      n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, 
      n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, 
      n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, 
      n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, 
      n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, 
      n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, 
      n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, 
      n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, 
      n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, 
      n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, 
      n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, 
      n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, 
      n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, 
      n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, 
      n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, 
      n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, 
      n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, 
      n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, 
      n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, 
      n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, 
      n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, 
      n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, 
      n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, 
      n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, 
      n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, 
      n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, 
      n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, 
      n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, 
      n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, 
      n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, 
      n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, 
      n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, 
      n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, 
      n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, 
      n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, 
      n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, 
      n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, 
      n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, 
      n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, 
      n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, 
      n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, 
      n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, 
      n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, 
      n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, 
      n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, 
      n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, 
      n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, 
      n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, 
      n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, 
      n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, 
      n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, 
      n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, 
      n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, 
      n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, 
      n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, 
      n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, 
      n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, 
      n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, 
      n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, 
      n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, 
      n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, 
      n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, 
      n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, 
      n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, 
      n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, 
      n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, 
      n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, 
      n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, 
      n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, 
      n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, 
      n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, 
      n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, 
      n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, 
      n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, 
      n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, 
      n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, 
      n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, 
      n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, 
      n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, 
      n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, 
      n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, 
      n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, 
      n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, 
      n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, 
      n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, 
      n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, 
      n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, 
      n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, 
      n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, 
      n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, 
      n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, 
      n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, 
      n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, 
      n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, 
      n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, 
      n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, 
      n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, 
      n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, 
      n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, 
      n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, 
      n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, 
      n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, 
      n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, 
      n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, 
      n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, 
      n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, 
      n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, 
      n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, 
      n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, 
      n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, 
      n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, 
      n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, 
      n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, 
      n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, 
      n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, 
      n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, 
      n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, 
      n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, 
      n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, 
      n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, 
      n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, 
      n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, 
      n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, 
      n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, 
      n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, 
      n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, 
      n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, 
      n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, 
      n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, 
      n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, 
      n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, 
      n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, 
      n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, 
      n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, 
      n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, 
      n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, 
      n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, 
      n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, 
      n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, 
      n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, 
      n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, 
      n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, 
      n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, 
      n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, 
      n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, 
      n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, 
      n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, 
      n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, 
      n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, 
      n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, 
      n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, 
      n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, 
      n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, 
      n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, 
      n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, 
      n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, 
      n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, 
      n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, 
      n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, 
      n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, 
      n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, 
      n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, 
      n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, 
      n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, 
      n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, 
      n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, 
      n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, 
      n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, 
      n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, 
      n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, 
      n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, 
      n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, 
      n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, 
      n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, 
      n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, 
      n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, 
      n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, 
      n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, 
      n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, 
      n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, 
      n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, 
      n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, 
      n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, 
      n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, 
      n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, 
      n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, 
      n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, 
      n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, 
      n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, 
      n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, 
      n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, 
      n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, 
      n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, 
      n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, 
      n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, 
      n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, 
      n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, 
      n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, 
      n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, 
      n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, 
      n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, 
      n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, 
      n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, 
      n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, 
      n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, 
      n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, 
      n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, 
      n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, 
      n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, 
      n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, 
      n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, 
      n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, 
      n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, 
      n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, 
      n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, 
      n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, 
      n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, 
      n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, 
      n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, 
      n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, 
      n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, 
      n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, 
      n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, 
      n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, 
      n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, 
      n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, 
      n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, 
      n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, 
      n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, 
      n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, 
      n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, 
      n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, 
      n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, 
      n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, 
      n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, 
      n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, 
      n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, 
      n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, 
      n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, 
      n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, 
      n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, 
      n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, 
      n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, 
      n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, 
      n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, 
      n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, 
      n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, 
      n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, 
      n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, 
      n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, 
      n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, 
      n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, 
      n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, 
      n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, 
      n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, 
      n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, 
      n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, 
      n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, 
      n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, 
      n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, 
      n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, 
      n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, 
      n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, 
      n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, 
      n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, 
      n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, 
      n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, 
      n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, 
      n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, 
      n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, 
      n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, 
      n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, 
      n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, 
      n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, 
      n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, 
      n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, 
      n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, 
      n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, 
      n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, 
      n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, 
      n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, 
      n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, 
      n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, 
      n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, 
      n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, 
      n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, 
      n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, 
      n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, 
      n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, 
      n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, 
      n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, 
      n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, 
      n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, 
      n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, 
      n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, 
      n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, 
      n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, 
      n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, 
      n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, 
      n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, 
      n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, 
      n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, 
      n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, 
      n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, 
      n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, 
      n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, 
      n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, 
      n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, 
      n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, 
      n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, 
      n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, 
      n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, 
      n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, 
      n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, 
      n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, 
      n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, 
      n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, 
      n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, 
      n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, 
      n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, 
      n14462, n14463, n14464, n14465, n14466, n_1046, n_1047, n_1048, n_1049, 
      n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, 
      n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, 
      n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, 
      n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, 
      n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, 
      n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, 
      n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, 
      n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, 
      n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, 
      n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, 
      n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, 
      n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, 
      n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, 
      n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, 
      n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, 
      n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, 
      n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, 
      n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, 
      n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, 
      n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, 
      n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, 
      n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, 
      n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, 
      n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, 
      n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, 
      n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, 
      n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, 
      n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, 
      n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, 
      n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, 
      n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, 
      n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, 
      n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, 
      n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, 
      n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, 
      n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, 
      n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, 
      n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, 
      n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, 
      n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, 
      n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, 
      n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, 
      n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, 
      n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, 
      n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, 
      n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, 
      n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, 
      n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, 
      n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, 
      n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, 
      n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, 
      n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, 
      n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, 
      n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, 
      n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, 
      n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, 
      n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, 
      n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, 
      n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, 
      n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, 
      n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, 
      n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, 
      n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, 
      n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, 
      n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, 
      n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, 
      n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, 
      n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, 
      n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, 
      n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, 
      n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, 
      n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, 
      n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, 
      n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, 
      n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, 
      n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, 
      n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, 
      n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, 
      n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, 
      n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, 
      n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, 
      n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, 
      n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, 
      n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, 
      n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, 
      n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, 
      n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, 
      n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, 
      n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, 
      n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, 
      n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, 
      n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, 
      n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, 
      n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, 
      n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, 
      n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, 
      n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, 
      n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, 
      n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, 
      n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, 
      n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, 
      n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, 
      n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, 
      n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, 
      n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, 
      n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, 
      n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, 
      n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, 
      n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, 
      n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, 
      n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, 
      n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, 
      n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, 
      n_2067, n_2068, n_2069 : std_logic;

begin
   
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n7037, CK => CLK, Q => 
                           n_1046, QN => n13392);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n7028, CK => CLK, Q => 
                           n_1047, QN => n13393);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n7027, CK => CLK, Q => 
                           n_1048, QN => n13394);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n7026, CK => CLK, Q => 
                           n_1049, QN => n13395);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n7025, CK => CLK, Q => 
                           n_1050, QN => n13396);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n7024, CK => CLK, Q => 
                           n_1051, QN => n13397);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n7023, CK => CLK, Q => 
                           n_1052, QN => n13398);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n7022, CK => CLK, Q => 
                           n_1053, QN => n13399);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n7021, CK => CLK, Q => 
                           n_1054, QN => n13400);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n7020, CK => CLK, Q => 
                           n_1055, QN => n13401);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n6938, CK => CLK, Q => 
                           n_1056, QN => n13402);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n6937, CK => CLK, Q => 
                           n_1057, QN => n13403);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n6936, CK => CLK, Q => 
                           n_1058, QN => n13404);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n6935, CK => CLK, Q => 
                           n_1059, QN => n13405);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n6934, CK => CLK, Q => 
                           n_1060, QN => n13406);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n6933, CK => CLK, Q => 
                           n_1061, QN => n13407);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n6932, CK => CLK, Q => 
                           n_1062, QN => n13408);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n6931, CK => CLK, Q => 
                           n_1063, QN => n13409);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n6930, CK => CLK, Q => 
                           n_1064, QN => n13410);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n6929, CK => CLK, Q => 
                           n_1065, QN => n13411);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n6928, CK => CLK, Q => 
                           n_1066, QN => n13412);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n6927, CK => CLK, Q => 
                           n_1067, QN => n13413);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n6926, CK => CLK, Q => 
                           n_1068, QN => n13414);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n6925, CK => CLK, Q => 
                           n_1069, QN => n13415);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n6924, CK => CLK, Q => 
                           n_1070, QN => n13416);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n6923, CK => CLK, Q => 
                           n_1071, QN => n13417);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n6922, CK => CLK, Q => 
                           n_1072, QN => n13418);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n6921, CK => CLK, Q => 
                           n_1073, QN => n13419);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n6920, CK => CLK, Q => 
                           n_1074, QN => n13420);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n6919, CK => CLK, Q => n_1075
                           , QN => n13421);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n6918, CK => CLK, Q => n_1076
                           , QN => n13422);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n6917, CK => CLK, Q => n_1077
                           , QN => n13423);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n6916, CK => CLK, Q => n_1078
                           , QN => n13424);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n6915, CK => CLK, Q => n_1079
                           , QN => n13425);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n6914, CK => CLK, Q => n_1080
                           , QN => n13426);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n6913, CK => CLK, Q => n_1081
                           , QN => n13427);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n6912, CK => CLK, Q => n_1082
                           , QN => n13428);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n6911, CK => CLK, Q => n_1083
                           , QN => n13429);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n6910, CK => CLK, Q => n_1084
                           , QN => n13430);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => n6393, CK => CLK, Q => 
                           n_1085, QN => n13435);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => n6392, CK => CLK, Q => 
                           n_1086, QN => n13436);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => n6391, CK => CLK, Q => 
                           n_1087, QN => n13437);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => n6390, CK => CLK, Q => 
                           n_1088, QN => n13438);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => n6389, CK => CLK, Q => 
                           n_1089, QN => n13439);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => n6388, CK => CLK, Q => 
                           n_1090, QN => n13440);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => n6387, CK => CLK, Q => 
                           n_1091, QN => n13441);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => n6386, CK => CLK, Q => 
                           n_1092, QN => n13442);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => n6385, CK => CLK, Q => 
                           n_1093, QN => n13443);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => n6384, CK => CLK, Q => 
                           n_1094, QN => n13444);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => n6383, CK => CLK, Q => 
                           n_1095, QN => n13445);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => n6382, CK => CLK, Q => 
                           n_1096, QN => n13446);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => n6381, CK => CLK, Q => 
                           n_1097, QN => n13447);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => n6380, CK => CLK, Q => 
                           n_1098, QN => n13448);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => n6379, CK => CLK, Q => 
                           n_1099, QN => n13449);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => n6378, CK => CLK, Q => 
                           n_1100, QN => n13450);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => n6377, CK => CLK, Q => 
                           n_1101, QN => n13451);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => n6376, CK => CLK, Q => 
                           n_1102, QN => n13452);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => n6375, CK => CLK, Q => 
                           n_1103, QN => n13453);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => n6374, CK => CLK, Q => 
                           n_1104, QN => n13454);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => n6373, CK => CLK, Q => 
                           n_1105, QN => n13455);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => n6372, CK => CLK, Q => 
                           n_1106, QN => n13456);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => n6371, CK => CLK, Q => 
                           n_1107, QN => n13457);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => n6370, CK => CLK, Q => 
                           n_1108, QN => n13458);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => n6369, CK => CLK, Q => 
                           n_1109, QN => n13459);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => n6368, CK => CLK, Q => 
                           n_1110, QN => n13460);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => n6367, CK => CLK, Q => 
                           n_1111, QN => n13461);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => n6366, CK => CLK, Q => 
                           n_1112, QN => n13462);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n6365, CK => CLK, Q => 
                           n_1113, QN => n13463);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n6364, CK => CLK, Q => 
                           n_1114, QN => n13464);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n6363, CK => CLK, Q => 
                           n_1115, QN => n13465);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n6362, CK => CLK, Q => 
                           n_1116, QN => n13466);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n6361, CK => CLK, Q => 
                           n_1117, QN => n13467);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n6360, CK => CLK, Q => 
                           n_1118, QN => n13468);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n6359, CK => CLK, Q => 
                           n_1119, QN => n13469);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n6358, CK => CLK, Q => 
                           n_1120, QN => n13470);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n6357, CK => CLK, Q => 
                           n_1121, QN => n13471);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n6356, CK => CLK, Q => 
                           n_1122, QN => n13472);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n6355, CK => CLK, Q => 
                           n_1123, QN => n13473);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n6354, CK => CLK, Q => 
                           n_1124, QN => n13474);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n6353, CK => CLK, Q => 
                           n_1125, QN => n13475);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n6352, CK => CLK, Q => 
                           n_1126, QN => n13476);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n6351, CK => CLK, Q => 
                           n_1127, QN => n13477);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n6350, CK => CLK, Q => 
                           n_1128, QN => n13478);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n6349, CK => CLK, Q => 
                           n_1129, QN => n13479);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n6348, CK => CLK, Q => 
                           n_1130, QN => n13480);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n6347, CK => CLK, Q => 
                           n_1131, QN => n13481);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n6346, CK => CLK, Q => 
                           n_1132, QN => n13482);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n6345, CK => CLK, Q => 
                           n_1133, QN => n13483);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n6344, CK => CLK, Q => 
                           n_1134, QN => n13484);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n6343, CK => CLK, Q => 
                           n_1135, QN => n13485);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n6342, CK => CLK, Q => 
                           n_1136, QN => n13486);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n6341, CK => CLK, Q => 
                           n_1137, QN => n13487);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n6340, CK => CLK, Q => 
                           n_1138, QN => n13488);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n6339, CK => CLK, Q => 
                           n_1139, QN => n13489);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n6338, CK => CLK, Q => 
                           n_1140, QN => n13490);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n6337, CK => CLK, Q => 
                           n_1141, QN => n13491);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n6336, CK => CLK, Q => 
                           n_1142, QN => n13492);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n6335, CK => CLK, Q => 
                           n_1143, QN => n13493);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n6334, CK => CLK, Q => 
                           n_1144, QN => n13494);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => n6329, CK => CLK, Q => 
                           n_1145, QN => n13499);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => n6328, CK => CLK, Q => 
                           n_1146, QN => n13500);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => n6327, CK => CLK, Q => 
                           n_1147, QN => n13501);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => n6326, CK => CLK, Q => 
                           n_1148, QN => n13502);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => n6325, CK => CLK, Q => 
                           n_1149, QN => n13503);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => n6324, CK => CLK, Q => 
                           n_1150, QN => n13504);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => n6323, CK => CLK, Q => 
                           n_1151, QN => n13505);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => n6322, CK => CLK, Q => 
                           n_1152, QN => n13506);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => n6321, CK => CLK, Q => 
                           n_1153, QN => n13507);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => n6320, CK => CLK, Q => 
                           n_1154, QN => n13508);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => n6319, CK => CLK, Q => 
                           n_1155, QN => n13509);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => n6318, CK => CLK, Q => 
                           n_1156, QN => n13510);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => n6317, CK => CLK, Q => 
                           n_1157, QN => n13511);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => n6316, CK => CLK, Q => 
                           n_1158, QN => n13512);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => n6315, CK => CLK, Q => 
                           n_1159, QN => n13513);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => n6314, CK => CLK, Q => 
                           n_1160, QN => n13514);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => n6313, CK => CLK, Q => 
                           n_1161, QN => n13515);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => n6308, CK => CLK, Q => 
                           n_1162, QN => n13516);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => n6307, CK => CLK, Q => 
                           n_1163, QN => n13517);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => n6306, CK => CLK, Q => 
                           n_1164, QN => n13518);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => n6305, CK => CLK, Q => 
                           n_1165, QN => n13519);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => n6304, CK => CLK, Q => 
                           n_1166, QN => n13520);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => n6303, CK => CLK, Q => 
                           n_1167, QN => n13521);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => n6302, CK => CLK, Q => 
                           n_1168, QN => n13522);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n6301, CK => CLK, Q => 
                           n_1169, QN => n13523);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n6300, CK => CLK, Q => 
                           n_1170, QN => n13524);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n6299, CK => CLK, Q => 
                           n_1171, QN => n13525);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n6298, CK => CLK, Q => 
                           n_1172, QN => n13526);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n6297, CK => CLK, Q => 
                           n_1173, QN => n13527);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n6296, CK => CLK, Q => 
                           n_1174, QN => n13528);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n6295, CK => CLK, Q => 
                           n_1175, QN => n13529);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n6294, CK => CLK, Q => 
                           n_1176, QN => n13530);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n6293, CK => CLK, Q => 
                           n_1177, QN => n13531);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n6292, CK => CLK, Q => 
                           n_1178, QN => n13532);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n6291, CK => CLK, Q => 
                           n_1179, QN => n13533);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n6290, CK => CLK, Q => 
                           n_1180, QN => n13534);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n6286, CK => CLK, Q => 
                           n_1181, QN => n13535);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n6273, CK => CLK, Q => 
                           n_1182, QN => n13536);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n6272, CK => CLK, Q => 
                           n_1183, QN => n13537);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n6271, CK => CLK, Q => 
                           n_1184, QN => n13538);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n6270, CK => CLK, Q => 
                           n_1185, QN => n13539);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => n6137, CK => CLK, Q => 
                           n_1186, QN => n13544);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => n6136, CK => CLK, Q => 
                           n_1187, QN => n13545);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => n6135, CK => CLK, Q => 
                           n_1188, QN => n13546);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => n6134, CK => CLK, Q => 
                           n_1189, QN => n13547);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => n6133, CK => CLK, Q => 
                           n_1190, QN => n13548);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => n6132, CK => CLK, Q => 
                           n_1191, QN => n13549);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => n6131, CK => CLK, Q => 
                           n_1192, QN => n13550);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => n6130, CK => CLK, Q => 
                           n_1193, QN => n13551);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => n6129, CK => CLK, Q => 
                           n_1194, QN => n13552);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => n6128, CK => CLK, Q => 
                           n_1195, QN => n13553);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => n6127, CK => CLK, Q => 
                           n_1196, QN => n13554);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => n6126, CK => CLK, Q => 
                           n_1197, QN => n13555);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => n6125, CK => CLK, Q => 
                           n_1198, QN => n13556);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => n6124, CK => CLK, Q => 
                           n_1199, QN => n13557);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => n6123, CK => CLK, Q => 
                           n_1200, QN => n13558);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => n6122, CK => CLK, Q => 
                           n_1201, QN => n13559);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => n6121, CK => CLK, Q => 
                           n_1202, QN => n13560);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => n6120, CK => CLK, Q => 
                           n_1203, QN => n13561);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => n6119, CK => CLK, Q => 
                           n_1204, QN => n13562);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => n6118, CK => CLK, Q => 
                           n_1205, QN => n13563);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => n6117, CK => CLK, Q => 
                           n_1206, QN => n13564);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => n6116, CK => CLK, Q => 
                           n_1207, QN => n13565);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => n6115, CK => CLK, Q => 
                           n_1208, QN => n13566);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => n6114, CK => CLK, Q => 
                           n_1209, QN => n13567);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => n6113, CK => CLK, Q => 
                           n_1210, QN => n13568);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => n6112, CK => CLK, Q => 
                           n_1211, QN => n13569);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => n6111, CK => CLK, Q => 
                           n_1212, QN => n13570);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => n6110, CK => CLK, Q => 
                           n_1213, QN => n13571);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n6109, CK => CLK, Q => 
                           n_1214, QN => n13572);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n6108, CK => CLK, Q => 
                           n_1215, QN => n13573);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n6107, CK => CLK, Q => 
                           n_1216, QN => n13574);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n6106, CK => CLK, Q => 
                           n_1217, QN => n13575);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n6105, CK => CLK, Q => 
                           n_1218, QN => n13576);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n6104, CK => CLK, Q => 
                           n_1219, QN => n13577);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n6103, CK => CLK, Q => 
                           n_1220, QN => n13578);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n6102, CK => CLK, Q => 
                           n_1221, QN => n13579);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n6101, CK => CLK, Q => 
                           n_1222, QN => n13580);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n6100, CK => CLK, Q => 
                           n_1223, QN => n13581);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n6099, CK => CLK, Q => 
                           n_1224, QN => n13582);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n6098, CK => CLK, Q => 
                           n_1225, QN => n13583);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n6097, CK => CLK, Q => 
                           n_1226, QN => n13584);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n6096, CK => CLK, Q => 
                           n_1227, QN => n13585);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n6095, CK => CLK, Q => 
                           n_1228, QN => n13586);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n6094, CK => CLK, Q => 
                           n_1229, QN => n13587);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n6093, CK => CLK, Q => 
                           n_1230, QN => n13588);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n6092, CK => CLK, Q => 
                           n_1231, QN => n13589);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n6091, CK => CLK, Q => 
                           n_1232, QN => n13590);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n6090, CK => CLK, Q => 
                           n_1233, QN => n13591);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n6089, CK => CLK, Q => 
                           n_1234, QN => n13592);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n6088, CK => CLK, Q => 
                           n_1235, QN => n13593);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n6087, CK => CLK, Q => 
                           n_1236, QN => n13594);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n6086, CK => CLK, Q => 
                           n_1237, QN => n13595);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n6085, CK => CLK, Q => 
                           n_1238, QN => n13596);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n6084, CK => CLK, Q => 
                           n_1239, QN => n13597);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n6083, CK => CLK, Q => 
                           n_1240, QN => n13598);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n6082, CK => CLK, Q => 
                           n_1241, QN => n13599);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n6081, CK => CLK, Q => 
                           n_1242, QN => n13600);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n6080, CK => CLK, Q => 
                           n_1243, QN => n13601);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n6079, CK => CLK, Q => 
                           n_1244, QN => n13602);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n6078, CK => CLK, Q => 
                           n_1245, QN => n13603);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => n6073, CK => CLK, Q => 
                           n_1246, QN => n13608);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => n6072, CK => CLK, Q => 
                           n_1247, QN => n13609);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => n6071, CK => CLK, Q => 
                           n_1248, QN => n13610);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => n6070, CK => CLK, Q => 
                           n_1249, QN => n13611);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => n6069, CK => CLK, Q => 
                           n_1250, QN => n13612);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => n6068, CK => CLK, Q => 
                           n_1251, QN => n13613);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => n6067, CK => CLK, Q => 
                           n_1252, QN => n13614);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => n6066, CK => CLK, Q => 
                           n_1253, QN => n13615);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => n6065, CK => CLK, Q => 
                           n_1254, QN => n13616);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => n6064, CK => CLK, Q => 
                           n_1255, QN => n13617);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => n6063, CK => CLK, Q => 
                           n_1256, QN => n13618);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => n6062, CK => CLK, Q => 
                           n_1257, QN => n13619);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => n6061, CK => CLK, Q => 
                           n_1258, QN => n13620);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => n6060, CK => CLK, Q => 
                           n_1259, QN => n13621);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => n6059, CK => CLK, Q => 
                           n_1260, QN => n13622);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => n6058, CK => CLK, Q => 
                           n_1261, QN => n13623);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => n6057, CK => CLK, Q => 
                           n_1262, QN => n13624);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => n6056, CK => CLK, Q => 
                           n_1263, QN => n13625);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => n6055, CK => CLK, Q => 
                           n_1264, QN => n13626);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => n6054, CK => CLK, Q => 
                           n_1265, QN => n13627);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => n6053, CK => CLK, Q => 
                           n_1266, QN => n13628);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => n6052, CK => CLK, Q => 
                           n_1267, QN => n13629);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => n6051, CK => CLK, Q => 
                           n_1268, QN => n13630);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => n6050, CK => CLK, Q => 
                           n_1269, QN => n13631);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => n6049, CK => CLK, Q => 
                           n_1270, QN => n13632);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => n6048, CK => CLK, Q => 
                           n_1271, QN => n13633);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => n6047, CK => CLK, Q => 
                           n_1272, QN => n13634);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => n6046, CK => CLK, Q => 
                           n_1273, QN => n13635);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n6045, CK => CLK, Q => 
                           n_1274, QN => n13636);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n6044, CK => CLK, Q => 
                           n_1275, QN => n13637);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n6043, CK => CLK, Q => 
                           n_1276, QN => n13638);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n6042, CK => CLK, Q => 
                           n_1277, QN => n13639);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n6041, CK => CLK, Q => 
                           n_1278, QN => n13640);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n6040, CK => CLK, Q => 
                           n_1279, QN => n13641);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n6039, CK => CLK, Q => 
                           n_1280, QN => n13642);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n6038, CK => CLK, Q => 
                           n_1281, QN => n13643);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n6037, CK => CLK, Q => 
                           n_1282, QN => n13644);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n6036, CK => CLK, Q => 
                           n_1283, QN => n13645);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n6030, CK => CLK, Q => 
                           n_1284, QN => n13646);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n6017, CK => CLK, Q => 
                           n_1285, QN => n13647);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n6016, CK => CLK, Q => 
                           n_1286, QN => n13648);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n6015, CK => CLK, Q => 
                           n_1287, QN => n13649);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n6014, CK => CLK, Q => 
                           n_1288, QN => n13650);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => n5881, CK => CLK, Q => 
                           n4682, QN => n12128);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => n5880, CK => CLK, Q => 
                           n4678, QN => n12127);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => n5879, CK => CLK, Q => 
                           n4676, QN => n12126);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => n5878, CK => CLK, Q => 
                           n4674, QN => n12125);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => n5877, CK => CLK, Q => 
                           n4672, QN => n12124);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => n5876, CK => CLK, Q => 
                           n4670, QN => n12123);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => n5875, CK => CLK, Q => 
                           n4668, QN => n12122);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => n5874, CK => CLK, Q => 
                           n4666, QN => n12121);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => n5873, CK => CLK, Q => 
                           n4664, QN => n12120);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => n5872, CK => CLK, Q => 
                           n4662, QN => n12119);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => n5871, CK => CLK, Q => 
                           n4660, QN => n12118);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => n5870, CK => CLK, Q => 
                           n4658, QN => n12117);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => n5869, CK => CLK, Q => 
                           n4656, QN => n12116);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => n5868, CK => CLK, Q => 
                           n8695, QN => n12115);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => n5867, CK => CLK, Q => 
                           n8693, QN => n12114);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => n5866, CK => CLK, Q => 
                           n8691, QN => n12113);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => n5865, CK => CLK, Q => 
                           n8689, QN => n12112);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => n5864, CK => CLK, Q => 
                           n8687, QN => n12111);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => n5863, CK => CLK, Q => 
                           n8685, QN => n12110);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => n5862, CK => CLK, Q => 
                           n8683, QN => n12109);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => n5861, CK => CLK, Q => 
                           n8681, QN => n12108);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => n5860, CK => CLK, Q => 
                           n8679, QN => n12107);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => n5859, CK => CLK, Q => 
                           n8677, QN => n12106);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => n5858, CK => CLK, Q => 
                           n8675, QN => n12105);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => n5857, CK => CLK, Q => 
                           n8673, QN => n12104);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => n5856, CK => CLK, Q => 
                           n8671, QN => n12103);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => n5855, CK => CLK, Q => 
                           n8669, QN => n12102);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => n5854, CK => CLK, Q => 
                           n8667, QN => n12101);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n5853, CK => CLK, Q => 
                           n8665, QN => n12100);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n5852, CK => CLK, Q => 
                           n8663, QN => n12099);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n5851, CK => CLK, Q => 
                           n8661, QN => n12098);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n5850, CK => CLK, Q => 
                           n8659, QN => n12097);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n5849, CK => CLK, Q => 
                           n8657, QN => n12096);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n5848, CK => CLK, Q => 
                           n8655, QN => n12095);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n5847, CK => CLK, Q => 
                           n8653, QN => n12094);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n5846, CK => CLK, Q => 
                           n8651, QN => n12093);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n5845, CK => CLK, Q => 
                           n8649, QN => n12045);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n5844, CK => CLK, Q => 
                           n8647, QN => n12044);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n5843, CK => CLK, Q => 
                           n8645, QN => n12043);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n5842, CK => CLK, Q => 
                           n8643, QN => n12042);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n5841, CK => CLK, Q => 
                           n8641, QN => n12041);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n5840, CK => CLK, Q => 
                           n8639, QN => n12040);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n5839, CK => CLK, Q => 
                           n8637, QN => n12039);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n5838, CK => CLK, Q => 
                           n8635, QN => n12038);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n5837, CK => CLK, Q => 
                           n8633, QN => n12037);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n5836, CK => CLK, Q => 
                           n8631, QN => n12036);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n5835, CK => CLK, Q => 
                           n8629, QN => n12035);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n5834, CK => CLK, Q => 
                           n8627, QN => n12034);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n5833, CK => CLK, Q => 
                           n8625, QN => n12033);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n5832, CK => CLK, Q => 
                           n8623, QN => n12032);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n5831, CK => CLK, Q => n8621
                           , QN => n12031);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n5830, CK => CLK, Q => n8619
                           , QN => n12030);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n5829, CK => CLK, Q => n8617
                           , QN => n12029);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n5828, CK => CLK, Q => n8611
                           , QN => n12028);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n5827, CK => CLK, Q => n8603
                           , QN => n12027);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n5826, CK => CLK, Q => n8599
                           , QN => n12026);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n5825, CK => CLK, Q => n4654
                           , QN => n12025);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n5824, CK => CLK, Q => n4652
                           , QN => n12024);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n5823, CK => CLK, Q => n4646
                           , QN => n12023);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n5822, CK => CLK, Q => n4642
                           , QN => n12022);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => n5817, CK => CLK, Q => 
                           n4683, QN => n11958);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => n5816, CK => CLK, Q => 
                           n4679, QN => n11957);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => n5815, CK => CLK, Q => 
                           n4677, QN => n11956);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => n5814, CK => CLK, Q => 
                           n4675, QN => n11955);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => n5813, CK => CLK, Q => 
                           n4673, QN => n11954);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => n5812, CK => CLK, Q => 
                           n4671, QN => n11953);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => n5811, CK => CLK, Q => 
                           n4669, QN => n11952);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => n5810, CK => CLK, Q => 
                           n4667, QN => n11951);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => n5809, CK => CLK, Q => 
                           n4665, QN => n11950);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => n5808, CK => CLK, Q => 
                           n4663, QN => n11949);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => n5807, CK => CLK, Q => 
                           n4661, QN => n11948);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => n5806, CK => CLK, Q => 
                           n4659, QN => n11947);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => n5805, CK => CLK, Q => 
                           n4657, QN => n11946);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n5761, CK => CLK, Q => n4655
                           , QN => n11850);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n5760, CK => CLK, Q => n4653
                           , QN => n11849);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n5759, CK => CLK, Q => n4647
                           , QN => n11848);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n5758, CK => CLK, Q => n4643
                           , QN => n11847);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => n5625, CK => CLK, Q => 
                           n4684, QN => n12092);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => n5624, CK => CLK, Q => 
                           n4502, QN => n12091);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => n5623, CK => CLK, Q => 
                           n4500, QN => n12090);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => n5622, CK => CLK, Q => 
                           n4498, QN => n12089);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => n5621, CK => CLK, Q => 
                           n4496, QN => n12088);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => n5620, CK => CLK, Q => 
                           n4494, QN => n12087);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => n5619, CK => CLK, Q => 
                           n4492, QN => n12086);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => n5618, CK => CLK, Q => 
                           n4490, QN => n12085);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => n5617, CK => CLK, Q => 
                           n4488, QN => n12084);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => n5616, CK => CLK, Q => 
                           n4486, QN => n12083);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => n5615, CK => CLK, Q => 
                           n7322, QN => n12082);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => n5614, CK => CLK, Q => 
                           n7318, QN => n12081);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => n5613, CK => CLK, Q => 
                           n7314, QN => n12080);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => n5612, CK => CLK, Q => 
                           n7310, QN => n12079);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => n5611, CK => CLK, Q => 
                           n7306, QN => n12078);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => n5610, CK => CLK, Q => 
                           n7302, QN => n12077);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => n5609, CK => CLK, Q => 
                           n7298, QN => n12076);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => n5608, CK => CLK, Q => 
                           n7294, QN => n12075);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => n5607, CK => CLK, Q => 
                           n7290, QN => n12074);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => n5606, CK => CLK, Q => 
                           n7286, QN => n12073);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => n5605, CK => CLK, Q => 
                           n7282, QN => n12072);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => n5604, CK => CLK, Q => 
                           n7278, QN => n12071);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => n5603, CK => CLK, Q => 
                           n7245, QN => n12070);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => n5602, CK => CLK, Q => 
                           n7232, QN => n12069);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => n5601, CK => CLK, Q => 
                           n7229, QN => n12068);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => n5600, CK => CLK, Q => 
                           n7226, QN => n12067);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => n5599, CK => CLK, Q => 
                           n7223, QN => n12066);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => n5598, CK => CLK, Q => 
                           n7220, QN => n12065);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n5597, CK => CLK, Q => 
                           n7217, QN => n12064);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n5596, CK => CLK, Q => 
                           n7214, QN => n12063);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n5595, CK => CLK, Q => 
                           n7211, QN => n12062);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n5594, CK => CLK, Q => 
                           n7208, QN => n12061);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n5593, CK => CLK, Q => 
                           n7205, QN => n12060);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n5592, CK => CLK, Q => 
                           n7202, QN => n12059);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n5591, CK => CLK, Q => 
                           n7198, QN => n12058);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n5590, CK => CLK, Q => 
                           n7194, QN => n12057);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n5589, CK => CLK, Q => 
                           n7190, QN => n12021);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n5588, CK => CLK, Q => 
                           n7186, QN => n12020);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n5587, CK => CLK, Q => 
                           n7182, QN => n12019);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n5586, CK => CLK, Q => 
                           n7178, QN => n12018);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n5585, CK => CLK, Q => 
                           n7174, QN => n12017);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n5584, CK => CLK, Q => 
                           n7170, QN => n12016);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n5583, CK => CLK, Q => 
                           n7166, QN => n12015);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n5582, CK => CLK, Q => 
                           n7162, QN => n12014);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n5581, CK => CLK, Q => 
                           n7158, QN => n12013);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n5580, CK => CLK, Q => 
                           n7154, QN => n12012);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n5579, CK => CLK, Q => 
                           n7130, QN => n12011);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n5578, CK => CLK, Q => 
                           n7104, QN => n12010);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n5577, CK => CLK, Q => 
                           n7100, QN => n12009);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n5576, CK => CLK, Q => 
                           n7096, QN => n12008);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n5575, CK => CLK, Q => n7092
                           , QN => n12007);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n5574, CK => CLK, Q => n7088
                           , QN => n12006);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n5573, CK => CLK, Q => n7084
                           , QN => n12005);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n5572, CK => CLK, Q => n8613
                           , QN => n12004);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n5571, CK => CLK, Q => n8605
                           , QN => n12003);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n5570, CK => CLK, Q => n7080
                           , QN => n12002);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n5569, CK => CLK, Q => n4484
                           , QN => n12001);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n5568, CK => CLK, Q => n4482
                           , QN => n12000);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n5567, CK => CLK, Q => n4648
                           , QN => n11999);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n5566, CK => CLK, Q => n4480
                           , QN => n11998);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => n5561, CK => CLK, Q => 
                           n4685, QN => n11945);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => n5560, CK => CLK, Q => 
                           n4503, QN => n11944);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => n5559, CK => CLK, Q => 
                           n4501, QN => n11943);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => n5558, CK => CLK, Q => 
                           n4499, QN => n11942);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => n5557, CK => CLK, Q => 
                           n4497, QN => n11941);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => n5556, CK => CLK, Q => 
                           n4495, QN => n11940);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => n5555, CK => CLK, Q => 
                           n4493, QN => n11939);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => n5554, CK => CLK, Q => 
                           n4491, QN => n11938);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => n5553, CK => CLK, Q => 
                           n4489, QN => n11937);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => n5552, CK => CLK, Q => 
                           n4487, QN => n11936);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n5505, CK => CLK, Q => n4485
                           , QN => n11846);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n5504, CK => CLK, Q => n4483
                           , QN => n11845);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n5503, CK => CLK, Q => n4649
                           , QN => n11844);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n5502, CK => CLK, Q => n4481
                           , QN => n11843);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => n5497, CK => CLK, Q => 
                           n_1289, QN => n13671);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => n5496, CK => CLK, Q => 
                           n_1290, QN => n13672);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => n5495, CK => CLK, Q => 
                           n_1291, QN => n13673);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => n5494, CK => CLK, Q => 
                           n_1292, QN => n13674);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => n5493, CK => CLK, Q => 
                           n_1293, QN => n13675);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => n5492, CK => CLK, Q => 
                           n_1294, QN => n13676);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => n5491, CK => CLK, Q => 
                           n_1295, QN => n13677);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => n5490, CK => CLK, Q => 
                           n_1296, QN => n13678);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => n5489, CK => CLK, Q => 
                           n_1297, QN => n13679);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => n5488, CK => CLK, Q => 
                           n_1298, QN => n13680);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => n5487, CK => CLK, Q => 
                           n_1299, QN => n13681);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => n5486, CK => CLK, Q => 
                           n_1300, QN => n13682);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => n5485, CK => CLK, Q => 
                           n_1301, QN => n13683);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => n5484, CK => CLK, Q => 
                           n_1302, QN => n13684);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => n5483, CK => CLK, Q => 
                           n_1303, QN => n13685);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => n5482, CK => CLK, Q => 
                           n_1304, QN => n13686);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => n5481, CK => CLK, Q => 
                           n_1305, QN => n13687);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => n5480, CK => CLK, Q => 
                           n_1306, QN => n13688);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => n5479, CK => CLK, Q => 
                           n_1307, QN => n13689);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => n5478, CK => CLK, Q => 
                           n_1308, QN => n13690);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => n5477, CK => CLK, Q => 
                           n_1309, QN => n13691);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => n5476, CK => CLK, Q => 
                           n_1310, QN => n13692);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => n5475, CK => CLK, Q => 
                           n_1311, QN => n13693);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => n5474, CK => CLK, Q => 
                           n_1312, QN => n13694);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => n5473, CK => CLK, Q => 
                           n_1313, QN => n13695);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => n5472, CK => CLK, Q => 
                           n_1314, QN => n13696);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => n5471, CK => CLK, Q => 
                           n_1315, QN => n13697);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => n5470, CK => CLK, Q => 
                           n_1316, QN => n13698);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n5469, CK => CLK, Q => 
                           n_1317, QN => n13699);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n5468, CK => CLK, Q => 
                           n_1318, QN => n13700);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n5467, CK => CLK, Q => 
                           n_1319, QN => n13701);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n5466, CK => CLK, Q => 
                           n_1320, QN => n13702);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n5465, CK => CLK, Q => 
                           n_1321, QN => n13703);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n5464, CK => CLK, Q => 
                           n_1322, QN => n13704);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n5463, CK => CLK, Q => 
                           n_1323, QN => n13705);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n5462, CK => CLK, Q => 
                           n_1324, QN => n13706);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n5461, CK => CLK, Q => 
                           n_1325, QN => n13707);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n5460, CK => CLK, Q => 
                           n_1326, QN => n13708);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n5459, CK => CLK, Q => 
                           n_1327, QN => n13709);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n5458, CK => CLK, Q => 
                           n_1328, QN => n13710);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n5457, CK => CLK, Q => 
                           n_1329, QN => n13711);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n5456, CK => CLK, Q => 
                           n_1330, QN => n13712);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n5455, CK => CLK, Q => 
                           n_1331, QN => n13713);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n5454, CK => CLK, Q => 
                           n_1332, QN => n13714);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n5453, CK => CLK, Q => 
                           n_1333, QN => n13715);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n5452, CK => CLK, Q => 
                           n_1334, QN => n13716);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n5451, CK => CLK, Q => 
                           n_1335, QN => n13717);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n5450, CK => CLK, Q => 
                           n_1336, QN => n13718);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n5449, CK => CLK, Q => 
                           n_1337, QN => n13719);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n5448, CK => CLK, Q => 
                           n_1338, QN => n13720);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n5447, CK => CLK, Q => 
                           n_1339, QN => n13721);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n5446, CK => CLK, Q => 
                           n_1340, QN => n13722);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n5445, CK => CLK, Q => 
                           n_1341, QN => n13723);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n5444, CK => CLK, Q => 
                           n_1342, QN => n13724);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n5443, CK => CLK, Q => 
                           n_1343, QN => n13725);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n5442, CK => CLK, Q => 
                           n_1344, QN => n13726);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n5441, CK => CLK, Q => 
                           n_1345, QN => n13727);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n5440, CK => CLK, Q => 
                           n_1346, QN => n13728);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n5439, CK => CLK, Q => 
                           n_1347, QN => n13729);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n5438, CK => CLK, Q => 
                           n_1348, QN => n13730);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => n5433, CK => CLK, Q => 
                           n_1349, QN => n13735);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => n5432, CK => CLK, Q => 
                           n_1350, QN => n13736);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => n5431, CK => CLK, Q => 
                           n_1351, QN => n13737);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => n5430, CK => CLK, Q => 
                           n_1352, QN => n13738);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => n5429, CK => CLK, Q => 
                           n_1353, QN => n13739);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => n5428, CK => CLK, Q => 
                           n_1354, QN => n13740);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => n5427, CK => CLK, Q => 
                           n_1355, QN => n13741);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => n5426, CK => CLK, Q => 
                           n_1356, QN => n13742);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n5377, CK => CLK, Q => 
                           n_1357, QN => n13743);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n5376, CK => CLK, Q => 
                           n_1358, QN => n13744);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n5375, CK => CLK, Q => 
                           n_1359, QN => n13745);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n5374, CK => CLK, Q => 
                           n_1360, QN => n13746);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => n5241, CK => CLK, Q => 
                           n_1361, QN => n13751);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => n5240, CK => CLK, Q => 
                           n_1362, QN => n13752);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => n5239, CK => CLK, Q => 
                           n_1363, QN => n13753);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => n5238, CK => CLK, Q => 
                           n_1364, QN => n13754);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => n5237, CK => CLK, Q => 
                           n_1365, QN => n13755);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => n5236, CK => CLK, Q => 
                           n_1366, QN => n13756);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => n5235, CK => CLK, Q => 
                           n_1367, QN => n13757);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => n5234, CK => CLK, Q => 
                           n_1368, QN => n13758);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => n5233, CK => CLK, Q => 
                           n_1369, QN => n13759);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => n5232, CK => CLK, Q => 
                           n_1370, QN => n13760);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => n5231, CK => CLK, Q => 
                           n_1371, QN => n13761);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => n5230, CK => CLK, Q => 
                           n_1372, QN => n13762);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => n5229, CK => CLK, Q => 
                           n_1373, QN => n13763);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => n5228, CK => CLK, Q => 
                           n_1374, QN => n13764);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => n5227, CK => CLK, Q => 
                           n_1375, QN => n13765);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => n5226, CK => CLK, Q => 
                           n_1376, QN => n13766);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => n5225, CK => CLK, Q => 
                           n_1377, QN => n13767);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => n5224, CK => CLK, Q => 
                           n_1378, QN => n13768);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => n5223, CK => CLK, Q => 
                           n_1379, QN => n13769);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => n5222, CK => CLK, Q => 
                           n_1380, QN => n13770);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => n5221, CK => CLK, Q => 
                           n_1381, QN => n13771);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => n5220, CK => CLK, Q => 
                           n_1382, QN => n13772);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => n5219, CK => CLK, Q => 
                           n_1383, QN => n13773);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => n5218, CK => CLK, Q => 
                           n_1384, QN => n13774);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => n5217, CK => CLK, Q => 
                           n_1385, QN => n13775);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => n5216, CK => CLK, Q => 
                           n_1386, QN => n13776);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => n5215, CK => CLK, Q => 
                           n_1387, QN => n13777);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => n5214, CK => CLK, Q => 
                           n_1388, QN => n13778);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n5213, CK => CLK, Q => 
                           n_1389, QN => n13779);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n5212, CK => CLK, Q => 
                           n_1390, QN => n13780);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n5211, CK => CLK, Q => 
                           n_1391, QN => n13781);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n5210, CK => CLK, Q => 
                           n_1392, QN => n13782);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n5209, CK => CLK, Q => 
                           n_1393, QN => n13783);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n5208, CK => CLK, Q => 
                           n_1394, QN => n13784);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n5207, CK => CLK, Q => 
                           n_1395, QN => n13785);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n5206, CK => CLK, Q => 
                           n_1396, QN => n13786);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n5205, CK => CLK, Q => 
                           n_1397, QN => n13787);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n5204, CK => CLK, Q => 
                           n_1398, QN => n13788);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n5203, CK => CLK, Q => 
                           n_1399, QN => n13789);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n5202, CK => CLK, Q => 
                           n_1400, QN => n13790);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n5201, CK => CLK, Q => 
                           n_1401, QN => n13791);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n5200, CK => CLK, Q => 
                           n_1402, QN => n13792);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n5199, CK => CLK, Q => 
                           n_1403, QN => n13793);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n5198, CK => CLK, Q => 
                           n_1404, QN => n13794);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n5197, CK => CLK, Q => 
                           n_1405, QN => n13795);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n5196, CK => CLK, Q => 
                           n_1406, QN => n13796);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n5195, CK => CLK, Q => 
                           n_1407, QN => n13797);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n5194, CK => CLK, Q => 
                           n_1408, QN => n13798);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n5193, CK => CLK, Q => 
                           n_1409, QN => n13799);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n5192, CK => CLK, Q => 
                           n_1410, QN => n13800);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n5191, CK => CLK, Q => 
                           n_1411, QN => n13801);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n5190, CK => CLK, Q => 
                           n_1412, QN => n13802);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n5189, CK => CLK, Q => 
                           n_1413, QN => n13803);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n5188, CK => CLK, Q => 
                           n_1414, QN => n13804);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n5187, CK => CLK, Q => 
                           n_1415, QN => n13805);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n5186, CK => CLK, Q => 
                           n_1416, QN => n13806);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n5185, CK => CLK, Q => 
                           n_1417, QN => n13807);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n5184, CK => CLK, Q => 
                           n_1418, QN => n13808);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n5183, CK => CLK, Q => 
                           n_1419, QN => n13809);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n5182, CK => CLK, Q => 
                           n_1420, QN => n13810);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n5122, CK => CLK, Q => 
                           n_1421, QN => n13811);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n5121, CK => CLK, Q => 
                           n_1422, QN => n13812);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n5120, CK => CLK, Q => 
                           n_1423, QN => n13813);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n5119, CK => CLK, Q => 
                           n_1424, QN => n13814);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n5118, CK => CLK, Q => 
                           n_1425, QN => n13815);
   OUT1_reg_63_inst : DFF_X1 port map( D => n4989, CK => CLK, Q => OUT1(63), QN
                           => n4765);
   OUT1_reg_62_inst : DFF_X1 port map( D => n4988, CK => CLK, Q => OUT1(62), QN
                           => n4766);
   OUT1_reg_61_inst : DFF_X1 port map( D => n4987, CK => CLK, Q => OUT1(61), QN
                           => n4767);
   OUT1_reg_60_inst : DFF_X1 port map( D => n4986, CK => CLK, Q => OUT1(60), QN
                           => n4768);
   OUT1_reg_59_inst : DFF_X1 port map( D => n4985, CK => CLK, Q => OUT1(59), QN
                           => n4769);
   OUT1_reg_58_inst : DFF_X1 port map( D => n4984, CK => CLK, Q => OUT1(58), QN
                           => n4770);
   OUT1_reg_57_inst : DFF_X1 port map( D => n4983, CK => CLK, Q => OUT1(57), QN
                           => n4771);
   OUT1_reg_56_inst : DFF_X1 port map( D => n4982, CK => CLK, Q => OUT1(56), QN
                           => n4772);
   OUT1_reg_55_inst : DFF_X1 port map( D => n4981, CK => CLK, Q => OUT1(55), QN
                           => n4773);
   OUT1_reg_54_inst : DFF_X1 port map( D => n4980, CK => CLK, Q => OUT1(54), QN
                           => n4774);
   OUT1_reg_53_inst : DFF_X1 port map( D => n4979, CK => CLK, Q => OUT1(53), QN
                           => n4775);
   OUT1_reg_52_inst : DFF_X1 port map( D => n4978, CK => CLK, Q => OUT1(52), QN
                           => n4776);
   OUT1_reg_51_inst : DFF_X1 port map( D => n4977, CK => CLK, Q => OUT1(51), QN
                           => n4777);
   OUT1_reg_50_inst : DFF_X1 port map( D => n4976, CK => CLK, Q => OUT1(50), QN
                           => n4778);
   OUT1_reg_49_inst : DFF_X1 port map( D => n4975, CK => CLK, Q => OUT1(49), QN
                           => n4779);
   OUT1_reg_48_inst : DFF_X1 port map( D => n4974, CK => CLK, Q => OUT1(48), QN
                           => n4780);
   OUT1_reg_47_inst : DFF_X1 port map( D => n4973, CK => CLK, Q => OUT1(47), QN
                           => n4781);
   OUT1_reg_46_inst : DFF_X1 port map( D => n4972, CK => CLK, Q => OUT1(46), QN
                           => n4782);
   OUT1_reg_45_inst : DFF_X1 port map( D => n4971, CK => CLK, Q => OUT1(45), QN
                           => n4783);
   OUT1_reg_44_inst : DFF_X1 port map( D => n4970, CK => CLK, Q => OUT1(44), QN
                           => n4784);
   OUT1_reg_43_inst : DFF_X1 port map( D => n4969, CK => CLK, Q => OUT1(43), QN
                           => n4785);
   OUT1_reg_42_inst : DFF_X1 port map( D => n4968, CK => CLK, Q => OUT1(42), QN
                           => n4786);
   OUT1_reg_41_inst : DFF_X1 port map( D => n4967, CK => CLK, Q => OUT1(41), QN
                           => n4787);
   OUT1_reg_40_inst : DFF_X1 port map( D => n4966, CK => CLK, Q => OUT1(40), QN
                           => n4788);
   OUT1_reg_39_inst : DFF_X1 port map( D => n4965, CK => CLK, Q => OUT1(39), QN
                           => n4789);
   OUT1_reg_38_inst : DFF_X1 port map( D => n4964, CK => CLK, Q => OUT1(38), QN
                           => n4790);
   OUT1_reg_37_inst : DFF_X1 port map( D => n4963, CK => CLK, Q => OUT1(37), QN
                           => n4791);
   OUT1_reg_36_inst : DFF_X1 port map( D => n4962, CK => CLK, Q => OUT1(36), QN
                           => n4792);
   OUT1_reg_35_inst : DFF_X1 port map( D => n4961, CK => CLK, Q => OUT1(35), QN
                           => n4793);
   OUT1_reg_34_inst : DFF_X1 port map( D => n4960, CK => CLK, Q => OUT1(34), QN
                           => n4794);
   OUT1_reg_33_inst : DFF_X1 port map( D => n4959, CK => CLK, Q => OUT1(33), QN
                           => n4795);
   OUT1_reg_32_inst : DFF_X1 port map( D => n4958, CK => CLK, Q => OUT1(32), QN
                           => n4796);
   OUT1_reg_31_inst : DFF_X1 port map( D => n4957, CK => CLK, Q => OUT1(31), QN
                           => n4797);
   OUT1_reg_30_inst : DFF_X1 port map( D => n4956, CK => CLK, Q => OUT1(30), QN
                           => n4803);
   OUT1_reg_29_inst : DFF_X1 port map( D => n4955, CK => CLK, Q => OUT1(29), QN
                           => n4804);
   OUT1_reg_28_inst : DFF_X1 port map( D => n4954, CK => CLK, Q => OUT1(28), QN
                           => n4805);
   OUT1_reg_27_inst : DFF_X1 port map( D => n4953, CK => CLK, Q => OUT1(27), QN
                           => n4806);
   OUT1_reg_26_inst : DFF_X1 port map( D => n4952, CK => CLK, Q => OUT1(26), QN
                           => n4807);
   OUT1_reg_25_inst : DFF_X1 port map( D => n4951, CK => CLK, Q => OUT1(25), QN
                           => n4808);
   OUT1_reg_24_inst : DFF_X1 port map( D => n4950, CK => CLK, Q => OUT1(24), QN
                           => n4809);
   OUT1_reg_23_inst : DFF_X1 port map( D => n4949, CK => CLK, Q => OUT1(23), QN
                           => n4810);
   OUT1_reg_22_inst : DFF_X1 port map( D => n4948, CK => CLK, Q => OUT1(22), QN
                           => n4811);
   OUT1_reg_21_inst : DFF_X1 port map( D => n4947, CK => CLK, Q => OUT1(21), QN
                           => n4812);
   OUT1_reg_20_inst : DFF_X1 port map( D => n4946, CK => CLK, Q => OUT1(20), QN
                           => n4813);
   OUT1_reg_19_inst : DFF_X1 port map( D => n4945, CK => CLK, Q => OUT1(19), QN
                           => n4814);
   OUT1_reg_18_inst : DFF_X1 port map( D => n4944, CK => CLK, Q => OUT1(18), QN
                           => n4815);
   OUT1_reg_17_inst : DFF_X1 port map( D => n4943, CK => CLK, Q => OUT1(17), QN
                           => n4816);
   OUT1_reg_16_inst : DFF_X1 port map( D => n4942, CK => CLK, Q => OUT1(16), QN
                           => n4817);
   OUT1_reg_15_inst : DFF_X1 port map( D => n4941, CK => CLK, Q => OUT1(15), QN
                           => n4818);
   OUT1_reg_14_inst : DFF_X1 port map( D => n4940, CK => CLK, Q => OUT1(14), QN
                           => n4819);
   OUT1_reg_13_inst : DFF_X1 port map( D => n4939, CK => CLK, Q => OUT1(13), QN
                           => n4820);
   OUT1_reg_12_inst : DFF_X1 port map( D => n4938, CK => CLK, Q => OUT1(12), QN
                           => n4821);
   OUT1_reg_11_inst : DFF_X1 port map( D => n4937, CK => CLK, Q => OUT1(11), QN
                           => n4822);
   OUT1_reg_10_inst : DFF_X1 port map( D => n4936, CK => CLK, Q => OUT1(10), QN
                           => n4823);
   OUT1_reg_9_inst : DFF_X1 port map( D => n4935, CK => CLK, Q => OUT1(9), QN 
                           => n4824);
   OUT1_reg_8_inst : DFF_X1 port map( D => n4934, CK => CLK, Q => OUT1(8), QN 
                           => n4825);
   OUT1_reg_7_inst : DFF_X1 port map( D => n4933, CK => CLK, Q => OUT1(7), QN 
                           => n4826);
   OUT1_reg_6_inst : DFF_X1 port map( D => n4932, CK => CLK, Q => OUT1(6), QN 
                           => n4827);
   OUT1_reg_5_inst : DFF_X1 port map( D => n4931, CK => CLK, Q => OUT1(5), QN 
                           => n4828);
   OUT1_reg_4_inst : DFF_X1 port map( D => n4930, CK => CLK, Q => OUT1(4), QN 
                           => n4829);
   OUT1_reg_3_inst : DFF_X1 port map( D => n4929, CK => CLK, Q => OUT1(3), QN 
                           => n4830);
   OUT1_reg_2_inst : DFF_X1 port map( D => n4928, CK => CLK, Q => OUT1(2), QN 
                           => n4831);
   OUT1_reg_1_inst : DFF_X1 port map( D => n4927, CK => CLK, Q => OUT1(1), QN 
                           => n4832);
   OUT1_reg_0_inst : DFF_X1 port map( D => n4926, CK => CLK, Q => OUT1(0), QN 
                           => n4833);
   OUT2_reg_63_inst : DFF_X1 port map( D => n4925, CK => CLK, Q => OUT2(63), QN
                           => n4834);
   OUT2_reg_62_inst : DFF_X1 port map( D => n4924, CK => CLK, Q => OUT2(62), QN
                           => n4851);
   OUT2_reg_61_inst : DFF_X1 port map( D => n4923, CK => CLK, Q => OUT2(61), QN
                           => n7112);
   OUT2_reg_60_inst : DFF_X1 port map( D => n4922, CK => CLK, Q => OUT2(60), QN
                           => n7129);
   OUT2_reg_59_inst : DFF_X1 port map( D => n4921, CK => CLK, Q => OUT2(59), QN
                           => n7146);
   OUT2_reg_58_inst : DFF_X1 port map( D => n4920, CK => CLK, Q => OUT2(58), QN
                           => n7243);
   OUT2_reg_57_inst : DFF_X1 port map( D => n4919, CK => CLK, Q => OUT2(57), QN
                           => n7260);
   OUT2_reg_56_inst : DFF_X1 port map( D => n4918, CK => CLK, Q => OUT2(56), QN
                           => n7277);
   OUT2_reg_55_inst : DFF_X1 port map( D => n4917, CK => CLK, Q => OUT2(55), QN
                           => n7376);
   OUT2_reg_54_inst : DFF_X1 port map( D => n4916, CK => CLK, Q => OUT2(54), QN
                           => n7393);
   OUT2_reg_53_inst : DFF_X1 port map( D => n4915, CK => CLK, Q => OUT2(53), QN
                           => n7495);
   OUT2_reg_52_inst : DFF_X1 port map( D => n4914, CK => CLK, Q => OUT2(52), QN
                           => n7512);
   OUT2_reg_51_inst : DFF_X1 port map( D => n4913, CK => CLK, Q => OUT2(51), QN
                           => n7529);
   OUT2_reg_50_inst : DFF_X1 port map( D => n4912, CK => CLK, Q => OUT2(50), QN
                           => n7633);
   OUT2_reg_49_inst : DFF_X1 port map( D => n4911, CK => CLK, Q => OUT2(49), QN
                           => n7650);
   OUT2_reg_48_inst : DFF_X1 port map( D => n4910, CK => CLK, Q => OUT2(48), QN
                           => n7752);
   OUT2_reg_47_inst : DFF_X1 port map( D => n4909, CK => CLK, Q => OUT2(47), QN
                           => n7769);
   OUT2_reg_46_inst : DFF_X1 port map( D => n4908, CK => CLK, Q => OUT2(46), QN
                           => n7786);
   OUT2_reg_45_inst : DFF_X1 port map( D => n4907, CK => CLK, Q => OUT2(45), QN
                           => n7803);
   OUT2_reg_44_inst : DFF_X1 port map( D => n4906, CK => CLK, Q => OUT2(44), QN
                           => n7820);
   OUT2_reg_43_inst : DFF_X1 port map( D => n4905, CK => CLK, Q => OUT2(43), QN
                           => n7837);
   OUT2_reg_42_inst : DFF_X1 port map( D => n4904, CK => CLK, Q => OUT2(42), QN
                           => n7854);
   OUT2_reg_41_inst : DFF_X1 port map( D => n4903, CK => CLK, Q => OUT2(41), QN
                           => n7871);
   OUT2_reg_40_inst : DFF_X1 port map( D => n4902, CK => CLK, Q => OUT2(40), QN
                           => n7888);
   OUT2_reg_39_inst : DFF_X1 port map( D => n4901, CK => CLK, Q => OUT2(39), QN
                           => n7905);
   OUT2_reg_38_inst : DFF_X1 port map( D => n4900, CK => CLK, Q => OUT2(38), QN
                           => n7922);
   OUT2_reg_37_inst : DFF_X1 port map( D => n4899, CK => CLK, Q => OUT2(37), QN
                           => n7939);
   OUT2_reg_36_inst : DFF_X1 port map( D => n4898, CK => CLK, Q => OUT2(36), QN
                           => n7956);
   OUT2_reg_35_inst : DFF_X1 port map( D => n4897, CK => CLK, Q => OUT2(35), QN
                           => n7973);
   OUT2_reg_34_inst : DFF_X1 port map( D => n4896, CK => CLK, Q => OUT2(34), QN
                           => n7990);
   OUT2_reg_33_inst : DFF_X1 port map( D => n4895, CK => CLK, Q => OUT2(33), QN
                           => n8007);
   OUT2_reg_32_inst : DFF_X1 port map( D => n4894, CK => CLK, Q => OUT2(32), QN
                           => n8024);
   OUT2_reg_31_inst : DFF_X1 port map( D => n4893, CK => CLK, Q => OUT2(31), QN
                           => n8041);
   OUT2_reg_30_inst : DFF_X1 port map( D => n4892, CK => CLK, Q => OUT2(30), QN
                           => n8058);
   OUT2_reg_29_inst : DFF_X1 port map( D => n4891, CK => CLK, Q => OUT2(29), QN
                           => n8075);
   OUT2_reg_28_inst : DFF_X1 port map( D => n4890, CK => CLK, Q => OUT2(28), QN
                           => n8092);
   OUT2_reg_27_inst : DFF_X1 port map( D => n4889, CK => CLK, Q => OUT2(27), QN
                           => n8109);
   OUT2_reg_26_inst : DFF_X1 port map( D => n4888, CK => CLK, Q => OUT2(26), QN
                           => n8126);
   OUT2_reg_25_inst : DFF_X1 port map( D => n4887, CK => CLK, Q => OUT2(25), QN
                           => n8143);
   OUT2_reg_24_inst : DFF_X1 port map( D => n4886, CK => CLK, Q => OUT2(24), QN
                           => n8160);
   OUT2_reg_23_inst : DFF_X1 port map( D => n4885, CK => CLK, Q => OUT2(23), QN
                           => n8177);
   OUT2_reg_22_inst : DFF_X1 port map( D => n4884, CK => CLK, Q => OUT2(22), QN
                           => n8194);
   OUT2_reg_21_inst : DFF_X1 port map( D => n4883, CK => CLK, Q => OUT2(21), QN
                           => n8211);
   OUT2_reg_20_inst : DFF_X1 port map( D => n4882, CK => CLK, Q => OUT2(20), QN
                           => n8228);
   OUT2_reg_19_inst : DFF_X1 port map( D => n4881, CK => CLK, Q => OUT2(19), QN
                           => n8245);
   OUT2_reg_18_inst : DFF_X1 port map( D => n4880, CK => CLK, Q => OUT2(18), QN
                           => n8262);
   OUT2_reg_17_inst : DFF_X1 port map( D => n4879, CK => CLK, Q => OUT2(17), QN
                           => n8279);
   OUT2_reg_16_inst : DFF_X1 port map( D => n4878, CK => CLK, Q => OUT2(16), QN
                           => n8296);
   OUT2_reg_15_inst : DFF_X1 port map( D => n4877, CK => CLK, Q => OUT2(15), QN
                           => n8313);
   OUT2_reg_14_inst : DFF_X1 port map( D => n4876, CK => CLK, Q => OUT2(14), QN
                           => n8330);
   OUT2_reg_13_inst : DFF_X1 port map( D => n4875, CK => CLK, Q => OUT2(13), QN
                           => n8347);
   OUT2_reg_12_inst : DFF_X1 port map( D => n4874, CK => CLK, Q => OUT2(12), QN
                           => n8364);
   OUT2_reg_11_inst : DFF_X1 port map( D => n4873, CK => CLK, Q => OUT2(11), QN
                           => n8381);
   OUT2_reg_10_inst : DFF_X1 port map( D => n4872, CK => CLK, Q => OUT2(10), QN
                           => n8398);
   OUT2_reg_9_inst : DFF_X1 port map( D => n4871, CK => CLK, Q => OUT2(9), QN 
                           => n8415);
   OUT2_reg_8_inst : DFF_X1 port map( D => n4870, CK => CLK, Q => OUT2(8), QN 
                           => n8432);
   OUT2_reg_7_inst : DFF_X1 port map( D => n4869, CK => CLK, Q => OUT2(7), QN 
                           => n8449);
   OUT2_reg_6_inst : DFF_X1 port map( D => n4868, CK => CLK, Q => OUT2(6), QN 
                           => n8466);
   OUT2_reg_5_inst : DFF_X1 port map( D => n4867, CK => CLK, Q => OUT2(5), QN 
                           => n8483);
   OUT2_reg_4_inst : DFF_X1 port map( D => n4866, CK => CLK, Q => OUT2(4), QN 
                           => n8500);
   OUT2_reg_3_inst : DFF_X1 port map( D => n4865, CK => CLK, Q => OUT2(3), QN 
                           => n8517);
   OUT2_reg_2_inst : DFF_X1 port map( D => n4864, CK => CLK, Q => OUT2(2), QN 
                           => n8534);
   OUT2_reg_1_inst : DFF_X1 port map( D => n4863, CK => CLK, Q => OUT2(1), QN 
                           => n8551);
   OUT2_reg_0_inst : DFF_X1 port map( D => n4862, CK => CLK, Q => OUT2(0), QN 
                           => n8568);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n6844, CK => CLK, Q => n9950
                           , QN => n11997);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n6843, CK => CLK, Q => n9951
                           , QN => n11996);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n6842, CK => CLK, Q => n9952
                           , QN => n11995);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n5401, CK => CLK, Q => 
                           n_1426, QN => n13869);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n5400, CK => CLK, Q => 
                           n_1427, QN => n13870);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n5399, CK => CLK, Q => 
                           n_1428, QN => n13871);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n5398, CK => CLK, Q => 
                           n_1429, QN => n13872);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n5397, CK => CLK, Q => 
                           n_1430, QN => n13873);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n5396, CK => CLK, Q => 
                           n_1431, QN => n13874);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n5395, CK => CLK, Q => 
                           n_1432, QN => n13875);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n5394, CK => CLK, Q => 
                           n_1433, QN => n13876);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n5393, CK => CLK, Q => 
                           n_1434, QN => n13877);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n5392, CK => CLK, Q => 
                           n_1435, QN => n13878);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n5391, CK => CLK, Q => 
                           n_1436, QN => n13879);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n5390, CK => CLK, Q => 
                           n_1437, QN => n13880);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n5389, CK => CLK, Q => 
                           n_1438, QN => n13881);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n5388, CK => CLK, Q => 
                           n_1439, QN => n13882);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n5387, CK => CLK, Q => 
                           n_1440, QN => n13883);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n5386, CK => CLK, Q => 
                           n_1441, QN => n13884);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n5385, CK => CLK, Q => 
                           n_1442, QN => n13885);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n5384, CK => CLK, Q => 
                           n_1443, QN => n13886);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n5383, CK => CLK, Q => 
                           n_1444, QN => n13887);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n5382, CK => CLK, Q => 
                           n_1445, QN => n13888);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n5381, CK => CLK, Q => 
                           n_1446, QN => n13889);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n5380, CK => CLK, Q => 
                           n_1447, QN => n13890);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n5379, CK => CLK, Q => 
                           n_1448, QN => n13891);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n5378, CK => CLK, Q => 
                           n_1449, QN => n13892);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => n5157, CK => CLK, Q => 
                           n_1450, QN => n13929);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => n5156, CK => CLK, Q => 
                           n_1451, QN => n13930);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => n5155, CK => CLK, Q => 
                           n_1452, QN => n13931);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => n5154, CK => CLK, Q => 
                           n_1453, QN => n13932);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => n5153, CK => CLK, Q => 
                           n_1454, QN => n13933);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => n5152, CK => CLK, Q => 
                           n_1455, QN => n13934);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => n5151, CK => CLK, Q => 
                           n_1456, QN => n13935);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => n5150, CK => CLK, Q => 
                           n_1457, QN => n13936);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n5149, CK => CLK, Q => 
                           n_1458, QN => n13937);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n5148, CK => CLK, Q => 
                           n_1459, QN => n13938);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n5147, CK => CLK, Q => 
                           n_1460, QN => n13939);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n5146, CK => CLK, Q => 
                           n_1461, QN => n13940);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n5145, CK => CLK, Q => 
                           n_1462, QN => n13941);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n5144, CK => CLK, Q => 
                           n_1463, QN => n13942);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n5143, CK => CLK, Q => 
                           n_1464, QN => n13943);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n5142, CK => CLK, Q => 
                           n_1465, QN => n13944);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n5141, CK => CLK, Q => 
                           n_1466, QN => n13945);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n5140, CK => CLK, Q => 
                           n_1467, QN => n13946);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n5139, CK => CLK, Q => 
                           n_1468, QN => n13947);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n5138, CK => CLK, Q => 
                           n_1469, QN => n13948);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n5137, CK => CLK, Q => 
                           n_1470, QN => n13949);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n5136, CK => CLK, Q => 
                           n_1471, QN => n13950);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n5135, CK => CLK, Q => 
                           n_1472, QN => n13951);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n5134, CK => CLK, Q => 
                           n_1473, QN => n13952);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n5133, CK => CLK, Q => 
                           n_1474, QN => n14025);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n5132, CK => CLK, Q => 
                           n_1475, QN => n14026);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n5131, CK => CLK, Q => 
                           n_1476, QN => n14027);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n5130, CK => CLK, Q => 
                           n_1477, QN => n14028);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n5129, CK => CLK, Q => 
                           n_1478, QN => n14029);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n5128, CK => CLK, Q => 
                           n_1479, QN => n14030);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n5127, CK => CLK, Q => 
                           n_1480, QN => n14031);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n5126, CK => CLK, Q => 
                           n_1481, QN => n14032);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n5125, CK => CLK, Q => 
                           n_1482, QN => n14033);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n5124, CK => CLK, Q => 
                           n_1483, QN => n14034);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n5123, CK => CLK, Q => 
                           n_1484, QN => n14035);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => n5425, CK => CLK, Q => 
                           n_1485, QN => n14036);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => n5424, CK => CLK, Q => 
                           n_1486, QN => n14037);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => n5423, CK => CLK, Q => 
                           n_1487, QN => n14038);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => n5422, CK => CLK, Q => 
                           n_1488, QN => n14039);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => n5421, CK => CLK, Q => 
                           n_1489, QN => n14040);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => n5420, CK => CLK, Q => 
                           n_1490, QN => n14041);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => n5419, CK => CLK, Q => 
                           n_1491, QN => n14042);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => n5418, CK => CLK, Q => 
                           n_1492, QN => n14043);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => n5417, CK => CLK, Q => 
                           n_1493, QN => n14044);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => n5416, CK => CLK, Q => 
                           n_1494, QN => n14045);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => n5415, CK => CLK, Q => 
                           n_1495, QN => n14046);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => n5414, CK => CLK, Q => 
                           n_1496, QN => n14047);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => n5413, CK => CLK, Q => 
                           n_1497, QN => n14048);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => n5412, CK => CLK, Q => 
                           n_1498, QN => n14049);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => n5411, CK => CLK, Q => 
                           n_1499, QN => n14050);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => n5410, CK => CLK, Q => 
                           n_1500, QN => n14051);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => n5409, CK => CLK, Q => 
                           n_1501, QN => n14052);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => n5408, CK => CLK, Q => 
                           n_1502, QN => n14053);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => n5407, CK => CLK, Q => 
                           n_1503, QN => n14054);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => n5406, CK => CLK, Q => 
                           n_1504, QN => n14055);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n5405, CK => CLK, Q => 
                           n_1505, QN => n14056);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n5404, CK => CLK, Q => 
                           n_1506, QN => n14057);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n5403, CK => CLK, Q => 
                           n_1507, QN => n14058);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n5402, CK => CLK, Q => 
                           n_1508, QN => n14059);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => n5177, CK => CLK, Q => 
                           n_1509, QN => n14087);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => n5176, CK => CLK, Q => 
                           n_1510, QN => n14088);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => n5175, CK => CLK, Q => 
                           n_1511, QN => n14089);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => n5174, CK => CLK, Q => 
                           n_1512, QN => n14090);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => n5173, CK => CLK, Q => 
                           n_1513, QN => n14091);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => n5172, CK => CLK, Q => 
                           n_1514, QN => n14092);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => n5171, CK => CLK, Q => 
                           n_1515, QN => n14093);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => n5170, CK => CLK, Q => 
                           n_1516, QN => n14094);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => n5169, CK => CLK, Q => 
                           n_1517, QN => n14095);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => n5168, CK => CLK, Q => 
                           n_1518, QN => n14096);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => n5167, CK => CLK, Q => 
                           n_1519, QN => n14097);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => n5166, CK => CLK, Q => 
                           n_1520, QN => n14098);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => n5165, CK => CLK, Q => 
                           n_1521, QN => n14099);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => n5164, CK => CLK, Q => 
                           n_1522, QN => n14100);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => n5163, CK => CLK, Q => 
                           n_1523, QN => n14101);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => n5162, CK => CLK, Q => 
                           n_1524, QN => n14102);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => n5161, CK => CLK, Q => 
                           n_1525, QN => n14103);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => n5160, CK => CLK, Q => 
                           n_1526, QN => n14104);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => n5159, CK => CLK, Q => 
                           n_1527, QN => n14105);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => n5158, CK => CLK, Q => 
                           n_1528, QN => n14106);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n5527, CK => CLK, Q => 
                           n7199, QN => n11935);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n5526, CK => CLK, Q => 
                           n7195, QN => n11934);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n5525, CK => CLK, Q => 
                           n7191, QN => n11842);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n5524, CK => CLK, Q => 
                           n7187, QN => n11841);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n5523, CK => CLK, Q => 
                           n7183, QN => n11840);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n5522, CK => CLK, Q => 
                           n7179, QN => n11839);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n5521, CK => CLK, Q => 
                           n7175, QN => n11838);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n5520, CK => CLK, Q => 
                           n7171, QN => n11837);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n5519, CK => CLK, Q => 
                           n7167, QN => n11836);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n5518, CK => CLK, Q => 
                           n7163, QN => n11835);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n5517, CK => CLK, Q => 
                           n7159, QN => n11834);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n5516, CK => CLK, Q => 
                           n7155, QN => n11833);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => n5664, CK => CLK, Q => 
                           n_1529, QN => n8001);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => n5663, CK => CLK, Q => 
                           n_1530, QN => n8018);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => n5662, CK => CLK, Q => 
                           n_1531, QN => n8035);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n5661, CK => CLK, Q => 
                           n_1532, QN => n8052);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n5660, CK => CLK, Q => 
                           n_1533, QN => n8069);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n5659, CK => CLK, Q => 
                           n_1534, QN => n8086);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n5658, CK => CLK, Q => 
                           n_1535, QN => n8103);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n5657, CK => CLK, Q => 
                           n_1536, QN => n8120);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n5656, CK => CLK, Q => 
                           n_1537, QN => n8137);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n5655, CK => CLK, Q => 
                           n_1538, QN => n8154);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n5654, CK => CLK, Q => 
                           n_1539, QN => n8171);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => n5753, CK => CLK, Q => 
                           n_1540, QN => n7238);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => n5752, CK => CLK, Q => 
                           n_1541, QN => n7255);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => n5751, CK => CLK, Q => 
                           n_1542, QN => n7272);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => n5750, CK => CLK, Q => 
                           n_1543, QN => n7371);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => n5749, CK => CLK, Q => 
                           n_1544, QN => n7388);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => n5748, CK => CLK, Q => 
                           n_1545, QN => n7490);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => n5747, CK => CLK, Q => 
                           n_1546, QN => n7507);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => n5746, CK => CLK, Q => 
                           n_1547, QN => n7524);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => n5745, CK => CLK, Q => 
                           n_1548, QN => n7628);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => n5744, CK => CLK, Q => 
                           n_1549, QN => n7645);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => n5743, CK => CLK, Q => 
                           n_1550, QN => n7747);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => n5742, CK => CLK, Q => 
                           n_1551, QN => n7764);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => n5741, CK => CLK, Q => 
                           n_1552, QN => n7781);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => n5740, CK => CLK, Q => 
                           n_1553, QN => n7798);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => n5739, CK => CLK, Q => 
                           n_1554, QN => n7815);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => n5738, CK => CLK, Q => 
                           n_1555, QN => n7832);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => n5737, CK => CLK, Q => 
                           n_1556, QN => n7849);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => n5736, CK => CLK, Q => 
                           n_1557, QN => n7866);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => n5735, CK => CLK, Q => 
                           n_1558, QN => n7883);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => n5734, CK => CLK, Q => 
                           n_1559, QN => n7900);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => n5733, CK => CLK, Q => 
                           n_1560, QN => n7917);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => n5732, CK => CLK, Q => 
                           n_1561, QN => n7934);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => n5731, CK => CLK, Q => 
                           n_1562, QN => n7951);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => n5730, CK => CLK, Q => 
                           n_1563, QN => n7968);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => n5729, CK => CLK, Q => 
                           n_1564, QN => n7985);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => n5728, CK => CLK, Q => 
                           n_1565, QN => n8002);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => n5727, CK => CLK, Q => 
                           n_1566, QN => n8019);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => n5726, CK => CLK, Q => 
                           n_1567, QN => n8036);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n5725, CK => CLK, Q => 
                           n_1568, QN => n8053);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n5724, CK => CLK, Q => 
                           n_1569, QN => n8070);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n5723, CK => CLK, Q => 
                           n_1570, QN => n8087);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n5722, CK => CLK, Q => 
                           n_1571, QN => n8104);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n5721, CK => CLK, Q => 
                           n_1572, QN => n8121);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n5720, CK => CLK, Q => 
                           n_1573, QN => n8138);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n5719, CK => CLK, Q => 
                           n_1574, QN => n8155);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n5718, CK => CLK, Q => 
                           n_1575, QN => n8172);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n5781, CK => CLK, Q => 
                           n8650, QN => n11832);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n5780, CK => CLK, Q => 
                           n8648, QN => n11831);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n5779, CK => CLK, Q => 
                           n8646, QN => n11830);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n5778, CK => CLK, Q => 
                           n8644, QN => n11829);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n5777, CK => CLK, Q => 
                           n8642, QN => n11828);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n5776, CK => CLK, Q => 
                           n8640, QN => n11827);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n5775, CK => CLK, Q => 
                           n8638, QN => n11826);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n5773, CK => CLK, Q => 
                           n8634, QN => n11825);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n5772, CK => CLK, Q => 
                           n8632, QN => n11824);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n5771, CK => CLK, Q => 
                           n8630, QN => n11823);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n5770, CK => CLK, Q => 
                           n8628, QN => n11822);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n5766, CK => CLK, Q => n8620
                           , QN => n11821);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => n5945, CK => CLK, Q => 
                           n_1576, QN => n7235);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => n5944, CK => CLK, Q => 
                           n_1577, QN => n7252);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => n5943, CK => CLK, Q => 
                           n_1578, QN => n7269);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => n5942, CK => CLK, Q => 
                           n_1579, QN => n7368);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => n5941, CK => CLK, Q => 
                           n_1580, QN => n7385);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => n5940, CK => CLK, Q => 
                           n_1581, QN => n7402);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => n5939, CK => CLK, Q => 
                           n_1582, QN => n7504);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => n5938, CK => CLK, Q => 
                           n_1583, QN => n7521);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => n5937, CK => CLK, Q => 
                           n_1584, QN => n7625);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => n5936, CK => CLK, Q => 
                           n_1585, QN => n7642);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => n5935, CK => CLK, Q => 
                           n_1586, QN => n7744);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => n5934, CK => CLK, Q => 
                           n_1587, QN => n7761);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => n5933, CK => CLK, Q => 
                           n_1588, QN => n7778);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => n5932, CK => CLK, Q => 
                           n_1589, QN => n7795);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => n5931, CK => CLK, Q => 
                           n_1590, QN => n7812);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => n5930, CK => CLK, Q => 
                           n_1591, QN => n7829);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => n5929, CK => CLK, Q => 
                           n_1592, QN => n7846);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => n5928, CK => CLK, Q => 
                           n_1593, QN => n7863);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => n5927, CK => CLK, Q => 
                           n_1594, QN => n7880);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => n5926, CK => CLK, Q => 
                           n_1595, QN => n7897);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => n5925, CK => CLK, Q => 
                           n_1596, QN => n7914);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => n5924, CK => CLK, Q => 
                           n_1597, QN => n7931);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => n5923, CK => CLK, Q => 
                           n_1598, QN => n7948);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => n5922, CK => CLK, Q => 
                           n_1599, QN => n7965);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => n5921, CK => CLK, Q => 
                           n_1600, QN => n7982);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => n5920, CK => CLK, Q => 
                           n_1601, QN => n7999);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => n5919, CK => CLK, Q => 
                           n_1602, QN => n8016);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => n5918, CK => CLK, Q => 
                           n_1603, QN => n8033);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n5917, CK => CLK, Q => 
                           n_1604, QN => n8050);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n5916, CK => CLK, Q => 
                           n_1605, QN => n8067);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n5915, CK => CLK, Q => 
                           n_1606, QN => n8084);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n5914, CK => CLK, Q => 
                           n_1607, QN => n8101);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n5913, CK => CLK, Q => 
                           n_1608, QN => n8118);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n5912, CK => CLK, Q => 
                           n_1609, QN => n8135);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n5911, CK => CLK, Q => 
                           n_1610, QN => n8152);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n5910, CK => CLK, Q => 
                           n_1611, QN => n8169);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => n6009, CK => CLK, Q => 
                           n_1612, QN => n7236);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => n6008, CK => CLK, Q => 
                           n_1613, QN => n7253);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => n6007, CK => CLK, Q => 
                           n_1614, QN => n7270);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => n6006, CK => CLK, Q => 
                           n_1615, QN => n7369);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => n6005, CK => CLK, Q => 
                           n_1616, QN => n7386);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => n6004, CK => CLK, Q => 
                           n_1617, QN => n7403);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => n6003, CK => CLK, Q => 
                           n_1618, QN => n7505);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => n6002, CK => CLK, Q => 
                           n_1619, QN => n7522);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => n6001, CK => CLK, Q => 
                           n_1620, QN => n7626);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => n6000, CK => CLK, Q => 
                           n_1621, QN => n7643);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => n5999, CK => CLK, Q => 
                           n_1622, QN => n7745);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => n5998, CK => CLK, Q => 
                           n_1623, QN => n7762);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => n5997, CK => CLK, Q => 
                           n_1624, QN => n7779);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => n5996, CK => CLK, Q => 
                           n_1625, QN => n7796);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => n5995, CK => CLK, Q => 
                           n_1626, QN => n7813);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => n5994, CK => CLK, Q => 
                           n_1627, QN => n7830);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => n5993, CK => CLK, Q => 
                           n_1628, QN => n7847);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => n5992, CK => CLK, Q => 
                           n_1629, QN => n7864);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => n5991, CK => CLK, Q => 
                           n_1630, QN => n7881);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => n5990, CK => CLK, Q => 
                           n_1631, QN => n7898);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => n5989, CK => CLK, Q => 
                           n_1632, QN => n7915);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => n5988, CK => CLK, Q => 
                           n_1633, QN => n7932);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => n5987, CK => CLK, Q => 
                           n_1634, QN => n7949);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => n5986, CK => CLK, Q => 
                           n_1635, QN => n7966);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => n5985, CK => CLK, Q => 
                           n_1636, QN => n7983);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => n5984, CK => CLK, Q => 
                           n_1637, QN => n8000);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => n5983, CK => CLK, Q => 
                           n_1638, QN => n8017);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => n5982, CK => CLK, Q => 
                           n_1639, QN => n8034);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n5981, CK => CLK, Q => 
                           n_1640, QN => n8051);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n5980, CK => CLK, Q => 
                           n_1641, QN => n8068);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n5979, CK => CLK, Q => 
                           n_1642, QN => n8085);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n5978, CK => CLK, Q => 
                           n_1643, QN => n8102);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n5977, CK => CLK, Q => 
                           n_1644, QN => n8119);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n5976, CK => CLK, Q => 
                           n_1645, QN => n8136);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n5975, CK => CLK, Q => 
                           n_1646, QN => n8153);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n5974, CK => CLK, Q => 
                           n_1647, QN => n8170);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n5515, CK => CLK, Q => 
                           n7131, QN => n11820);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n5514, CK => CLK, Q => 
                           n7105, QN => n11819);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n5513, CK => CLK, Q => 
                           n7101, QN => n11818);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n5512, CK => CLK, Q => 
                           n7097, QN => n11817);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n5511, CK => CLK, Q => n7093
                           , QN => n11816);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n5510, CK => CLK, Q => n7089
                           , QN => n11815);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n5509, CK => CLK, Q => n7085
                           , QN => n11814);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n5508, CK => CLK, Q => n8614
                           , QN => n11813);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n5507, CK => CLK, Q => n8606
                           , QN => n11812);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n5506, CK => CLK, Q => n7081
                           , QN => n11811);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n5769, CK => CLK, Q => 
                           n8626, QN => n11810);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n5768, CK => CLK, Q => 
                           n8624, QN => n11809);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n5767, CK => CLK, Q => n8622
                           , QN => n11808);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n5765, CK => CLK, Q => n8618
                           , QN => n11807);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n5764, CK => CLK, Q => n8612
                           , QN => n11806);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n5763, CK => CLK, Q => n8604
                           , QN => n11805);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n5762, CK => CLK, Q => n8600
                           , QN => n11804);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => n5551, CK => CLK, Q => 
                           n7323, QN => n11933);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => n5550, CK => CLK, Q => 
                           n7319, QN => n11932);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => n5549, CK => CLK, Q => 
                           n7315, QN => n11931);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => n5548, CK => CLK, Q => 
                           n7311, QN => n11930);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => n5547, CK => CLK, Q => 
                           n7307, QN => n11929);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => n5546, CK => CLK, Q => 
                           n7303, QN => n11928);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => n5545, CK => CLK, Q => 
                           n7299, QN => n11927);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => n5544, CK => CLK, Q => 
                           n7295, QN => n11926);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => n5543, CK => CLK, Q => 
                           n7291, QN => n11925);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => n5542, CK => CLK, Q => 
                           n7287, QN => n11924);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => n5541, CK => CLK, Q => 
                           n7283, QN => n11923);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => n5540, CK => CLK, Q => 
                           n7279, QN => n11922);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => n5539, CK => CLK, Q => 
                           n8697, QN => n11921);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => n5538, CK => CLK, Q => 
                           n8698, QN => n11920);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => n5537, CK => CLK, Q => 
                           n8699, QN => n11919);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => n5536, CK => CLK, Q => 
                           n8700, QN => n11918);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => n5535, CK => CLK, Q => 
                           n8701, QN => n11917);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => n5534, CK => CLK, Q => 
                           n8702, QN => n11916);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n5533, CK => CLK, Q => 
                           n8703, QN => n11915);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n5532, CK => CLK, Q => 
                           n8704, QN => n11914);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n5531, CK => CLK, Q => 
                           n8705, QN => n11913);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n5530, CK => CLK, Q => 
                           n8706, QN => n11912);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n5529, CK => CLK, Q => 
                           n8707, QN => n11911);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n5528, CK => CLK, Q => 
                           n8708, QN => n11910);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n5653, CK => CLK, Q => 
                           n_1648, QN => n8188);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n5652, CK => CLK, Q => 
                           n_1649, QN => n8205);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n5651, CK => CLK, Q => 
                           n_1650, QN => n8222);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n5650, CK => CLK, Q => 
                           n_1651, QN => n8239);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n5649, CK => CLK, Q => 
                           n_1652, QN => n8256);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n5648, CK => CLK, Q => 
                           n_1653, QN => n8273);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n5647, CK => CLK, Q => 
                           n_1654, QN => n8290);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n5646, CK => CLK, Q => 
                           n_1655, QN => n8307);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n5645, CK => CLK, Q => 
                           n_1656, QN => n8324);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n5644, CK => CLK, Q => 
                           n_1657, QN => n8341);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n5643, CK => CLK, Q => 
                           n_1658, QN => n8358);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n5642, CK => CLK, Q => 
                           n_1659, QN => n8375);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n5641, CK => CLK, Q => 
                           n_1660, QN => n8392);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n5640, CK => CLK, Q => 
                           n_1661, QN => n8409);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n5639, CK => CLK, Q => 
                           n_1662, QN => n8426);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n5638, CK => CLK, Q => 
                           n_1663, QN => n8443);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n5637, CK => CLK, Q => 
                           n_1664, QN => n8460);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n5636, CK => CLK, Q => 
                           n_1665, QN => n8477);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n5635, CK => CLK, Q => 
                           n_1666, QN => n8494);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n5634, CK => CLK, Q => 
                           n_1667, QN => n8511);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n5633, CK => CLK, Q => 
                           n_1668, QN => n8528);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n5632, CK => CLK, Q => 
                           n_1669, QN => n8545);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n5631, CK => CLK, Q => 
                           n_1670, QN => n8562);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n5630, CK => CLK, Q => 
                           n_1671, QN => n8579);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n5717, CK => CLK, Q => 
                           n_1672, QN => n8189);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n5716, CK => CLK, Q => 
                           n_1673, QN => n8206);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n5715, CK => CLK, Q => 
                           n_1674, QN => n8223);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n5714, CK => CLK, Q => 
                           n_1675, QN => n8240);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n5713, CK => CLK, Q => 
                           n_1676, QN => n8257);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n5712, CK => CLK, Q => 
                           n_1677, QN => n8274);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n5711, CK => CLK, Q => 
                           n_1678, QN => n8291);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n5710, CK => CLK, Q => 
                           n_1679, QN => n8308);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n5709, CK => CLK, Q => 
                           n_1680, QN => n8325);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n5708, CK => CLK, Q => 
                           n_1681, QN => n8342);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n5707, CK => CLK, Q => 
                           n_1682, QN => n8359);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n5706, CK => CLK, Q => 
                           n_1683, QN => n8376);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n5705, CK => CLK, Q => 
                           n_1684, QN => n8393);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n5704, CK => CLK, Q => 
                           n_1685, QN => n8410);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n5703, CK => CLK, Q => 
                           n_1686, QN => n8427);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n5702, CK => CLK, Q => 
                           n_1687, QN => n8444);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n5701, CK => CLK, Q => 
                           n_1688, QN => n8461);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n5700, CK => CLK, Q => 
                           n_1689, QN => n8478);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n5699, CK => CLK, Q => 
                           n_1690, QN => n8495);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n5698, CK => CLK, Q => 
                           n_1691, QN => n8512);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n5697, CK => CLK, Q => 
                           n_1692, QN => n8529);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n5696, CK => CLK, Q => 
                           n_1693, QN => n8546);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n5695, CK => CLK, Q => 
                           n_1694, QN => n8563);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n5694, CK => CLK, Q => 
                           n_1695, QN => n8580);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => n5804, CK => CLK, Q => 
                           n8696, QN => n11909);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => n5803, CK => CLK, Q => 
                           n8694, QN => n11908);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => n5802, CK => CLK, Q => 
                           n8692, QN => n11907);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => n5801, CK => CLK, Q => 
                           n8690, QN => n11906);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => n5800, CK => CLK, Q => 
                           n8688, QN => n11905);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => n5799, CK => CLK, Q => 
                           n8686, QN => n11904);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => n5798, CK => CLK, Q => 
                           n8684, QN => n11903);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => n5797, CK => CLK, Q => 
                           n8682, QN => n11902);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => n5796, CK => CLK, Q => 
                           n8680, QN => n11901);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => n5795, CK => CLK, Q => 
                           n8678, QN => n11900);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => n5794, CK => CLK, Q => 
                           n8676, QN => n11899);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => n5793, CK => CLK, Q => 
                           n8674, QN => n11898);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => n5792, CK => CLK, Q => 
                           n8672, QN => n11897);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => n5791, CK => CLK, Q => 
                           n8670, QN => n11896);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => n5790, CK => CLK, Q => 
                           n8668, QN => n11895);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n5789, CK => CLK, Q => 
                           n8666, QN => n11894);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n5788, CK => CLK, Q => 
                           n8664, QN => n11893);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n5787, CK => CLK, Q => 
                           n8662, QN => n11892);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n5786, CK => CLK, Q => 
                           n8660, QN => n11891);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n5785, CK => CLK, Q => 
                           n8658, QN => n11890);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n5784, CK => CLK, Q => 
                           n8656, QN => n11889);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n5783, CK => CLK, Q => 
                           n8654, QN => n11888);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n5782, CK => CLK, Q => 
                           n8652, QN => n11887);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n5774, CK => CLK, Q => 
                           n8636, QN => n11803);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n5909, CK => CLK, Q => 
                           n_1696, QN => n8186);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n5908, CK => CLK, Q => 
                           n_1697, QN => n8203);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n5907, CK => CLK, Q => 
                           n_1698, QN => n8220);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n5906, CK => CLK, Q => 
                           n_1699, QN => n8237);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n5905, CK => CLK, Q => 
                           n_1700, QN => n8254);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n5904, CK => CLK, Q => 
                           n_1701, QN => n8271);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n5903, CK => CLK, Q => 
                           n_1702, QN => n8288);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n5902, CK => CLK, Q => 
                           n_1703, QN => n8305);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n5901, CK => CLK, Q => 
                           n_1704, QN => n8322);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n5900, CK => CLK, Q => 
                           n_1705, QN => n8339);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n5899, CK => CLK, Q => 
                           n_1706, QN => n8356);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n5898, CK => CLK, Q => 
                           n_1707, QN => n8373);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n5897, CK => CLK, Q => 
                           n_1708, QN => n8390);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n5896, CK => CLK, Q => 
                           n_1709, QN => n8407);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n5895, CK => CLK, Q => 
                           n_1710, QN => n8424);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n5894, CK => CLK, Q => 
                           n_1711, QN => n8441);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n5893, CK => CLK, Q => 
                           n_1712, QN => n8458);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n5892, CK => CLK, Q => 
                           n_1713, QN => n8475);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n5891, CK => CLK, Q => 
                           n_1714, QN => n8492);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n5890, CK => CLK, Q => 
                           n_1715, QN => n8509);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n5889, CK => CLK, Q => 
                           n_1716, QN => n8526);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n5888, CK => CLK, Q => 
                           n_1717, QN => n8543);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n5887, CK => CLK, Q => 
                           n_1718, QN => n8560);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n5886, CK => CLK, Q => 
                           n_1719, QN => n8577);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n5973, CK => CLK, Q => 
                           n_1720, QN => n8187);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n5972, CK => CLK, Q => 
                           n_1721, QN => n8204);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n5971, CK => CLK, Q => 
                           n_1722, QN => n8221);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n5970, CK => CLK, Q => 
                           n_1723, QN => n8238);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n5969, CK => CLK, Q => 
                           n_1724, QN => n8255);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n5968, CK => CLK, Q => 
                           n_1725, QN => n8272);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n5967, CK => CLK, Q => 
                           n_1726, QN => n8289);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n5966, CK => CLK, Q => 
                           n_1727, QN => n8306);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n5965, CK => CLK, Q => 
                           n_1728, QN => n8323);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n5964, CK => CLK, Q => 
                           n_1729, QN => n8340);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n5963, CK => CLK, Q => 
                           n_1730, QN => n8357);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n5962, CK => CLK, Q => 
                           n_1731, QN => n8374);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n5961, CK => CLK, Q => 
                           n_1732, QN => n8391);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n5960, CK => CLK, Q => 
                           n_1733, QN => n8408);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n5959, CK => CLK, Q => 
                           n_1734, QN => n8425);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n5958, CK => CLK, Q => 
                           n_1735, QN => n8442);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n5957, CK => CLK, Q => 
                           n_1736, QN => n8459);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n5956, CK => CLK, Q => 
                           n_1737, QN => n8476);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n5955, CK => CLK, Q => 
                           n_1738, QN => n8493);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n5954, CK => CLK, Q => 
                           n_1739, QN => n8510);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n5953, CK => CLK, Q => 
                           n_1740, QN => n8527);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n5952, CK => CLK, Q => 
                           n_1741, QN => n8544);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n5951, CK => CLK, Q => 
                           n_1742, QN => n8561);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n5950, CK => CLK, Q => 
                           n_1743, QN => n8578);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n6974, CK => CLK, Q => n_1744
                           , QN => n14216);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => n6585, CK => CLK, Q => 
                           n11765, QN => n7150);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => n6584, CK => CLK, Q => 
                           n11641, QN => n7247);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => n6583, CK => CLK, Q => 
                           n11640, QN => n7264);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => n6582, CK => CLK, Q => 
                           n11639, QN => n7363);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => n6581, CK => CLK, Q => 
                           n11638, QN => n7380);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => n6580, CK => CLK, Q => 
                           n11637, QN => n7397);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => n6579, CK => CLK, Q => 
                           n11636, QN => n7499);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => n6578, CK => CLK, Q => 
                           n11635, QN => n7516);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => n6577, CK => CLK, Q => 
                           n11634, QN => n7620);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => n6576, CK => CLK, Q => 
                           n11633, QN => n7637);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => n6575, CK => CLK, Q => 
                           n11632, QN => n7654);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => n6574, CK => CLK, Q => 
                           n11631, QN => n7756);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => n6573, CK => CLK, Q => 
                           n11630, QN => n7773);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => n6572, CK => CLK, Q => 
                           n11629, QN => n7790);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => n6571, CK => CLK, Q => 
                           n11628, QN => n7807);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => n6570, CK => CLK, Q => 
                           n11627, QN => n7824);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => n6569, CK => CLK, Q => 
                           n11626, QN => n7841);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => n6568, CK => CLK, Q => 
                           n11625, QN => n7858);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => n6567, CK => CLK, Q => 
                           n11624, QN => n7875);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => n6566, CK => CLK, Q => 
                           n11623, QN => n7892);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => n6565, CK => CLK, Q => 
                           n11622, QN => n7909);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => n6564, CK => CLK, Q => 
                           n11621, QN => n7926);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => n6563, CK => CLK, Q => 
                           n11620, QN => n7943);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => n6562, CK => CLK, Q => 
                           n11619, QN => n7960);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => n6561, CK => CLK, Q => 
                           n11618, QN => n7977);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => n6560, CK => CLK, Q => 
                           n11617, QN => n7994);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => n6559, CK => CLK, Q => 
                           n11616, QN => n8011);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => n6558, CK => CLK, Q => 
                           n11615, QN => n8028);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n6557, CK => CLK, Q => 
                           n11614, QN => n8045);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n6556, CK => CLK, Q => 
                           n11613, QN => n8062);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n6555, CK => CLK, Q => 
                           n11612, QN => n8079);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n6554, CK => CLK, Q => 
                           n11611, QN => n8096);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n6553, CK => CLK, Q => 
                           n11610, QN => n8113);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n6552, CK => CLK, Q => 
                           n11609, QN => n8130);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n6551, CK => CLK, Q => 
                           n11608, QN => n8147);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n6550, CK => CLK, Q => 
                           n11607, QN => n8164);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => n6649, CK => CLK, Q => 
                           n11585, QN => n7149);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => n6648, CK => CLK, Q => 
                           n11461, QN => n7246);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => n6647, CK => CLK, Q => 
                           n11460, QN => n7263);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => n6646, CK => CLK, Q => 
                           n11459, QN => n7362);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => n6645, CK => CLK, Q => 
                           n11458, QN => n7379);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => n6644, CK => CLK, Q => 
                           n11457, QN => n7396);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => n6643, CK => CLK, Q => 
                           n11456, QN => n7498);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => n6642, CK => CLK, Q => 
                           n11455, QN => n7515);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => n6641, CK => CLK, Q => 
                           n11454, QN => n7619);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => n6640, CK => CLK, Q => 
                           n11453, QN => n7636);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => n6639, CK => CLK, Q => 
                           n11452, QN => n7653);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => n6638, CK => CLK, Q => 
                           n11451, QN => n7755);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => n6637, CK => CLK, Q => 
                           n11450, QN => n7772);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => n6636, CK => CLK, Q => 
                           n11449, QN => n7789);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => n6635, CK => CLK, Q => 
                           n11448, QN => n7806);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => n6634, CK => CLK, Q => 
                           n11447, QN => n7823);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => n6633, CK => CLK, Q => 
                           n11446, QN => n7840);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => n6632, CK => CLK, Q => 
                           n11445, QN => n7857);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => n6631, CK => CLK, Q => 
                           n11444, QN => n7874);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => n6630, CK => CLK, Q => 
                           n11443, QN => n7891);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => n6629, CK => CLK, Q => 
                           n11442, QN => n7908);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => n6628, CK => CLK, Q => 
                           n11441, QN => n7925);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => n6627, CK => CLK, Q => 
                           n11440, QN => n7942);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => n6626, CK => CLK, Q => 
                           n11439, QN => n7959);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => n6625, CK => CLK, Q => 
                           n11438, QN => n7976);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => n6624, CK => CLK, Q => 
                           n11437, QN => n7993);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => n6623, CK => CLK, Q => 
                           n11436, QN => n8010);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => n6622, CK => CLK, Q => 
                           n11435, QN => n8027);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n6621, CK => CLK, Q => 
                           n11434, QN => n8044);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n6620, CK => CLK, Q => 
                           n11433, QN => n8061);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n6619, CK => CLK, Q => 
                           n11432, QN => n8078);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n6618, CK => CLK, Q => 
                           n11431, QN => n8095);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n6617, CK => CLK, Q => 
                           n11430, QN => n8112);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n6616, CK => CLK, Q => 
                           n11429, QN => n8129);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n6615, CK => CLK, Q => 
                           n11428, QN => n8146);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n6614, CK => CLK, Q => 
                           n11427, QN => n8163);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => n6713, CK => CLK, Q => 
                           n_1745, QN => n14217);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => n6712, CK => CLK, Q => 
                           n_1746, QN => n14218);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => n6711, CK => CLK, Q => 
                           n_1747, QN => n14219);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => n6710, CK => CLK, Q => 
                           n_1748, QN => n14220);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => n6709, CK => CLK, Q => 
                           n_1749, QN => n14221);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => n6708, CK => CLK, Q => 
                           n_1750, QN => n14222);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => n6707, CK => CLK, Q => 
                           n_1751, QN => n14223);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => n6706, CK => CLK, Q => 
                           n_1752, QN => n14224);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => n6705, CK => CLK, Q => 
                           n_1753, QN => n14225);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => n6704, CK => CLK, Q => 
                           n_1754, QN => n14226);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => n6703, CK => CLK, Q => 
                           n_1755, QN => n14227);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => n6702, CK => CLK, Q => 
                           n_1756, QN => n14228);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => n6701, CK => CLK, Q => 
                           n_1757, QN => n14229);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => n6700, CK => CLK, Q => 
                           n_1758, QN => n14230);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => n6699, CK => CLK, Q => 
                           n_1759, QN => n14231);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => n6698, CK => CLK, Q => 
                           n_1760, QN => n14232);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => n6697, CK => CLK, Q => 
                           n_1761, QN => n14233);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => n6696, CK => CLK, Q => 
                           n_1762, QN => n14234);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => n6695, CK => CLK, Q => 
                           n_1763, QN => n14235);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => n6694, CK => CLK, Q => 
                           n_1764, QN => n14236);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => n6693, CK => CLK, Q => 
                           n_1765, QN => n14237);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => n6692, CK => CLK, Q => 
                           n_1766, QN => n14238);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => n6691, CK => CLK, Q => 
                           n_1767, QN => n14239);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => n6690, CK => CLK, Q => 
                           n_1768, QN => n14240);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => n6689, CK => CLK, Q => 
                           n_1769, QN => n14241);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => n6688, CK => CLK, Q => 
                           n_1770, QN => n14242);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => n6687, CK => CLK, Q => 
                           n_1771, QN => n14243);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => n6686, CK => CLK, Q => 
                           n_1772, QN => n14244);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n6685, CK => CLK, Q => 
                           n_1773, QN => n14245);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n6684, CK => CLK, Q => 
                           n_1774, QN => n14246);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n6683, CK => CLK, Q => 
                           n_1775, QN => n14247);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n6682, CK => CLK, Q => 
                           n_1776, QN => n14248);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n6681, CK => CLK, Q => 
                           n_1777, QN => n14249);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n6680, CK => CLK, Q => 
                           n_1778, QN => n14250);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n6679, CK => CLK, Q => 
                           n_1779, QN => n14251);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n6678, CK => CLK, Q => 
                           n_1780, QN => n14252);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => n6777, CK => CLK, Q => 
                           n_1781, QN => n14253);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => n6776, CK => CLK, Q => 
                           n_1782, QN => n14254);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => n6775, CK => CLK, Q => 
                           n_1783, QN => n14255);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => n6774, CK => CLK, Q => 
                           n_1784, QN => n14256);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => n6773, CK => CLK, Q => 
                           n_1785, QN => n14257);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => n6772, CK => CLK, Q => 
                           n_1786, QN => n14258);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => n6771, CK => CLK, Q => 
                           n_1787, QN => n14259);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => n6770, CK => CLK, Q => 
                           n_1788, QN => n14260);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => n6769, CK => CLK, Q => 
                           n_1789, QN => n14261);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => n6768, CK => CLK, Q => 
                           n_1790, QN => n14262);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => n6767, CK => CLK, Q => 
                           n_1791, QN => n14263);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => n6766, CK => CLK, Q => 
                           n_1792, QN => n14264);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => n6765, CK => CLK, Q => 
                           n_1793, QN => n14265);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => n6764, CK => CLK, Q => 
                           n_1794, QN => n14266);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => n6763, CK => CLK, Q => 
                           n_1795, QN => n14267);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => n6762, CK => CLK, Q => 
                           n_1796, QN => n14268);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => n6761, CK => CLK, Q => 
                           n_1797, QN => n14269);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => n6760, CK => CLK, Q => 
                           n_1798, QN => n14270);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => n6759, CK => CLK, Q => 
                           n_1799, QN => n14271);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => n6758, CK => CLK, Q => 
                           n_1800, QN => n14272);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => n6757, CK => CLK, Q => 
                           n_1801, QN => n14273);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => n6756, CK => CLK, Q => 
                           n_1802, QN => n14274);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => n6755, CK => CLK, Q => 
                           n_1803, QN => n14275);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => n6754, CK => CLK, Q => 
                           n_1804, QN => n14276);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => n6753, CK => CLK, Q => 
                           n_1805, QN => n14277);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => n6752, CK => CLK, Q => 
                           n_1806, QN => n14278);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => n6751, CK => CLK, Q => 
                           n_1807, QN => n14279);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => n6750, CK => CLK, Q => 
                           n_1808, QN => n14280);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n6749, CK => CLK, Q => 
                           n_1809, QN => n14281);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n6748, CK => CLK, Q => 
                           n_1810, QN => n14282);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n6747, CK => CLK, Q => 
                           n_1811, QN => n14283);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n6746, CK => CLK, Q => 
                           n_1812, QN => n14284);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n6745, CK => CLK, Q => 
                           n_1813, QN => n14285);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n6744, CK => CLK, Q => 
                           n_1814, QN => n14286);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n6743, CK => CLK, Q => 
                           n_1815, QN => n14287);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n6742, CK => CLK, Q => 
                           n_1816, QN => n14288);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n6841, CK => CLK, Q => n9953
                           , QN => n11994);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n6840, CK => CLK, Q => n9954
                           , QN => n11993);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n6839, CK => CLK, Q => n9955
                           , QN => n11992);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n6838, CK => CLK, Q => n9956
                           , QN => n11991);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n6837, CK => CLK, Q => n9957
                           , QN => n11990);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n6836, CK => CLK, Q => n9958
                           , QN => n11989);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n6835, CK => CLK, Q => n9959
                           , QN => n11988);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n6834, CK => CLK, Q => n9960
                           , QN => n11987);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n6833, CK => CLK, Q => n9961
                           , QN => n11986);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n6832, CK => CLK, Q => n9962
                           , QN => n11985);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n6831, CK => CLK, Q => n9963
                           , QN => n11984);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n6830, CK => CLK, Q => n9964
                           , QN => n11983);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n6829, CK => CLK, Q => n9965
                           , QN => n11982);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n6828, CK => CLK, Q => n9966
                           , QN => n11981);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n6827, CK => CLK, Q => n9967
                           , QN => n11980);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n6826, CK => CLK, Q => n9968
                           , QN => n11979);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n6825, CK => CLK, Q => n9969
                           , QN => n11978);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n6824, CK => CLK, Q => n9970
                           , QN => n11977);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n6823, CK => CLK, Q => n9971
                           , QN => n11976);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n6822, CK => CLK, Q => n9972
                           , QN => n11975);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n6821, CK => CLK, Q => n9973
                           , QN => n11974);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n6820, CK => CLK, Q => n9974
                           , QN => n11973);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n6819, CK => CLK, Q => n9975
                           , QN => n11972);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n6818, CK => CLK, Q => n9976
                           , QN => n11971);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n6817, CK => CLK, Q => n9977
                           , QN => n11970);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n6816, CK => CLK, Q => n9978
                           , QN => n11969);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n6815, CK => CLK, Q => n9979
                           , QN => n11968);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n6814, CK => CLK, Q => n9980
                           , QN => n11967);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n6813, CK => CLK, Q => n9981
                           , QN => n11966);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n6812, CK => CLK, Q => n9982
                           , QN => n11965);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n6811, CK => CLK, Q => n9983
                           , QN => n11964);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n6810, CK => CLK, Q => n9984
                           , QN => n11963);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n6809, CK => CLK, Q => n9985
                           , QN => n11962);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n6808, CK => CLK, Q => n9986
                           , QN => n11961);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n6807, CK => CLK, Q => n9987
                           , QN => n11960);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n6806, CK => CLK, Q => n9988
                           , QN => n11959);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n6905, CK => CLK, Q => n9889
                           , QN => n11886);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n6904, CK => CLK, Q => n9890
                           , QN => n11885);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n6903, CK => CLK, Q => n9891
                           , QN => n11884);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n6902, CK => CLK, Q => n9892
                           , QN => n11883);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n6901, CK => CLK, Q => n9893
                           , QN => n11882);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n6900, CK => CLK, Q => n9894
                           , QN => n11881);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n6899, CK => CLK, Q => n9895
                           , QN => n11880);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n6898, CK => CLK, Q => n9896
                           , QN => n11879);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n6897, CK => CLK, Q => n9897
                           , QN => n11878);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n6896, CK => CLK, Q => n9898
                           , QN => n11877);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n6895, CK => CLK, Q => n9899
                           , QN => n11876);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n6894, CK => CLK, Q => n9900
                           , QN => n11875);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n6893, CK => CLK, Q => n9901
                           , QN => n11874);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n6892, CK => CLK, Q => n9902
                           , QN => n11873);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n6891, CK => CLK, Q => n9903
                           , QN => n11872);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n6890, CK => CLK, Q => n9904
                           , QN => n11871);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n6889, CK => CLK, Q => n9905
                           , QN => n11870);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n6888, CK => CLK, Q => n9906
                           , QN => n11869);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n6887, CK => CLK, Q => n9907
                           , QN => n11868);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n6886, CK => CLK, Q => n9908
                           , QN => n11867);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n6885, CK => CLK, Q => n9909
                           , QN => n11866);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n6884, CK => CLK, Q => n9910
                           , QN => n11865);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n6883, CK => CLK, Q => n9911
                           , QN => n11864);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n6882, CK => CLK, Q => n9912
                           , QN => n11863);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n6881, CK => CLK, Q => n9913
                           , QN => n11862);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n6880, CK => CLK, Q => n9914
                           , QN => n11861);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n6879, CK => CLK, Q => n9915
                           , QN => n11860);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n6878, CK => CLK, Q => n9916
                           , QN => n11859);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n6877, CK => CLK, Q => n9917
                           , QN => n11858);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n6876, CK => CLK, Q => n9918
                           , QN => n11857);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n6875, CK => CLK, Q => n9919
                           , QN => n11856);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n6874, CK => CLK, Q => n9920
                           , QN => n11855);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n6873, CK => CLK, Q => n9921
                           , QN => n11854);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n6872, CK => CLK, Q => n9922
                           , QN => n11853);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n6871, CK => CLK, Q => n9923
                           , QN => n11852);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n6870, CK => CLK, Q => n9924
                           , QN => n11851);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n7003, CK => CLK, Q => 
                           n_1817, QN => n14289);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n7002, CK => CLK, Q => 
                           n_1818, QN => n14290);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n7001, CK => CLK, Q => 
                           n_1819, QN => n14291);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n7000, CK => CLK, Q => 
                           n_1820, QN => n14292);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n6999, CK => CLK, Q => 
                           n_1821, QN => n14293);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n6998, CK => CLK, Q => 
                           n_1822, QN => n14294);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n6997, CK => CLK, Q => 
                           n_1823, QN => n14295);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n6996, CK => CLK, Q => 
                           n_1824, QN => n14296);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n6995, CK => CLK, Q => 
                           n_1825, QN => n14297);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n6994, CK => CLK, Q => 
                           n_1826, QN => n14298);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n6993, CK => CLK, Q => 
                           n_1827, QN => n14299);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n6992, CK => CLK, Q => 
                           n_1828, QN => n14300);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n6991, CK => CLK, Q => 
                           n_1829, QN => n14301);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n6990, CK => CLK, Q => 
                           n_1830, QN => n14302);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n6989, CK => CLK, Q => 
                           n_1831, QN => n14303);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n6988, CK => CLK, Q => 
                           n_1832, QN => n14304);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n6987, CK => CLK, Q => 
                           n_1833, QN => n14305);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n6986, CK => CLK, Q => 
                           n_1834, QN => n14306);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n6985, CK => CLK, Q => 
                           n_1835, QN => n14307);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n6984, CK => CLK, Q => 
                           n_1836, QN => n14308);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n6983, CK => CLK, Q => n_1837
                           , QN => n14309);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n6981, CK => CLK, Q => n_1838
                           , QN => n14310);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n6980, CK => CLK, Q => n_1839
                           , QN => n14311);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n6949, CK => CLK, Q => 
                           n_1840, QN => n14312);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n6948, CK => CLK, Q => 
                           n_1841, QN => n14313);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n6947, CK => CLK, Q => 
                           n_1842, QN => n14314);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n6946, CK => CLK, Q => 
                           n_1843, QN => n14315);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n6945, CK => CLK, Q => 
                           n_1844, QN => n14316);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n6944, CK => CLK, Q => 
                           n_1845, QN => n14317);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n6943, CK => CLK, Q => 
                           n_1846, QN => n14318);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n6942, CK => CLK, Q => 
                           n_1847, QN => n14319);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n6941, CK => CLK, Q => 
                           n_1848, QN => n14320);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n6940, CK => CLK, Q => 
                           n_1849, QN => n14321);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n6939, CK => CLK, Q => 
                           n_1850, QN => n14322);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n6982, CK => CLK, Q => n_1851
                           , QN => n14323);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n6979, CK => CLK, Q => n_1852
                           , QN => n14324);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n6978, CK => CLK, Q => n_1853
                           , QN => n14325);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n6977, CK => CLK, Q => n_1854
                           , QN => n14326);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n6976, CK => CLK, Q => n_1855
                           , QN => n14327);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n6975, CK => CLK, Q => n_1856
                           , QN => n14328);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => n6457, CK => CLK, Q => 
                           n11521, QN => n7151);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => n6456, CK => CLK, Q => 
                           n11520, QN => n7248);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => n6455, CK => CLK, Q => 
                           n11519, QN => n7265);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => n6454, CK => CLK, Q => 
                           n11518, QN => n7364);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => n6453, CK => CLK, Q => 
                           n11517, QN => n7381);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => n6452, CK => CLK, Q => 
                           n11516, QN => n7398);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => n6451, CK => CLK, Q => 
                           n11515, QN => n7500);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => n6450, CK => CLK, Q => 
                           n11514, QN => n7517);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => n6449, CK => CLK, Q => 
                           n11513, QN => n7621);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => n6448, CK => CLK, Q => 
                           n11512, QN => n7638);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => n6447, CK => CLK, Q => 
                           n11511, QN => n7655);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => n6446, CK => CLK, Q => 
                           n11510, QN => n7757);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => n6445, CK => CLK, Q => 
                           n11509, QN => n7774);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => n6444, CK => CLK, Q => 
                           n11508, QN => n7791);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => n6443, CK => CLK, Q => 
                           n11507, QN => n7808);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => n6442, CK => CLK, Q => 
                           n11506, QN => n7825);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => n6441, CK => CLK, Q => 
                           n11505, QN => n7842);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => n6440, CK => CLK, Q => 
                           n11504, QN => n7859);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => n6439, CK => CLK, Q => 
                           n11503, QN => n7876);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => n6438, CK => CLK, Q => 
                           n11502, QN => n7893);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => n6437, CK => CLK, Q => 
                           n11501, QN => n7910);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => n6436, CK => CLK, Q => 
                           n11500, QN => n7927);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => n6435, CK => CLK, Q => 
                           n11499, QN => n7944);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => n6434, CK => CLK, Q => 
                           n11498, QN => n7961);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => n6433, CK => CLK, Q => 
                           n11497, QN => n7978);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => n6432, CK => CLK, Q => 
                           n11496, QN => n7995);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => n6431, CK => CLK, Q => 
                           n11495, QN => n8012);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => n6430, CK => CLK, Q => 
                           n11494, QN => n8029);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n6429, CK => CLK, Q => 
                           n11493, QN => n8046);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n6428, CK => CLK, Q => 
                           n11492, QN => n8063);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n6427, CK => CLK, Q => 
                           n11491, QN => n8080);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n6426, CK => CLK, Q => 
                           n11490, QN => n8097);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n6425, CK => CLK, Q => 
                           n11489, QN => n8114);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n6424, CK => CLK, Q => 
                           n11488, QN => n8131);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n6423, CK => CLK, Q => 
                           n11487, QN => n8148);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n6422, CK => CLK, Q => 
                           n11486, QN => n8165);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => n6521, CK => CLK, Q => 
                           n11701, QN => n7152);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => n6520, CK => CLK, Q => 
                           n11700, QN => n7249);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => n6519, CK => CLK, Q => 
                           n11699, QN => n7266);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => n6518, CK => CLK, Q => 
                           n11698, QN => n7365);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => n6517, CK => CLK, Q => 
                           n11697, QN => n7382);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => n6516, CK => CLK, Q => 
                           n11696, QN => n7399);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => n6515, CK => CLK, Q => 
                           n11695, QN => n7501);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => n6514, CK => CLK, Q => 
                           n11694, QN => n7518);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => n6513, CK => CLK, Q => 
                           n11693, QN => n7622);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => n6512, CK => CLK, Q => 
                           n11692, QN => n7639);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => n6511, CK => CLK, Q => 
                           n11691, QN => n7656);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => n6510, CK => CLK, Q => 
                           n11690, QN => n7758);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => n6509, CK => CLK, Q => 
                           n11689, QN => n7775);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => n6508, CK => CLK, Q => 
                           n11688, QN => n7792);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => n6507, CK => CLK, Q => 
                           n11687, QN => n7809);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => n6506, CK => CLK, Q => 
                           n11686, QN => n7826);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => n6505, CK => CLK, Q => 
                           n11685, QN => n7843);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => n6504, CK => CLK, Q => 
                           n11684, QN => n7860);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => n6503, CK => CLK, Q => 
                           n11683, QN => n7877);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => n6502, CK => CLK, Q => 
                           n11682, QN => n7894);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => n6501, CK => CLK, Q => 
                           n11681, QN => n7911);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => n6500, CK => CLK, Q => 
                           n11680, QN => n7928);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => n6499, CK => CLK, Q => 
                           n11679, QN => n7945);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => n6498, CK => CLK, Q => 
                           n11678, QN => n7962);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => n6497, CK => CLK, Q => 
                           n11677, QN => n7979);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => n6496, CK => CLK, Q => 
                           n11676, QN => n7996);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => n6495, CK => CLK, Q => 
                           n11675, QN => n8013);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => n6494, CK => CLK, Q => 
                           n11674, QN => n8030);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n6493, CK => CLK, Q => 
                           n11673, QN => n8047);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n6492, CK => CLK, Q => 
                           n11672, QN => n8064);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n6491, CK => CLK, Q => 
                           n11671, QN => n8081);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n6490, CK => CLK, Q => 
                           n11670, QN => n8098);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n6489, CK => CLK, Q => 
                           n11669, QN => n8115);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n6488, CK => CLK, Q => 
                           n11668, QN => n8132);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n6487, CK => CLK, Q => 
                           n11667, QN => n8149);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n6486, CK => CLK, Q => 
                           n11666, QN => n8166);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => n6265, CK => CLK, Q => 
                           n11761, QN => n7234);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => n6264, CK => CLK, Q => 
                           n11760, QN => n7251);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => n6263, CK => CLK, Q => 
                           n11759, QN => n7268);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => n6262, CK => CLK, Q => 
                           n11758, QN => n7367);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => n6261, CK => CLK, Q => 
                           n11757, QN => n7384);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => n6260, CK => CLK, Q => 
                           n11756, QN => n7401);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => n6259, CK => CLK, Q => 
                           n11755, QN => n7503);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => n6258, CK => CLK, Q => 
                           n11754, QN => n7520);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => n6257, CK => CLK, Q => 
                           n11753, QN => n7624);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => n6256, CK => CLK, Q => 
                           n11752, QN => n7641);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => n6255, CK => CLK, Q => 
                           n11751, QN => n7743);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => n6254, CK => CLK, Q => 
                           n11750, QN => n7760);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => n6253, CK => CLK, Q => 
                           n11749, QN => n7777);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => n6252, CK => CLK, Q => 
                           n11748, QN => n7794);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => n6251, CK => CLK, Q => 
                           n11747, QN => n7811);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => n6250, CK => CLK, Q => 
                           n11746, QN => n7828);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => n6249, CK => CLK, Q => 
                           n11745, QN => n7845);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => n6248, CK => CLK, Q => 
                           n11744, QN => n7862);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => n6247, CK => CLK, Q => 
                           n11743, QN => n7879);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => n6246, CK => CLK, Q => 
                           n11742, QN => n7896);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => n6245, CK => CLK, Q => 
                           n11741, QN => n7913);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => n6244, CK => CLK, Q => 
                           n11740, QN => n7930);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => n6243, CK => CLK, Q => 
                           n11739, QN => n7947);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => n6242, CK => CLK, Q => 
                           n11738, QN => n7964);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => n6241, CK => CLK, Q => 
                           n11737, QN => n7981);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => n6240, CK => CLK, Q => 
                           n11736, QN => n7998);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => n6239, CK => CLK, Q => 
                           n11735, QN => n8015);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => n6238, CK => CLK, Q => 
                           n11734, QN => n8032);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n6237, CK => CLK, Q => 
                           n11733, QN => n8049);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n6236, CK => CLK, Q => 
                           n11732, QN => n8066);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n6235, CK => CLK, Q => 
                           n11731, QN => n8083);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n6234, CK => CLK, Q => 
                           n11730, QN => n8100);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n6233, CK => CLK, Q => 
                           n11729, QN => n8117);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n6232, CK => CLK, Q => 
                           n11728, QN => n8134);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n6231, CK => CLK, Q => 
                           n11727, QN => n8151);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n6230, CK => CLK, Q => 
                           n11726, QN => n8168);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => n6201, CK => CLK, Q => 
                           n11581, QN => n7153);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => n6200, CK => CLK, Q => 
                           n11580, QN => n7250);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => n6199, CK => CLK, Q => 
                           n11579, QN => n7267);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => n6198, CK => CLK, Q => 
                           n11578, QN => n7366);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => n6197, CK => CLK, Q => 
                           n11577, QN => n7383);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => n6196, CK => CLK, Q => 
                           n11576, QN => n7400);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => n6195, CK => CLK, Q => 
                           n11575, QN => n7502);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => n6194, CK => CLK, Q => 
                           n11574, QN => n7519);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => n6193, CK => CLK, Q => 
                           n11573, QN => n7623);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => n6192, CK => CLK, Q => 
                           n11572, QN => n7640);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => n6191, CK => CLK, Q => 
                           n11571, QN => n7742);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => n6190, CK => CLK, Q => 
                           n11570, QN => n7759);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => n6189, CK => CLK, Q => 
                           n11569, QN => n7776);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => n6188, CK => CLK, Q => 
                           n11568, QN => n7793);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => n6187, CK => CLK, Q => 
                           n11567, QN => n7810);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => n6186, CK => CLK, Q => 
                           n11566, QN => n7827);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => n6185, CK => CLK, Q => 
                           n11565, QN => n7844);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => n6184, CK => CLK, Q => 
                           n11564, QN => n7861);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => n6183, CK => CLK, Q => 
                           n11563, QN => n7878);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => n6182, CK => CLK, Q => 
                           n11562, QN => n7895);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => n6181, CK => CLK, Q => 
                           n11561, QN => n7912);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => n6180, CK => CLK, Q => 
                           n11560, QN => n7929);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => n6179, CK => CLK, Q => 
                           n11559, QN => n7946);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => n6178, CK => CLK, Q => 
                           n11558, QN => n7963);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => n6177, CK => CLK, Q => 
                           n11557, QN => n7980);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => n6176, CK => CLK, Q => 
                           n11556, QN => n7997);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => n6175, CK => CLK, Q => 
                           n11555, QN => n8014);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => n6174, CK => CLK, Q => 
                           n11554, QN => n8031);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n6173, CK => CLK, Q => 
                           n11553, QN => n8048);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n6172, CK => CLK, Q => 
                           n11552, QN => n8065);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n6171, CK => CLK, Q => 
                           n11551, QN => n8082);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n6170, CK => CLK, Q => 
                           n11550, QN => n8099);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n6169, CK => CLK, Q => 
                           n11549, QN => n8116);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n6168, CK => CLK, Q => 
                           n11548, QN => n8133);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n6167, CK => CLK, Q => 
                           n11547, QN => n8150);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n6166, CK => CLK, Q => 
                           n11546, QN => n8167);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n6289, CK => CLK, Q => 
                           n_1857, QN => n14329);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n6288, CK => CLK, Q => 
                           n_1858, QN => n14330);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n6287, CK => CLK, Q => 
                           n_1859, QN => n14331);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n6285, CK => CLK, Q => 
                           n_1860, QN => n14332);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n6284, CK => CLK, Q => 
                           n_1861, QN => n14333);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n6283, CK => CLK, Q => 
                           n_1862, QN => n14334);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n6282, CK => CLK, Q => 
                           n_1863, QN => n14335);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n6281, CK => CLK, Q => 
                           n_1864, QN => n14336);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n6280, CK => CLK, Q => 
                           n_1865, QN => n14337);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n6279, CK => CLK, Q => 
                           n_1866, QN => n14338);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n6278, CK => CLK, Q => 
                           n_1867, QN => n14339);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n6277, CK => CLK, Q => 
                           n_1868, QN => n14340);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n6035, CK => CLK, Q => 
                           n_1869, QN => n14341);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n6034, CK => CLK, Q => 
                           n_1870, QN => n14342);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n6033, CK => CLK, Q => 
                           n_1871, QN => n14343);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n6032, CK => CLK, Q => 
                           n_1872, QN => n14344);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n6031, CK => CLK, Q => 
                           n_1873, QN => n14345);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n6029, CK => CLK, Q => 
                           n_1874, QN => n14346);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n6028, CK => CLK, Q => 
                           n_1875, QN => n14347);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n6027, CK => CLK, Q => 
                           n_1876, QN => n14348);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n6026, CK => CLK, Q => 
                           n_1877, QN => n14349);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n6025, CK => CLK, Q => 
                           n_1878, QN => n14350);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n6024, CK => CLK, Q => 
                           n_1879, QN => n14351);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n6023, CK => CLK, Q => 
                           n_1880, QN => n14352);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n6022, CK => CLK, Q => 
                           n_1881, QN => n14353);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n6021, CK => CLK, Q => 
                           n_1882, QN => n14354);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n6020, CK => CLK, Q => 
                           n_1883, QN => n14355);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n6019, CK => CLK, Q => 
                           n_1884, QN => n14356);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n6018, CK => CLK, Q => 
                           n_1885, QN => n14357);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n6276, CK => CLK, Q => 
                           n_1886, QN => n14358);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n6275, CK => CLK, Q => 
                           n_1887, QN => n14359);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n6274, CK => CLK, Q => 
                           n_1888, QN => n14360);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n6526, CK => CLK, Q => n11586
                           , QN => n8572);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n6590, CK => CLK, Q => n11406
                           , QN => n8571);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n6654, CK => CLK, Q => n_1889
                           , QN => n14361);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n6718, CK => CLK, Q => n_1890
                           , QN => n14362);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n6782, CK => CLK, Q => n11766
                           , QN => n8570);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n6846, CK => CLK, Q => n9948,
                           QN => n11802);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n6549, CK => CLK, Q => 
                           n11606, QN => n8181);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n6548, CK => CLK, Q => 
                           n11605, QN => n8198);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n6547, CK => CLK, Q => 
                           n11604, QN => n8215);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n6546, CK => CLK, Q => 
                           n11603, QN => n8232);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n6545, CK => CLK, Q => 
                           n11602, QN => n8249);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n6544, CK => CLK, Q => 
                           n11601, QN => n8266);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n6543, CK => CLK, Q => 
                           n11600, QN => n8283);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n6542, CK => CLK, Q => 
                           n11599, QN => n8300);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n6541, CK => CLK, Q => 
                           n11598, QN => n8317);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n6540, CK => CLK, Q => 
                           n11597, QN => n8334);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n6539, CK => CLK, Q => 
                           n11596, QN => n8351);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n6538, CK => CLK, Q => 
                           n11595, QN => n8368);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n6537, CK => CLK, Q => 
                           n11594, QN => n8385);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n6536, CK => CLK, Q => 
                           n11593, QN => n8402);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n6535, CK => CLK, Q => n11592
                           , QN => n8419);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n6534, CK => CLK, Q => n11591
                           , QN => n8436);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n6533, CK => CLK, Q => n11590
                           , QN => n8453);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n6532, CK => CLK, Q => n11764
                           , QN => n8470);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n6531, CK => CLK, Q => n11763
                           , QN => n8487);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n6530, CK => CLK, Q => n11589
                           , QN => n8504);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n6529, CK => CLK, Q => n11588
                           , QN => n8521);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n6528, CK => CLK, Q => n11587
                           , QN => n8538);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n6527, CK => CLK, Q => n11762
                           , QN => n8555);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n6613, CK => CLK, Q => 
                           n11426, QN => n8180);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n6612, CK => CLK, Q => 
                           n11425, QN => n8197);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n6611, CK => CLK, Q => 
                           n11424, QN => n8214);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n6610, CK => CLK, Q => 
                           n11423, QN => n8231);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n6609, CK => CLK, Q => 
                           n11422, QN => n8248);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n6608, CK => CLK, Q => 
                           n11421, QN => n8265);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n6607, CK => CLK, Q => 
                           n11420, QN => n8282);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n6606, CK => CLK, Q => 
                           n11419, QN => n8299);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n6605, CK => CLK, Q => 
                           n11418, QN => n8316);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n6604, CK => CLK, Q => 
                           n11417, QN => n8333);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n6603, CK => CLK, Q => 
                           n11416, QN => n8350);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n6602, CK => CLK, Q => 
                           n11415, QN => n8367);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n6601, CK => CLK, Q => 
                           n11414, QN => n8384);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n6600, CK => CLK, Q => 
                           n11413, QN => n8401);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n6599, CK => CLK, Q => n11412
                           , QN => n8418);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n6598, CK => CLK, Q => n11411
                           , QN => n8435);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n6597, CK => CLK, Q => n11410
                           , QN => n8452);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n6596, CK => CLK, Q => n11584
                           , QN => n8469);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n6595, CK => CLK, Q => n11583
                           , QN => n8486);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n6594, CK => CLK, Q => n11409
                           , QN => n8503);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n6593, CK => CLK, Q => n11408
                           , QN => n8520);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n6592, CK => CLK, Q => n11407
                           , QN => n8537);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n6591, CK => CLK, Q => n11582
                           , QN => n8554);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n6677, CK => CLK, Q => 
                           n_1891, QN => n14363);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n6676, CK => CLK, Q => 
                           n_1892, QN => n14364);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n6675, CK => CLK, Q => 
                           n_1893, QN => n14365);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n6674, CK => CLK, Q => 
                           n_1894, QN => n14366);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n6673, CK => CLK, Q => 
                           n_1895, QN => n14367);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n6672, CK => CLK, Q => 
                           n_1896, QN => n14368);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n6671, CK => CLK, Q => 
                           n_1897, QN => n14369);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n6670, CK => CLK, Q => 
                           n_1898, QN => n14370);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n6669, CK => CLK, Q => 
                           n_1899, QN => n14371);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n6668, CK => CLK, Q => 
                           n_1900, QN => n14372);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n6667, CK => CLK, Q => 
                           n_1901, QN => n14373);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n6666, CK => CLK, Q => 
                           n_1902, QN => n14374);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n6665, CK => CLK, Q => 
                           n_1903, QN => n14375);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n6664, CK => CLK, Q => 
                           n_1904, QN => n14376);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n6663, CK => CLK, Q => n_1905
                           , QN => n14377);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n6662, CK => CLK, Q => n_1906
                           , QN => n14378);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n6661, CK => CLK, Q => n_1907
                           , QN => n14379);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n6660, CK => CLK, Q => n_1908
                           , QN => n14380);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n6659, CK => CLK, Q => n_1909
                           , QN => n14381);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n6658, CK => CLK, Q => n_1910
                           , QN => n14382);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n6657, CK => CLK, Q => n_1911
                           , QN => n14383);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n6656, CK => CLK, Q => n_1912
                           , QN => n14384);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n6655, CK => CLK, Q => n_1913
                           , QN => n14385);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n6741, CK => CLK, Q => 
                           n_1914, QN => n14386);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n6740, CK => CLK, Q => 
                           n_1915, QN => n14387);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n6739, CK => CLK, Q => 
                           n_1916, QN => n14388);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n6738, CK => CLK, Q => 
                           n_1917, QN => n14389);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n6737, CK => CLK, Q => 
                           n_1918, QN => n14390);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n6736, CK => CLK, Q => 
                           n_1919, QN => n14391);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n6735, CK => CLK, Q => 
                           n_1920, QN => n14392);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n6734, CK => CLK, Q => 
                           n_1921, QN => n14393);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n6733, CK => CLK, Q => 
                           n_1922, QN => n14394);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n6732, CK => CLK, Q => 
                           n_1923, QN => n14395);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n6731, CK => CLK, Q => 
                           n_1924, QN => n14396);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n6730, CK => CLK, Q => 
                           n_1925, QN => n14397);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n6729, CK => CLK, Q => 
                           n_1926, QN => n14398);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n6728, CK => CLK, Q => 
                           n_1927, QN => n14399);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n6727, CK => CLK, Q => n_1928
                           , QN => n14400);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n6726, CK => CLK, Q => n_1929
                           , QN => n14401);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n6725, CK => CLK, Q => n_1930
                           , QN => n14402);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n6724, CK => CLK, Q => n_1931
                           , QN => n14403);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n6723, CK => CLK, Q => n_1932
                           , QN => n14404);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n6722, CK => CLK, Q => n_1933
                           , QN => n14405);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n6721, CK => CLK, Q => n_1934
                           , QN => n14406);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n6720, CK => CLK, Q => n_1935
                           , QN => n14407);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n6719, CK => CLK, Q => n_1936
                           , QN => n14408);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n6805, CK => CLK, Q => n9989
                           , QN => n12056);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n6804, CK => CLK, Q => n9990
                           , QN => n12055);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n6803, CK => CLK, Q => n9991
                           , QN => n12054);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n6802, CK => CLK, Q => n9992
                           , QN => n12053);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n6801, CK => CLK, Q => n9993
                           , QN => n12052);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n6800, CK => CLK, Q => n9994
                           , QN => n12051);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n6799, CK => CLK, Q => n9995
                           , QN => n12050);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n6798, CK => CLK, Q => n9996
                           , QN => n12049);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n6797, CK => CLK, Q => n9997
                           , QN => n12048);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n6796, CK => CLK, Q => n9998
                           , QN => n12047);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n6795, CK => CLK, Q => n9999
                           , QN => n12046);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n6794, CK => CLK, Q => 
                           n11778, QN => n8366);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n6793, CK => CLK, Q => 
                           n11777, QN => n8383);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n6792, CK => CLK, Q => 
                           n11776, QN => n8400);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n6791, CK => CLK, Q => n11775
                           , QN => n8417);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n6790, CK => CLK, Q => n11774
                           , QN => n8434);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n6789, CK => CLK, Q => n11773
                           , QN => n8451);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n6788, CK => CLK, Q => n11772
                           , QN => n8468);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n6787, CK => CLK, Q => n11771
                           , QN => n8485);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n6786, CK => CLK, Q => n11770
                           , QN => n8502);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n6785, CK => CLK, Q => n11769
                           , QN => n8519);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n6784, CK => CLK, Q => n11768
                           , QN => n8536);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n6783, CK => CLK, Q => n11767
                           , QN => n8553);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n6869, CK => CLK, Q => n9925
                           , QN => n11801);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n6868, CK => CLK, Q => n9926
                           , QN => n11800);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n6867, CK => CLK, Q => n9927
                           , QN => n11799);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n6866, CK => CLK, Q => n9928
                           , QN => n11798);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n6865, CK => CLK, Q => n9929
                           , QN => n11797);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n6864, CK => CLK, Q => n9930
                           , QN => n11796);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n6863, CK => CLK, Q => n9931
                           , QN => n11795);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n6862, CK => CLK, Q => n9932
                           , QN => n11794);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n6861, CK => CLK, Q => n9933
                           , QN => n11793);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n6860, CK => CLK, Q => n9934
                           , QN => n11792);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n6859, CK => CLK, Q => n9935
                           , QN => n11791);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n6858, CK => CLK, Q => n9936
                           , QN => n11790);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n6857, CK => CLK, Q => n9937
                           , QN => n11789);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n6856, CK => CLK, Q => n9938
                           , QN => n11788);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n6855, CK => CLK, Q => n9939,
                           QN => n11787);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n6854, CK => CLK, Q => n9940,
                           QN => n11786);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n6853, CK => CLK, Q => n9941,
                           QN => n11785);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n6852, CK => CLK, Q => n9942,
                           QN => n11784);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n6851, CK => CLK, Q => n9943,
                           QN => n11783);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n6850, CK => CLK, Q => n9944,
                           QN => n11782);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n6849, CK => CLK, Q => n9945,
                           QN => n11781);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n6848, CK => CLK, Q => n9946,
                           QN => n11780);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n6847, CK => CLK, Q => n9947,
                           QN => n11779);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n6970, CK => CLK, Q => 
                           n_1937, QN => n14412);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n6969, CK => CLK, Q => 
                           n_1938, QN => n14413);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n6968, CK => CLK, Q => 
                           n_1939, QN => n14414);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n6967, CK => CLK, Q => 
                           n_1940, QN => n14415);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n6966, CK => CLK, Q => 
                           n_1941, QN => n14416);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n6965, CK => CLK, Q => 
                           n_1942, QN => n14417);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n6964, CK => CLK, Q => 
                           n_1943, QN => n14418);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n6963, CK => CLK, Q => 
                           n_1944, QN => n14419);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n6962, CK => CLK, Q => 
                           n_1945, QN => n14420);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n6961, CK => CLK, Q => 
                           n_1946, QN => n14421);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n6960, CK => CLK, Q => 
                           n_1947, QN => n14422);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n6959, CK => CLK, Q => 
                           n_1948, QN => n14423);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n6958, CK => CLK, Q => 
                           n_1949, QN => n14424);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n6957, CK => CLK, Q => 
                           n_1950, QN => n14425);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n6956, CK => CLK, Q => 
                           n_1951, QN => n14426);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n6955, CK => CLK, Q => 
                           n_1952, QN => n14427);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n6954, CK => CLK, Q => 
                           n_1953, QN => n14428);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n6953, CK => CLK, Q => 
                           n_1954, QN => n14429);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n6952, CK => CLK, Q => 
                           n_1955, QN => n14430);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n6951, CK => CLK, Q => 
                           n_1956, QN => n14431);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n6950, CK => CLK, Q => 
                           n_1957, QN => n14432);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n7036, CK => CLK, Q => 
                           n_1958, QN => n14433);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n7035, CK => CLK, Q => 
                           n_1959, QN => n14434);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n7034, CK => CLK, Q => 
                           n_1960, QN => n14435);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n7033, CK => CLK, Q => 
                           n_1961, QN => n14436);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n7032, CK => CLK, Q => 
                           n_1962, QN => n14437);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n7031, CK => CLK, Q => 
                           n_1963, QN => n14438);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n7030, CK => CLK, Q => 
                           n_1964, QN => n14439);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n7029, CK => CLK, Q => 
                           n_1965, QN => n14440);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n7019, CK => CLK, Q => 
                           n_1966, QN => n14441);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n7018, CK => CLK, Q => 
                           n_1967, QN => n14442);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n7017, CK => CLK, Q => 
                           n_1968, QN => n14443);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n7016, CK => CLK, Q => 
                           n_1969, QN => n14444);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n7015, CK => CLK, Q => 
                           n_1970, QN => n14445);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n7014, CK => CLK, Q => 
                           n_1971, QN => n14446);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n7013, CK => CLK, Q => 
                           n_1972, QN => n14447);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n7012, CK => CLK, Q => 
                           n_1973, QN => n14448);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n7011, CK => CLK, Q => 
                           n_1974, QN => n14449);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n7010, CK => CLK, Q => 
                           n_1975, QN => n14450);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n7009, CK => CLK, Q => 
                           n_1976, QN => n14451);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n7008, CK => CLK, Q => 
                           n_1977, QN => n14452);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n7007, CK => CLK, Q => 
                           n_1978, QN => n14453);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n7006, CK => CLK, Q => 
                           n_1979, QN => n14454);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n7005, CK => CLK, Q => 
                           n_1980, QN => n14455);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n7004, CK => CLK, Q => 
                           n_1981, QN => n14456);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n6421, CK => CLK, Q => 
                           n11485, QN => n8182);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n6420, CK => CLK, Q => 
                           n11484, QN => n8199);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n6419, CK => CLK, Q => 
                           n11483, QN => n8216);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n6418, CK => CLK, Q => 
                           n11482, QN => n8233);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n6417, CK => CLK, Q => 
                           n11481, QN => n8250);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n6416, CK => CLK, Q => 
                           n11480, QN => n8267);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n6415, CK => CLK, Q => 
                           n11479, QN => n8284);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n6414, CK => CLK, Q => 
                           n11478, QN => n8301);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n6413, CK => CLK, Q => 
                           n11477, QN => n8318);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n6412, CK => CLK, Q => 
                           n11476, QN => n8335);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n6411, CK => CLK, Q => 
                           n11475, QN => n8352);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n6410, CK => CLK, Q => 
                           n11474, QN => n8369);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n6409, CK => CLK, Q => 
                           n11473, QN => n8386);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n6408, CK => CLK, Q => 
                           n11472, QN => n8403);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n6407, CK => CLK, Q => n11471
                           , QN => n8420);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n6406, CK => CLK, Q => n11470
                           , QN => n8437);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n6405, CK => CLK, Q => n11469
                           , QN => n8454);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n6404, CK => CLK, Q => n11468
                           , QN => n8471);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n6403, CK => CLK, Q => n11467
                           , QN => n8488);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n6402, CK => CLK, Q => n11466
                           , QN => n8505);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n6401, CK => CLK, Q => n11465
                           , QN => n8522);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n6400, CK => CLK, Q => n11464
                           , QN => n8539);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n6399, CK => CLK, Q => n11463
                           , QN => n8556);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n6398, CK => CLK, Q => n11462
                           , QN => n8573);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n6485, CK => CLK, Q => 
                           n11665, QN => n8183);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n6484, CK => CLK, Q => 
                           n11664, QN => n8200);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n6483, CK => CLK, Q => 
                           n11663, QN => n8217);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n6482, CK => CLK, Q => 
                           n11662, QN => n8234);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n6481, CK => CLK, Q => 
                           n11661, QN => n8251);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n6480, CK => CLK, Q => 
                           n11660, QN => n8268);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n6479, CK => CLK, Q => 
                           n11659, QN => n8285);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n6478, CK => CLK, Q => 
                           n11658, QN => n8302);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n6477, CK => CLK, Q => 
                           n11657, QN => n8319);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n6476, CK => CLK, Q => 
                           n11656, QN => n8336);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n6475, CK => CLK, Q => 
                           n11655, QN => n8353);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n6474, CK => CLK, Q => 
                           n11654, QN => n8370);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n6473, CK => CLK, Q => 
                           n11653, QN => n8387);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n6472, CK => CLK, Q => 
                           n11652, QN => n8404);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n6471, CK => CLK, Q => n11651
                           , QN => n8421);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n6470, CK => CLK, Q => n11650
                           , QN => n8438);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n6469, CK => CLK, Q => n11649
                           , QN => n8455);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n6468, CK => CLK, Q => n11648
                           , QN => n8472);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n6467, CK => CLK, Q => n11647
                           , QN => n8489);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n6466, CK => CLK, Q => n11646
                           , QN => n8506);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n6465, CK => CLK, Q => n11645
                           , QN => n8523);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n6464, CK => CLK, Q => n11644
                           , QN => n8540);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n6463, CK => CLK, Q => n11643
                           , QN => n8557);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n6462, CK => CLK, Q => n11642
                           , QN => n8574);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n6229, CK => CLK, Q => 
                           n11725, QN => n8185);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n6228, CK => CLK, Q => 
                           n11724, QN => n8202);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n6227, CK => CLK, Q => 
                           n11723, QN => n8219);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n6226, CK => CLK, Q => 
                           n11722, QN => n8236);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n6225, CK => CLK, Q => 
                           n11721, QN => n8253);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n6224, CK => CLK, Q => 
                           n11720, QN => n8270);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n6223, CK => CLK, Q => 
                           n11719, QN => n8287);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n6222, CK => CLK, Q => 
                           n11718, QN => n8304);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n6221, CK => CLK, Q => 
                           n11717, QN => n8321);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n6220, CK => CLK, Q => 
                           n11716, QN => n8338);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n6219, CK => CLK, Q => 
                           n11715, QN => n8355);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n6218, CK => CLK, Q => 
                           n11714, QN => n8372);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n6217, CK => CLK, Q => 
                           n11713, QN => n8389);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n6216, CK => CLK, Q => 
                           n11712, QN => n8406);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n6215, CK => CLK, Q => 
                           n11711, QN => n8423);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n6214, CK => CLK, Q => 
                           n11710, QN => n8440);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n6213, CK => CLK, Q => 
                           n11709, QN => n8457);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n6212, CK => CLK, Q => 
                           n11708, QN => n8474);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n6211, CK => CLK, Q => 
                           n11707, QN => n8491);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n6210, CK => CLK, Q => 
                           n11706, QN => n8508);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n6209, CK => CLK, Q => 
                           n11705, QN => n8525);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n6208, CK => CLK, Q => 
                           n11704, QN => n8542);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n6207, CK => CLK, Q => 
                           n11703, QN => n8559);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n6206, CK => CLK, Q => 
                           n11702, QN => n8576);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n6165, CK => CLK, Q => 
                           n11545, QN => n8184);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n6164, CK => CLK, Q => 
                           n11544, QN => n8201);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n6163, CK => CLK, Q => 
                           n11543, QN => n8218);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n6162, CK => CLK, Q => 
                           n11542, QN => n8235);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n6161, CK => CLK, Q => 
                           n11541, QN => n8252);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n6160, CK => CLK, Q => 
                           n11540, QN => n8269);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n6159, CK => CLK, Q => 
                           n11539, QN => n8286);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n6158, CK => CLK, Q => 
                           n11538, QN => n8303);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n6157, CK => CLK, Q => 
                           n11537, QN => n8320);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n6156, CK => CLK, Q => 
                           n11536, QN => n8337);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n6155, CK => CLK, Q => 
                           n11535, QN => n8354);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n6154, CK => CLK, Q => 
                           n11534, QN => n8371);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n6153, CK => CLK, Q => 
                           n11533, QN => n8388);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n6152, CK => CLK, Q => 
                           n11532, QN => n8405);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n6151, CK => CLK, Q => 
                           n11531, QN => n8422);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n6150, CK => CLK, Q => 
                           n11530, QN => n8439);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n6149, CK => CLK, Q => 
                           n11529, QN => n8456);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n6148, CK => CLK, Q => 
                           n11528, QN => n8473);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n6147, CK => CLK, Q => 
                           n11527, QN => n8490);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n6146, CK => CLK, Q => 
                           n11526, QN => n8507);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n6145, CK => CLK, Q => 
                           n11525, QN => n8524);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n6144, CK => CLK, Q => 
                           n11524, QN => n8541);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n6143, CK => CLK, Q => 
                           n11523, QN => n8558);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n6142, CK => CLK, Q => 
                           n11522, QN => n8575);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => n6312, CK => CLK, Q => 
                           n_1982, QN => n14457);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => n6311, CK => CLK, Q => 
                           n_1983, QN => n14458);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => n6310, CK => CLK, Q => 
                           n_1984, QN => n14459);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => n6309, CK => CLK, Q => 
                           n_1985, QN => n14460);
   U6638 : NAND3_X1 port map( A1 => n13383, A2 => n13382, A3 => n1922, ZN => 
                           n1906);
   U6640 : NAND3_X1 port map( A1 => n1922, A2 => n13383, A3 => ADD_WR(4), ZN =>
                           n1933);
   U6641 : NAND3_X1 port map( A1 => n13385, A2 => n13384, A3 => n13386, ZN => 
                           n1907);
   U6642 : NAND3_X1 port map( A1 => n13385, A2 => n13384, A3 => ADD_WR(0), ZN 
                           => n1909);
   U6643 : NAND3_X1 port map( A1 => n13386, A2 => n13384, A3 => ADD_WR(1), ZN 
                           => n1911);
   U6644 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n13384, A3 => ADD_WR(1), 
                           ZN => n1913);
   U6645 : NAND3_X1 port map( A1 => n13386, A2 => n13385, A3 => ADD_WR(2), ZN 
                           => n1915);
   U6646 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n13385, A3 => ADD_WR(2), 
                           ZN => n1917);
   U6647 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n13386, A3 => ADD_WR(2), 
                           ZN => n1919);
   U6649 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n1921);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => n5437, CK => CLK, Q => 
                           n_1986, QN => n13731);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => n5436, CK => CLK, Q => 
                           n_1987, QN => n13732);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => n5435, CK => CLK, Q => 
                           n_1988, QN => n13733);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => n5434, CK => CLK, Q => 
                           n_1989, QN => n13734);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => n5501, CK => CLK, Q => 
                           n_1990, QN => n13667);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => n5500, CK => CLK, Q => 
                           n_1991, QN => n13668);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => n5499, CK => CLK, Q => 
                           n_1992, QN => n13669);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => n5498, CK => CLK, Q => 
                           n_1993, QN => n13670);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => n5245, CK => CLK, Q => 
                           n_1994, QN => n13747);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => n5244, CK => CLK, Q => 
                           n_1995, QN => n13748);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => n5243, CK => CLK, Q => 
                           n_1996, QN => n13749);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => n5242, CK => CLK, Q => 
                           n_1997, QN => n13750);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => n5181, CK => CLK, Q => 
                           n_1998, QN => n14083);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => n5180, CK => CLK, Q => 
                           n_1999, QN => n14084);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => n5179, CK => CLK, Q => 
                           n_2000, QN => n14085);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => n5178, CK => CLK, Q => 
                           n_2001, QN => n14086);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => n5565, CK => CLK, Q => 
                           n4511, QN => n13663);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => n5564, CK => CLK, Q => 
                           n4509, QN => n13664);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => n5563, CK => CLK, Q => 
                           n4507, QN => n13665);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => n5562, CK => CLK, Q => 
                           n4505, QN => n13666);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => n5629, CK => CLK, Q => 
                           n4510, QN => n13659);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => n5628, CK => CLK, Q => 
                           n4508, QN => n13660);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => n5627, CK => CLK, Q => 
                           n4506, QN => n13661);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => n5626, CK => CLK, Q => 
                           n4504, QN => n13662);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => n5821, CK => CLK, Q => 
                           n4479, QN => n13655);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => n5820, CK => CLK, Q => 
                           n4477, QN => n13656);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => n5819, CK => CLK, Q => 
                           n4475, QN => n13657);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => n5818, CK => CLK, Q => 
                           n4473, QN => n13658);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => n5885, CK => CLK, Q => 
                           n4478, QN => n13651);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => n5884, CK => CLK, Q => 
                           n4476, QN => n13652);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => n5883, CK => CLK, Q => 
                           n4474, QN => n13653);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => n5882, CK => CLK, Q => 
                           n4472, QN => n13654);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n6845, CK => CLK, Q => n9949
                           , QN => n13848);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => n6397, CK => CLK, Q => 
                           n_2002, QN => n13431);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => n6396, CK => CLK, Q => 
                           n_2003, QN => n13432);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => n6395, CK => CLK, Q => 
                           n_2004, QN => n13433);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => n6394, CK => CLK, Q => 
                           n_2005, QN => n13434);
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => n6333, CK => CLK, Q => 
                           n_2006, QN => n13495);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => n6332, CK => CLK, Q => 
                           n_2007, QN => n13496);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => n6331, CK => CLK, Q => 
                           n_2008, QN => n13497);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => n6330, CK => CLK, Q => 
                           n_2009, QN => n13498);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => n6077, CK => CLK, Q => 
                           n_2010, QN => n13604);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => n6076, CK => CLK, Q => 
                           n_2011, QN => n13605);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => n6075, CK => CLK, Q => 
                           n_2012, QN => n13606);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => n6074, CK => CLK, Q => 
                           n_2013, QN => n13607);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => n6141, CK => CLK, Q => 
                           n_2014, QN => n13540);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => n6140, CK => CLK, Q => 
                           n_2015, QN => n13541);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => n6139, CK => CLK, Q => 
                           n_2016, QN => n13542);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => n6138, CK => CLK, Q => 
                           n_2017, QN => n13543);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => n6717, CK => CLK, Q => 
                           n_2018, QN => n13840);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => n6716, CK => CLK, Q => 
                           n_2019, QN => n13841);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => n6715, CK => CLK, Q => 
                           n_2020, QN => n13842);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => n6714, CK => CLK, Q => 
                           n_2021, QN => n13843);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => n6781, CK => CLK, Q => 
                           n_2022, QN => n13844);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => n6780, CK => CLK, Q => 
                           n_2023, QN => n13845);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => n6779, CK => CLK, Q => 
                           n_2024, QN => n13846);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => n6778, CK => CLK, Q => 
                           n_2025, QN => n13847);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n6909, CK => CLK, Q => n9885
                           , QN => n13849);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n6908, CK => CLK, Q => n9886
                           , QN => n13850);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n6907, CK => CLK, Q => n9887
                           , QN => n13851);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n6906, CK => CLK, Q => n9888
                           , QN => n13852);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n6973, CK => CLK, Q => 
                           n_2026, QN => n14409);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n6972, CK => CLK, Q => 
                           n_2027, QN => n14410);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n6971, CK => CLK, Q => 
                           n_2028, QN => n14411);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => n5373, CK => CLK, Q => 
                           n13816, QN => n4848);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => n5372, CK => CLK, Q => 
                           n13817, QN => n7109);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => n5371, CK => CLK, Q => 
                           n13818, QN => n7126);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => n5370, CK => CLK, Q => 
                           n13819, QN => n7143);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => n5309, CK => CLK, Q => 
                           n13820, QN => n4847);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => n5308, CK => CLK, Q => 
                           n13821, QN => n7108);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => n5307, CK => CLK, Q => 
                           n13822, QN => n7125);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => n5306, CK => CLK, Q => 
                           n13823, QN => n7142);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => n5117, CK => CLK, Q => 
                           n13824, QN => n4850);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => n5116, CK => CLK, Q => 
                           n13825, QN => n7111);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => n5115, CK => CLK, Q => 
                           n13826, QN => n7128);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => n5114, CK => CLK, Q => 
                           n13827, QN => n7145);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => n5053, CK => CLK, Q => 
                           n14156, QN => n4849);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => n5052, CK => CLK, Q => 
                           n14157, QN => n7110);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => n5051, CK => CLK, Q => 
                           n14158, QN => n7127);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => n5050, CK => CLK, Q => 
                           n14159, QN => n7144);
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => n5693, CK => CLK, Q => 
                           n_2029, QN => n4845);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => n5692, CK => CLK, Q => 
                           n_2030, QN => n7106);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => n5691, CK => CLK, Q => 
                           n_2031, QN => n7123);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => n5690, CK => CLK, Q => 
                           n_2032, QN => n7140);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => n5757, CK => CLK, Q => 
                           n_2033, QN => n4846);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => n5756, CK => CLK, Q => 
                           n_2034, QN => n7107);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => n5755, CK => CLK, Q => 
                           n_2035, QN => n7124);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => n5754, CK => CLK, Q => 
                           n_2036, QN => n7141);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => n5949, CK => CLK, Q => 
                           n_2037, QN => n4843);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => n5948, CK => CLK, Q => 
                           n_2038, QN => n4860);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => n5947, CK => CLK, Q => 
                           n_2039, QN => n7121);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => n5946, CK => CLK, Q => 
                           n_2040, QN => n7138);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => n6013, CK => CLK, Q => 
                           n_2041, QN => n4844);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => n6012, CK => CLK, Q => 
                           n_2042, QN => n4861);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => n6011, CK => CLK, Q => 
                           n_2043, QN => n7122);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => n6010, CK => CLK, Q => 
                           n_2044, QN => n7139);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => n6461, CK => CLK, Q => 
                           n13853, QN => n4839);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => n6460, CK => CLK, Q => 
                           n13854, QN => n4856);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => n6459, CK => CLK, Q => 
                           n13855, QN => n7117);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => n6458, CK => CLK, Q => 
                           n13856, QN => n7134);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => n6525, CK => CLK, Q => 
                           n13857, QN => n4840);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => n6524, CK => CLK, Q => 
                           n13858, QN => n4857);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => n6523, CK => CLK, Q => 
                           n13859, QN => n7118);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => n6522, CK => CLK, Q => 
                           n13860, QN => n7135);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => n6205, CK => CLK, Q => 
                           n13865, QN => n4841);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => n6204, CK => CLK, Q => 
                           n13866, QN => n4858);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => n6203, CK => CLK, Q => 
                           n13867, QN => n7119);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => n6202, CK => CLK, Q => 
                           n13868, QN => n7136);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => n6269, CK => CLK, Q => 
                           n13861, QN => n4842);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => n6268, CK => CLK, Q => 
                           n13862, QN => n4859);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => n6267, CK => CLK, Q => 
                           n13863, QN => n7120);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => n6266, CK => CLK, Q => 
                           n13864, QN => n7137);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => n6589, CK => CLK, Q => 
                           n13832, QN => n4838);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => n6588, CK => CLK, Q => 
                           n13833, QN => n4855);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => n6587, CK => CLK, Q => 
                           n13834, QN => n7116);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => n6586, CK => CLK, Q => 
                           n13835, QN => n7133);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => n6653, CK => CLK, Q => 
                           n13836, QN => n4837);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => n6652, CK => CLK, Q => 
                           n13837, QN => n4854);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => n6651, CK => CLK, Q => 
                           n13838, QN => n7115);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => n6650, CK => CLK, Q => 
                           n13839, QN => n7132);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => n5369, CK => CLK, Q => 
                           n13893, QN => n7240);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => n5368, CK => CLK, Q => 
                           n13894, QN => n7257);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => n5367, CK => CLK, Q => 
                           n13895, QN => n7274);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => n5366, CK => CLK, Q => 
                           n13896, QN => n7373);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => n5365, CK => CLK, Q => 
                           n13897, QN => n7390);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => n5364, CK => CLK, Q => 
                           n13898, QN => n7492);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => n5363, CK => CLK, Q => 
                           n13899, QN => n7509);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => n5362, CK => CLK, Q => 
                           n13900, QN => n7526);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => n5361, CK => CLK, Q => 
                           n13901, QN => n7630);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => n5360, CK => CLK, Q => 
                           n13902, QN => n7647);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => n5359, CK => CLK, Q => 
                           n13903, QN => n7749);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => n5358, CK => CLK, Q => 
                           n13904, QN => n7766);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => n5357, CK => CLK, Q => 
                           n13905, QN => n7783);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => n5356, CK => CLK, Q => 
                           n13906, QN => n7800);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => n5355, CK => CLK, Q => 
                           n13907, QN => n7817);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => n5354, CK => CLK, Q => 
                           n13908, QN => n7834);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => n5353, CK => CLK, Q => 
                           n13909, QN => n7851);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => n5352, CK => CLK, Q => 
                           n13910, QN => n7868);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => n5351, CK => CLK, Q => 
                           n13911, QN => n7885);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => n5350, CK => CLK, Q => 
                           n13912, QN => n7902);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => n5349, CK => CLK, Q => 
                           n13913, QN => n7919);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => n5348, CK => CLK, Q => 
                           n13914, QN => n7936);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => n5347, CK => CLK, Q => 
                           n13915, QN => n7953);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => n5346, CK => CLK, Q => 
                           n13916, QN => n7970);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => n5345, CK => CLK, Q => 
                           n13917, QN => n7987);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => n5344, CK => CLK, Q => 
                           n13918, QN => n8004);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => n5343, CK => CLK, Q => 
                           n13919, QN => n8021);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => n5342, CK => CLK, Q => 
                           n13920, QN => n8038);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n5341, CK => CLK, Q => 
                           n13921, QN => n8055);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n5340, CK => CLK, Q => 
                           n13922, QN => n8072);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n5339, CK => CLK, Q => 
                           n13923, QN => n8089);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n5338, CK => CLK, Q => 
                           n13924, QN => n8106);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n5337, CK => CLK, Q => 
                           n13925, QN => n8123);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n5336, CK => CLK, Q => 
                           n13926, QN => n8140);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n5335, CK => CLK, Q => 
                           n13927, QN => n8157);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n5334, CK => CLK, Q => 
                           n13928, QN => n8174);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => n5305, CK => CLK, Q => 
                           n13953, QN => n7239);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => n5304, CK => CLK, Q => 
                           n13954, QN => n7256);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => n5303, CK => CLK, Q => 
                           n13955, QN => n7273);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => n5302, CK => CLK, Q => 
                           n13956, QN => n7372);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => n5301, CK => CLK, Q => 
                           n13957, QN => n7389);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => n5300, CK => CLK, Q => 
                           n13958, QN => n7491);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => n5299, CK => CLK, Q => 
                           n13959, QN => n7508);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => n5298, CK => CLK, Q => 
                           n13960, QN => n7525);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => n5297, CK => CLK, Q => 
                           n13961, QN => n7629);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => n5296, CK => CLK, Q => 
                           n13962, QN => n7646);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => n5295, CK => CLK, Q => 
                           n13963, QN => n7748);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => n5294, CK => CLK, Q => 
                           n13964, QN => n7765);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => n5293, CK => CLK, Q => 
                           n13965, QN => n7782);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => n5292, CK => CLK, Q => 
                           n13966, QN => n7799);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => n5291, CK => CLK, Q => 
                           n13967, QN => n7816);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => n5290, CK => CLK, Q => 
                           n13968, QN => n7833);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => n5289, CK => CLK, Q => 
                           n13969, QN => n7850);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => n5288, CK => CLK, Q => 
                           n13970, QN => n7867);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => n5287, CK => CLK, Q => 
                           n13971, QN => n7884);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => n5286, CK => CLK, Q => 
                           n13972, QN => n7901);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => n5285, CK => CLK, Q => 
                           n13973, QN => n7918);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => n5284, CK => CLK, Q => 
                           n13974, QN => n7935);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => n5283, CK => CLK, Q => 
                           n13975, QN => n7952);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => n5282, CK => CLK, Q => 
                           n13976, QN => n7969);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => n5281, CK => CLK, Q => 
                           n13977, QN => n7986);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => n5280, CK => CLK, Q => 
                           n13978, QN => n8003);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => n5279, CK => CLK, Q => 
                           n13979, QN => n8020);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => n5278, CK => CLK, Q => 
                           n13980, QN => n8037);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n5277, CK => CLK, Q => 
                           n13981, QN => n8054);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n5276, CK => CLK, Q => 
                           n13982, QN => n8071);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n5275, CK => CLK, Q => 
                           n13983, QN => n8088);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n5274, CK => CLK, Q => 
                           n13984, QN => n8105);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n5273, CK => CLK, Q => 
                           n13985, QN => n8122);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n5272, CK => CLK, Q => 
                           n13986, QN => n8139);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n5271, CK => CLK, Q => 
                           n13987, QN => n8156);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n5270, CK => CLK, Q => 
                           n13988, QN => n8173);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => n5113, CK => CLK, Q => 
                           n13989, QN => n7242);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => n5112, CK => CLK, Q => 
                           n13990, QN => n7259);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => n5111, CK => CLK, Q => 
                           n13991, QN => n7276);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => n5110, CK => CLK, Q => 
                           n13992, QN => n7375);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => n5109, CK => CLK, Q => 
                           n13993, QN => n7392);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => n5108, CK => CLK, Q => 
                           n13994, QN => n7494);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => n5107, CK => CLK, Q => 
                           n13995, QN => n7511);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => n5106, CK => CLK, Q => 
                           n13996, QN => n7528);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => n5105, CK => CLK, Q => 
                           n13997, QN => n7632);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => n5104, CK => CLK, Q => 
                           n13998, QN => n7649);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => n5103, CK => CLK, Q => 
                           n13999, QN => n7751);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => n5102, CK => CLK, Q => 
                           n14000, QN => n7768);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => n5101, CK => CLK, Q => 
                           n14001, QN => n7785);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => n5100, CK => CLK, Q => 
                           n14002, QN => n7802);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => n5099, CK => CLK, Q => 
                           n14003, QN => n7819);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => n5098, CK => CLK, Q => 
                           n14004, QN => n7836);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => n5097, CK => CLK, Q => 
                           n14005, QN => n7853);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => n5096, CK => CLK, Q => 
                           n14006, QN => n7870);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => n5095, CK => CLK, Q => 
                           n14007, QN => n7887);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => n5094, CK => CLK, Q => 
                           n14008, QN => n7904);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => n5093, CK => CLK, Q => 
                           n14009, QN => n7921);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => n5092, CK => CLK, Q => 
                           n14010, QN => n7938);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => n5091, CK => CLK, Q => 
                           n14011, QN => n7955);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => n5090, CK => CLK, Q => 
                           n14012, QN => n7972);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => n5089, CK => CLK, Q => 
                           n14013, QN => n7989);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => n5088, CK => CLK, Q => 
                           n14014, QN => n8006);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => n5087, CK => CLK, Q => 
                           n14015, QN => n8023);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => n5086, CK => CLK, Q => 
                           n14016, QN => n8040);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n5085, CK => CLK, Q => 
                           n14017, QN => n8057);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n5084, CK => CLK, Q => 
                           n14018, QN => n8074);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n5083, CK => CLK, Q => 
                           n14019, QN => n8091);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n5082, CK => CLK, Q => 
                           n14020, QN => n8108);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n5081, CK => CLK, Q => 
                           n14021, QN => n8125);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n5080, CK => CLK, Q => 
                           n14022, QN => n8142);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n5079, CK => CLK, Q => 
                           n14023, QN => n8159);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n5078, CK => CLK, Q => 
                           n14024, QN => n8176);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n5333, CK => CLK, Q => 
                           n14060, QN => n8191);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n5332, CK => CLK, Q => 
                           n14061, QN => n8208);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n5331, CK => CLK, Q => 
                           n14062, QN => n8225);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n5330, CK => CLK, Q => 
                           n14063, QN => n8242);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n5329, CK => CLK, Q => 
                           n14064, QN => n8259);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n5328, CK => CLK, Q => 
                           n14065, QN => n8276);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n5327, CK => CLK, Q => 
                           n14066, QN => n8293);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n5326, CK => CLK, Q => 
                           n14067, QN => n8310);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n5325, CK => CLK, Q => 
                           n14068, QN => n8327);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n5324, CK => CLK, Q => 
                           n14069, QN => n8344);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n5323, CK => CLK, Q => 
                           n14070, QN => n8361);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n5322, CK => CLK, Q => 
                           n14071, QN => n8378);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n5321, CK => CLK, Q => 
                           n14072, QN => n8395);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n5320, CK => CLK, Q => 
                           n14073, QN => n8412);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n5319, CK => CLK, Q => 
                           n14074, QN => n8429);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n5318, CK => CLK, Q => 
                           n14075, QN => n8446);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n5317, CK => CLK, Q => 
                           n14076, QN => n8463);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n5316, CK => CLK, Q => 
                           n14077, QN => n8480);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n5315, CK => CLK, Q => 
                           n14078, QN => n8497);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n5313, CK => CLK, Q => 
                           n14079, QN => n8531);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n5314, CK => CLK, Q => 
                           n14080, QN => n8514);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n5312, CK => CLK, Q => 
                           n14081, QN => n8548);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n5311, CK => CLK, Q => 
                           n14082, QN => n8565);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n5310, CK => CLK, Q => 
                           n14153, QN => n8582);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n5269, CK => CLK, Q => 
                           n14107, QN => n8190);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n5268, CK => CLK, Q => 
                           n14108, QN => n8207);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n5267, CK => CLK, Q => 
                           n14109, QN => n8224);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n5266, CK => CLK, Q => 
                           n14110, QN => n8241);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n5265, CK => CLK, Q => 
                           n14111, QN => n8258);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n5264, CK => CLK, Q => 
                           n14112, QN => n8275);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n5263, CK => CLK, Q => 
                           n14113, QN => n8292);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n5262, CK => CLK, Q => 
                           n14114, QN => n8309);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n5261, CK => CLK, Q => 
                           n14115, QN => n8326);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n5260, CK => CLK, Q => 
                           n14116, QN => n8343);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n5259, CK => CLK, Q => 
                           n14117, QN => n8360);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n5258, CK => CLK, Q => 
                           n14118, QN => n8377);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n5257, CK => CLK, Q => 
                           n14119, QN => n8394);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n5256, CK => CLK, Q => 
                           n14120, QN => n8411);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n5255, CK => CLK, Q => 
                           n14121, QN => n8428);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n5254, CK => CLK, Q => 
                           n14122, QN => n8445);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n5253, CK => CLK, Q => 
                           n14123, QN => n8462);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n5252, CK => CLK, Q => 
                           n14124, QN => n8479);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n5251, CK => CLK, Q => 
                           n14125, QN => n8496);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n5249, CK => CLK, Q => 
                           n14126, QN => n8530);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n5250, CK => CLK, Q => 
                           n14127, QN => n8513);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n5248, CK => CLK, Q => 
                           n14128, QN => n8547);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n5247, CK => CLK, Q => 
                           n14129, QN => n8564);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n5246, CK => CLK, Q => 
                           n14154, QN => n8581);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n5077, CK => CLK, Q => 
                           n14130, QN => n8193);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n5076, CK => CLK, Q => 
                           n14131, QN => n8210);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n5075, CK => CLK, Q => 
                           n14132, QN => n8227);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n5074, CK => CLK, Q => 
                           n14133, QN => n8244);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n5073, CK => CLK, Q => 
                           n14134, QN => n8261);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n5072, CK => CLK, Q => 
                           n14135, QN => n8278);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n5071, CK => CLK, Q => 
                           n14136, QN => n8295);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n5070, CK => CLK, Q => 
                           n14137, QN => n8312);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n5069, CK => CLK, Q => 
                           n14138, QN => n8329);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n5068, CK => CLK, Q => 
                           n14139, QN => n8346);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n5067, CK => CLK, Q => 
                           n14140, QN => n8363);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n5066, CK => CLK, Q => 
                           n14141, QN => n8380);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n5065, CK => CLK, Q => 
                           n14142, QN => n8397);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n5064, CK => CLK, Q => 
                           n14143, QN => n8414);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n5063, CK => CLK, Q => 
                           n14144, QN => n8431);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n5062, CK => CLK, Q => 
                           n14145, QN => n8448);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n5061, CK => CLK, Q => 
                           n14146, QN => n8465);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n5060, CK => CLK, Q => 
                           n14147, QN => n8482);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n5059, CK => CLK, Q => 
                           n14148, QN => n8499);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n5057, CK => CLK, Q => 
                           n14149, QN => n8533);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n5058, CK => CLK, Q => 
                           n14150, QN => n8516);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n5056, CK => CLK, Q => 
                           n14151, QN => n8550);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n5055, CK => CLK, Q => 
                           n14152, QN => n8567);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n5054, CK => CLK, Q => 
                           n14155, QN => n8584);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => n5049, CK => CLK, Q => 
                           n14160, QN => n7241);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => n5048, CK => CLK, Q => 
                           n14161, QN => n7258);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => n5047, CK => CLK, Q => 
                           n14162, QN => n7275);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => n5046, CK => CLK, Q => 
                           n14163, QN => n7374);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => n5045, CK => CLK, Q => 
                           n14164, QN => n7391);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => n5044, CK => CLK, Q => 
                           n14165, QN => n7493);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => n5043, CK => CLK, Q => 
                           n14166, QN => n7510);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => n5042, CK => CLK, Q => 
                           n14167, QN => n7527);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => n5041, CK => CLK, Q => 
                           n14168, QN => n7631);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => n5040, CK => CLK, Q => 
                           n14169, QN => n7648);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => n5039, CK => CLK, Q => 
                           n14170, QN => n7750);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => n5038, CK => CLK, Q => 
                           n14171, QN => n7767);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => n5037, CK => CLK, Q => 
                           n14172, QN => n7784);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => n5036, CK => CLK, Q => 
                           n14173, QN => n7801);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => n5035, CK => CLK, Q => 
                           n14174, QN => n7818);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => n5034, CK => CLK, Q => 
                           n14175, QN => n7835);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => n5033, CK => CLK, Q => 
                           n14176, QN => n7852);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => n5032, CK => CLK, Q => 
                           n14177, QN => n7869);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => n5031, CK => CLK, Q => 
                           n14178, QN => n7886);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => n5030, CK => CLK, Q => 
                           n14179, QN => n7903);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => n5029, CK => CLK, Q => 
                           n14180, QN => n7920);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => n5028, CK => CLK, Q => 
                           n14181, QN => n7937);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => n5027, CK => CLK, Q => 
                           n14182, QN => n7954);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => n5026, CK => CLK, Q => 
                           n14183, QN => n7971);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => n5025, CK => CLK, Q => 
                           n14184, QN => n7988);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => n5024, CK => CLK, Q => 
                           n14185, QN => n8005);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => n5023, CK => CLK, Q => 
                           n14186, QN => n8022);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => n5022, CK => CLK, Q => 
                           n14187, QN => n8039);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n5021, CK => CLK, Q => 
                           n14188, QN => n8056);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n5020, CK => CLK, Q => 
                           n14189, QN => n8073);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n5019, CK => CLK, Q => 
                           n14190, QN => n8090);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n5018, CK => CLK, Q => 
                           n14191, QN => n8107);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n5017, CK => CLK, Q => 
                           n14192, QN => n8124);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n5016, CK => CLK, Q => 
                           n14193, QN => n8141);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n5015, CK => CLK, Q => 
                           n14194, QN => n8158);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n5014, CK => CLK, Q => 
                           n14195, QN => n8175);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n5013, CK => CLK, Q => 
                           n14196, QN => n8192);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n5012, CK => CLK, Q => 
                           n14197, QN => n8209);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n5011, CK => CLK, Q => 
                           n14198, QN => n8226);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n5010, CK => CLK, Q => 
                           n14199, QN => n8243);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n5009, CK => CLK, Q => 
                           n14200, QN => n8260);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n5008, CK => CLK, Q => 
                           n14201, QN => n8277);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n5007, CK => CLK, Q => 
                           n14202, QN => n8294);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n5006, CK => CLK, Q => 
                           n14203, QN => n8311);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n5005, CK => CLK, Q => 
                           n14204, QN => n8328);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n5004, CK => CLK, Q => 
                           n14205, QN => n8345);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n5003, CK => CLK, Q => 
                           n14206, QN => n8362);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n5002, CK => CLK, Q => 
                           n14207, QN => n8379);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n5001, CK => CLK, Q => 
                           n14208, QN => n8396);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n5000, CK => CLK, Q => 
                           n14209, QN => n8413);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n4999, CK => CLK, Q => 
                           n14210, QN => n8430);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n4998, CK => CLK, Q => 
                           n14211, QN => n8447);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n4997, CK => CLK, Q => 
                           n14212, QN => n8464);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n4996, CK => CLK, Q => 
                           n14213, QN => n8481);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n4995, CK => CLK, Q => 
                           n14214, QN => n8498);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n4994, CK => CLK, Q => 
                           n14215, QN => n8515);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n4993, CK => CLK, Q => 
                           n13828, QN => n8532);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n4992, CK => CLK, Q => 
                           n13829, QN => n8549);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n4991, CK => CLK, Q => 
                           n13830, QN => n8566);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n4990, CK => CLK, Q => 
                           n13831, QN => n8583);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => n5689, CK => CLK, Q => 
                           n_2045, QN => n7237);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => n5688, CK => CLK, Q => 
                           n_2046, QN => n7254);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => n5687, CK => CLK, Q => 
                           n_2047, QN => n7271);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => n5686, CK => CLK, Q => 
                           n_2048, QN => n7370);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => n5685, CK => CLK, Q => 
                           n_2049, QN => n7387);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => n5684, CK => CLK, Q => 
                           n_2050, QN => n7404);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => n5683, CK => CLK, Q => 
                           n_2051, QN => n7506);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => n5682, CK => CLK, Q => 
                           n_2052, QN => n7523);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => n5681, CK => CLK, Q => 
                           n_2053, QN => n7627);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => n5680, CK => CLK, Q => 
                           n_2054, QN => n7644);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => n5679, CK => CLK, Q => 
                           n_2055, QN => n7746);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => n5678, CK => CLK, Q => 
                           n_2056, QN => n7763);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => n5677, CK => CLK, Q => 
                           n_2057, QN => n7780);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => n5676, CK => CLK, Q => 
                           n_2058, QN => n7797);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => n5675, CK => CLK, Q => 
                           n_2059, QN => n7814);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => n5674, CK => CLK, Q => 
                           n_2060, QN => n7831);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => n5673, CK => CLK, Q => 
                           n_2061, QN => n7848);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => n5672, CK => CLK, Q => 
                           n_2062, QN => n7865);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => n5671, CK => CLK, Q => 
                           n_2063, QN => n7882);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => n5670, CK => CLK, Q => 
                           n_2064, QN => n7899);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => n5669, CK => CLK, Q => 
                           n_2065, QN => n7916);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => n5668, CK => CLK, Q => 
                           n_2066, QN => n7933);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => n5667, CK => CLK, Q => 
                           n_2067, QN => n7950);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => n5666, CK => CLK, Q => 
                           n_2068, QN => n7967);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => n5665, CK => CLK, Q => 
                           n_2069, QN => n7984);
   U3 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n4450);
   U4 : NOR2_X1 port map( A1 => n13389, A2 => ADD_RD2(1), ZN => n4454);
   U5 : AND3_X1 port map( A1 => ENABLE, A2 => n12139, A3 => RD2, ZN => n3211);
   U6 : NAND2_X1 port map( A1 => n3209, A2 => n3189, ZN => n1995);
   U7 : CLKBUF_X1 port map( A => n12614, Z => n12612);
   U8 : CLKBUF_X1 port map( A => n12690, Z => n12688);
   U9 : CLKBUF_X1 port map( A => n12633, Z => n12631);
   U10 : CLKBUF_X1 port map( A => n12709, Z => n12707);
   U11 : CLKBUF_X1 port map( A => n12595, Z => n12593);
   U12 : CLKBUF_X1 port map( A => n12652, Z => n12650);
   U13 : CLKBUF_X1 port map( A => n12671, Z => n12669);
   U14 : BUF_X1 port map( A => n1910, Z => n13130);
   U15 : BUF_X1 port map( A => n1912, Z => n13110);
   U16 : BUF_X1 port map( A => n1914, Z => n13090);
   U17 : BUF_X1 port map( A => n1916, Z => n13070);
   U18 : BUF_X1 port map( A => n1918, Z => n13050);
   U19 : BUF_X1 port map( A => n1920, Z => n13030);
   U20 : BUF_X1 port map( A => n1908, Z => n13150);
   U21 : BUF_X1 port map( A => n1842, Z => n13359);
   U22 : BUF_X1 port map( A => n1932, Z => n12850);
   U23 : BUF_X1 port map( A => n1934, Z => n12830);
   U24 : BUF_X1 port map( A => n1937, Z => n12770);
   U25 : BUF_X1 port map( A => n1938, Z => n12750);
   U26 : BUF_X1 port map( A => n1940, Z => n12710);
   U27 : BUF_X1 port map( A => n1939, Z => n12730);
   U28 : BUF_X1 port map( A => n1936, Z => n12790);
   U29 : BUF_X1 port map( A => n1935, Z => n12810);
   U30 : BUF_X1 port map( A => n1928, Z => n12930);
   U31 : BUF_X1 port map( A => n1923, Z => n13010);
   U32 : BUF_X1 port map( A => n1925, Z => n12990);
   U33 : BUF_X1 port map( A => n1929, Z => n12910);
   U34 : BUF_X1 port map( A => n1948, Z => n12577);
   U35 : BUF_X1 port map( A => n1945, Z => n12634);
   U36 : BUF_X1 port map( A => n1947, Z => n12596);
   U37 : BUF_X1 port map( A => n1931, Z => n12870);
   U38 : BUF_X1 port map( A => n1930, Z => n12890);
   U39 : BUF_X1 port map( A => n1927, Z => n12950);
   U40 : BUF_X1 port map( A => n1944, Z => n12653);
   U41 : BUF_X1 port map( A => n1946, Z => n12615);
   U42 : BUF_X1 port map( A => n1943, Z => n12672);
   U43 : BUF_X1 port map( A => n1941, Z => n12691);
   U44 : BUF_X1 port map( A => n1926, Z => n12970);
   U45 : INV_X1 port map( A => n12573, ZN => n12552);
   U46 : INV_X1 port map( A => n12573, ZN => n12553);
   U47 : INV_X1 port map( A => n12573, ZN => n12554);
   U48 : INV_X1 port map( A => n12573, ZN => n12555);
   U49 : INV_X1 port map( A => n12573, ZN => n12551);
   U50 : INV_X1 port map( A => n13128, ZN => n13112);
   U51 : INV_X1 port map( A => n13128, ZN => n13113);
   U52 : INV_X1 port map( A => n13128, ZN => n13114);
   U53 : INV_X1 port map( A => n13007, ZN => n12991);
   U54 : INV_X1 port map( A => n12847, ZN => n12831);
   U55 : INV_X1 port map( A => n12787, ZN => n12771);
   U56 : INV_X1 port map( A => n12767, ZN => n12751);
   U57 : INV_X1 port map( A => n12927, ZN => n12911);
   U58 : INV_X1 port map( A => n13027, ZN => n13011);
   U59 : INV_X1 port map( A => n13067, ZN => n13051);
   U60 : INV_X1 port map( A => n13047, ZN => n13031);
   U61 : INV_X1 port map( A => n12928, ZN => n12912);
   U62 : INV_X1 port map( A => n12928, ZN => n12913);
   U63 : INV_X1 port map( A => n12928, ZN => n12914);
   U64 : INV_X1 port map( A => n12948, ZN => n12932);
   U65 : INV_X1 port map( A => n12948, ZN => n12933);
   U66 : INV_X1 port map( A => n12948, ZN => n12934);
   U67 : INV_X1 port map( A => n13028, ZN => n13012);
   U68 : INV_X1 port map( A => n13028, ZN => n13013);
   U69 : INV_X1 port map( A => n13028, ZN => n13014);
   U70 : INV_X1 port map( A => n13008, ZN => n12992);
   U71 : INV_X1 port map( A => n13008, ZN => n12993);
   U72 : INV_X1 port map( A => n13008, ZN => n12994);
   U73 : INV_X1 port map( A => n13068, ZN => n13052);
   U74 : INV_X1 port map( A => n13068, ZN => n13053);
   U75 : INV_X1 port map( A => n13068, ZN => n13054);
   U76 : INV_X1 port map( A => n13048, ZN => n13032);
   U77 : INV_X1 port map( A => n13048, ZN => n13033);
   U78 : INV_X1 port map( A => n13048, ZN => n13034);
   U79 : INV_X1 port map( A => n12867, ZN => n12851);
   U80 : INV_X1 port map( A => n12868, ZN => n12852);
   U81 : INV_X1 port map( A => n12868, ZN => n12853);
   U82 : INV_X1 port map( A => n12868, ZN => n12854);
   U83 : INV_X1 port map( A => n12848, ZN => n12832);
   U84 : INV_X1 port map( A => n12848, ZN => n12833);
   U85 : INV_X1 port map( A => n12848, ZN => n12834);
   U86 : INV_X1 port map( A => n12788, ZN => n12772);
   U87 : INV_X1 port map( A => n12788, ZN => n12773);
   U88 : INV_X1 port map( A => n12788, ZN => n12774);
   U89 : INV_X1 port map( A => n12768, ZN => n12752);
   U90 : INV_X1 port map( A => n12768, ZN => n12753);
   U91 : INV_X1 port map( A => n12768, ZN => n12754);
   U92 : INV_X1 port map( A => n12594, ZN => n12578);
   U93 : INV_X1 port map( A => n12594, ZN => n12579);
   U94 : INV_X1 port map( A => n12594, ZN => n12580);
   U95 : INV_X1 port map( A => n12651, ZN => n12635);
   U96 : INV_X1 port map( A => n12651, ZN => n12636);
   U97 : INV_X1 port map( A => n12651, ZN => n12637);
   U98 : INV_X1 port map( A => n12670, ZN => n12654);
   U99 : INV_X1 port map( A => n12670, ZN => n12655);
   U100 : INV_X1 port map( A => n12670, ZN => n12656);
   U101 : INV_X1 port map( A => n13127, ZN => n13111);
   U102 : INV_X1 port map( A => n13147, ZN => n13131);
   U103 : INV_X1 port map( A => n13107, ZN => n13091);
   U104 : INV_X1 port map( A => n13087, ZN => n13071);
   U105 : INV_X1 port map( A => n13376, ZN => n13360);
   U106 : INV_X1 port map( A => n12807, ZN => n12791);
   U107 : INV_X1 port map( A => n12727, ZN => n12711);
   U108 : INV_X1 port map( A => n12747, ZN => n12731);
   U109 : INV_X1 port map( A => n12827, ZN => n12811);
   U110 : INV_X1 port map( A => n12887, ZN => n12871);
   U111 : INV_X1 port map( A => n12907, ZN => n12891);
   U112 : INV_X1 port map( A => n12967, ZN => n12951);
   U113 : INV_X1 port map( A => n12987, ZN => n12971);
   U114 : INV_X1 port map( A => n13167, ZN => n13151);
   U115 : INV_X1 port map( A => n13168, ZN => n13154);
   U116 : INV_X1 port map( A => n13168, ZN => n13153);
   U117 : INV_X1 port map( A => n13377, ZN => n13361);
   U118 : INV_X1 port map( A => n13148, ZN => n13132);
   U119 : INV_X1 port map( A => n13148, ZN => n13133);
   U120 : INV_X1 port map( A => n13148, ZN => n13134);
   U121 : INV_X1 port map( A => n13108, ZN => n13092);
   U122 : INV_X1 port map( A => n13108, ZN => n13093);
   U123 : INV_X1 port map( A => n13108, ZN => n13094);
   U124 : INV_X1 port map( A => n13088, ZN => n13072);
   U125 : INV_X1 port map( A => n13088, ZN => n13073);
   U126 : INV_X1 port map( A => n13088, ZN => n13074);
   U127 : INV_X1 port map( A => n12808, ZN => n12792);
   U128 : INV_X1 port map( A => n12728, ZN => n12713);
   U129 : INV_X1 port map( A => n12728, ZN => n12712);
   U130 : INV_X1 port map( A => n12613, ZN => n12599);
   U131 : INV_X1 port map( A => n12689, ZN => n12674);
   U132 : INV_X1 port map( A => n12613, ZN => n12597);
   U133 : INV_X1 port map( A => n12613, ZN => n12598);
   U134 : INV_X1 port map( A => n12689, ZN => n12673);
   U135 : INV_X1 port map( A => n12632, ZN => n12616);
   U136 : INV_X1 port map( A => n12632, ZN => n12617);
   U137 : INV_X1 port map( A => n12632, ZN => n12618);
   U138 : INV_X1 port map( A => n12689, ZN => n12675);
   U139 : INV_X1 port map( A => n12708, ZN => n12692);
   U140 : INV_X1 port map( A => n12708, ZN => n12693);
   U141 : INV_X1 port map( A => n12708, ZN => n12694);
   U142 : INV_X1 port map( A => n12728, ZN => n12714);
   U143 : INV_X1 port map( A => n12748, ZN => n12732);
   U144 : INV_X1 port map( A => n12748, ZN => n12733);
   U145 : INV_X1 port map( A => n12748, ZN => n12734);
   U146 : INV_X1 port map( A => n12808, ZN => n12793);
   U147 : INV_X1 port map( A => n12808, ZN => n12794);
   U148 : INV_X1 port map( A => n12828, ZN => n12812);
   U149 : INV_X1 port map( A => n12828, ZN => n12813);
   U150 : INV_X1 port map( A => n12828, ZN => n12814);
   U151 : INV_X1 port map( A => n12888, ZN => n12872);
   U152 : INV_X1 port map( A => n12888, ZN => n12873);
   U153 : INV_X1 port map( A => n12888, ZN => n12874);
   U154 : INV_X1 port map( A => n12908, ZN => n12892);
   U155 : INV_X1 port map( A => n12908, ZN => n12893);
   U156 : INV_X1 port map( A => n12908, ZN => n12894);
   U157 : INV_X1 port map( A => n12968, ZN => n12952);
   U158 : INV_X1 port map( A => n12968, ZN => n12953);
   U159 : INV_X1 port map( A => n12968, ZN => n12954);
   U160 : INV_X1 port map( A => n12988, ZN => n12972);
   U161 : INV_X1 port map( A => n12988, ZN => n12973);
   U162 : INV_X1 port map( A => n12988, ZN => n12974);
   U163 : INV_X1 port map( A => n13168, ZN => n13152);
   U164 : INV_X1 port map( A => n13377, ZN => n13362);
   U165 : INV_X1 port map( A => n13377, ZN => n13363);
   U166 : INV_X1 port map( A => n12947, ZN => n12931);
   U167 : BUF_X1 port map( A => n12575, Z => n12573);
   U168 : BUF_X1 port map( A => n12576, Z => n12571);
   U169 : BUF_X1 port map( A => n12574, Z => n12570);
   U170 : BUF_X1 port map( A => n12575, Z => n12569);
   U171 : BUF_X1 port map( A => n12574, Z => n12568);
   U172 : BUF_X1 port map( A => n12574, Z => n12567);
   U173 : BUF_X1 port map( A => n12574, Z => n12566);
   U174 : BUF_X1 port map( A => n12574, Z => n12565);
   U175 : BUF_X1 port map( A => n12575, Z => n12564);
   U176 : BUF_X1 port map( A => n12575, Z => n12563);
   U177 : BUF_X1 port map( A => n12575, Z => n12562);
   U178 : BUF_X1 port map( A => n12576, Z => n12561);
   U179 : BUF_X1 port map( A => n12576, Z => n12560);
   U180 : BUF_X1 port map( A => n12576, Z => n12559);
   U181 : BUF_X1 port map( A => n12574, Z => n12572);
   U182 : BUF_X1 port map( A => n12576, Z => n12558);
   U183 : BUF_X1 port map( A => n12576, Z => n12557);
   U184 : BUF_X1 port map( A => n1998, Z => n12357);
   U185 : BUF_X1 port map( A => n1998, Z => n12358);
   U186 : BUF_X1 port map( A => n1998, Z => n12359);
   U187 : BUF_X1 port map( A => n1998, Z => n12360);
   U188 : BUF_X1 port map( A => n1998, Z => n12361);
   U189 : BUF_X1 port map( A => n12929, Z => n12927);
   U190 : BUF_X1 port map( A => n12949, Z => n12947);
   U191 : BUF_X1 port map( A => n13009, Z => n13007);
   U192 : BUF_X1 port map( A => n13149, Z => n13147);
   U193 : BUF_X1 port map( A => n13109, Z => n13107);
   U194 : BUF_X1 port map( A => n13089, Z => n13087);
   U195 : BUF_X1 port map( A => n13378, Z => n13376);
   U196 : BUF_X1 port map( A => n12849, Z => n12847);
   U197 : BUF_X1 port map( A => n12789, Z => n12787);
   U198 : BUF_X1 port map( A => n12769, Z => n12767);
   U199 : BUF_X1 port map( A => n12729, Z => n12727);
   U200 : BUF_X1 port map( A => n12749, Z => n12747);
   U201 : BUF_X1 port map( A => n12809, Z => n12807);
   U202 : BUF_X1 port map( A => n12829, Z => n12827);
   U203 : BUF_X1 port map( A => n12889, Z => n12887);
   U204 : BUF_X1 port map( A => n12909, Z => n12907);
   U205 : BUF_X1 port map( A => n12969, Z => n12967);
   U206 : BUF_X1 port map( A => n12989, Z => n12987);
   U207 : BUF_X1 port map( A => n13169, Z => n13167);
   U208 : BUF_X1 port map( A => n13021, Z => n13024);
   U209 : BUF_X1 port map( A => n13020, Z => n13023);
   U210 : BUF_X1 port map( A => n13041, Z => n13044);
   U211 : BUF_X1 port map( A => n13040, Z => n13043);
   U212 : BUF_X1 port map( A => n13015, Z => n13022);
   U213 : BUF_X1 port map( A => n13029, Z => n13021);
   U214 : BUF_X1 port map( A => n13029, Z => n13020);
   U215 : BUF_X1 port map( A => n13029, Z => n13019);
   U216 : BUF_X1 port map( A => n13029, Z => n13018);
   U217 : BUF_X1 port map( A => n13029, Z => n13017);
   U218 : BUF_X1 port map( A => n13029, Z => n13016);
   U219 : BUF_X1 port map( A => n13035, Z => n13042);
   U220 : BUF_X1 port map( A => n13049, Z => n13041);
   U221 : BUF_X1 port map( A => n13049, Z => n13040);
   U222 : BUF_X1 port map( A => n13049, Z => n13039);
   U223 : BUF_X1 port map( A => n13049, Z => n13038);
   U224 : BUF_X1 port map( A => n13049, Z => n13037);
   U225 : BUF_X1 port map( A => n13049, Z => n13036);
   U226 : BUF_X1 port map( A => n13029, Z => n13015);
   U227 : BUF_X1 port map( A => n13049, Z => n13035);
   U228 : BUF_X1 port map( A => n12929, Z => n12926);
   U229 : BUF_X1 port map( A => n12929, Z => n12925);
   U230 : BUF_X1 port map( A => n12929, Z => n12924);
   U231 : BUF_X1 port map( A => n12929, Z => n12923);
   U232 : BUF_X1 port map( A => n12941, Z => n12944);
   U233 : BUF_X1 port map( A => n13009, Z => n13006);
   U234 : BUF_X1 port map( A => n13009, Z => n13005);
   U235 : BUF_X1 port map( A => n13009, Z => n13004);
   U236 : BUF_X1 port map( A => n13009, Z => n13003);
   U237 : BUF_X1 port map( A => n13371, Z => n13369);
   U238 : BUF_X1 port map( A => n13375, Z => n13368);
   U239 : BUF_X1 port map( A => n13162, Z => n13158);
   U240 : BUF_X1 port map( A => n13166, Z => n13157);
   U241 : BUF_X1 port map( A => n13165, Z => n13156);
   U242 : BUF_X1 port map( A => n13164, Z => n13155);
   U243 : BUF_X1 port map( A => n13149, Z => n13146);
   U244 : BUF_X1 port map( A => n13149, Z => n13145);
   U245 : BUF_X1 port map( A => n13149, Z => n13144);
   U246 : BUF_X1 port map( A => n13149, Z => n13143);
   U247 : BUF_X1 port map( A => n13121, Z => n13124);
   U248 : BUF_X1 port map( A => n13120, Z => n13123);
   U249 : BUF_X1 port map( A => n13109, Z => n13106);
   U250 : BUF_X1 port map( A => n13109, Z => n13105);
   U251 : BUF_X1 port map( A => n13109, Z => n13104);
   U252 : BUF_X1 port map( A => n13109, Z => n13103);
   U253 : BUF_X1 port map( A => n13089, Z => n13086);
   U254 : BUF_X1 port map( A => n13089, Z => n13085);
   U255 : BUF_X1 port map( A => n13089, Z => n13084);
   U256 : BUF_X1 port map( A => n13089, Z => n13083);
   U257 : BUF_X1 port map( A => n13061, Z => n13064);
   U258 : BUF_X1 port map( A => n13060, Z => n13063);
   U259 : BUF_X1 port map( A => n12889, Z => n12886);
   U260 : BUF_X1 port map( A => n12889, Z => n12885);
   U261 : BUF_X1 port map( A => n12969, Z => n12966);
   U262 : BUF_X1 port map( A => n12969, Z => n12965);
   U263 : BUF_X1 port map( A => n12929, Z => n12922);
   U264 : BUF_X1 port map( A => n12922, Z => n12921);
   U265 : BUF_X1 port map( A => n12926, Z => n12920);
   U266 : BUF_X1 port map( A => n12925, Z => n12919);
   U267 : BUF_X1 port map( A => n12924, Z => n12918);
   U268 : BUF_X1 port map( A => n12923, Z => n12917);
   U269 : BUF_X1 port map( A => n12922, Z => n12916);
   U270 : BUF_X1 port map( A => n12940, Z => n12942);
   U271 : BUF_X1 port map( A => n12949, Z => n12941);
   U272 : BUF_X1 port map( A => n12949, Z => n12940);
   U273 : BUF_X1 port map( A => n12949, Z => n12939);
   U274 : BUF_X1 port map( A => n12949, Z => n12938);
   U275 : BUF_X1 port map( A => n12949, Z => n12937);
   U276 : BUF_X1 port map( A => n12949, Z => n12936);
   U277 : BUF_X1 port map( A => n13009, Z => n13002);
   U278 : BUF_X1 port map( A => n13002, Z => n13001);
   U279 : BUF_X1 port map( A => n13006, Z => n13000);
   U280 : BUF_X1 port map( A => n13005, Z => n12999);
   U281 : BUF_X1 port map( A => n13004, Z => n12998);
   U282 : BUF_X1 port map( A => n13003, Z => n12997);
   U283 : BUF_X1 port map( A => n13002, Z => n12996);
   U284 : BUF_X1 port map( A => n13163, Z => n13161);
   U285 : BUF_X1 port map( A => n13162, Z => n13160);
   U286 : BUF_X1 port map( A => n13166, Z => n13159);
   U287 : BUF_X1 port map( A => n13378, Z => n13375);
   U288 : BUF_X1 port map( A => n13378, Z => n13374);
   U289 : BUF_X1 port map( A => n13378, Z => n13373);
   U290 : BUF_X1 port map( A => n13378, Z => n13372);
   U291 : BUF_X1 port map( A => n13378, Z => n13371);
   U292 : BUF_X1 port map( A => n13374, Z => n13370);
   U293 : BUF_X1 port map( A => n13149, Z => n13142);
   U294 : BUF_X1 port map( A => n13142, Z => n13141);
   U295 : BUF_X1 port map( A => n13146, Z => n13140);
   U296 : BUF_X1 port map( A => n13145, Z => n13139);
   U297 : BUF_X1 port map( A => n13144, Z => n13138);
   U298 : BUF_X1 port map( A => n13143, Z => n13137);
   U299 : BUF_X1 port map( A => n13142, Z => n13136);
   U300 : BUF_X1 port map( A => n13119, Z => n13122);
   U301 : BUF_X1 port map( A => n13129, Z => n13121);
   U302 : BUF_X1 port map( A => n13129, Z => n13120);
   U303 : BUF_X1 port map( A => n13129, Z => n13119);
   U304 : BUF_X1 port map( A => n13129, Z => n13118);
   U305 : BUF_X1 port map( A => n13129, Z => n13117);
   U306 : BUF_X1 port map( A => n13129, Z => n13116);
   U307 : BUF_X1 port map( A => n13109, Z => n13102);
   U308 : BUF_X1 port map( A => n13102, Z => n13101);
   U309 : BUF_X1 port map( A => n13106, Z => n13100);
   U310 : BUF_X1 port map( A => n13105, Z => n13099);
   U311 : BUF_X1 port map( A => n13104, Z => n13098);
   U312 : BUF_X1 port map( A => n13103, Z => n13097);
   U313 : BUF_X1 port map( A => n13102, Z => n13096);
   U314 : BUF_X1 port map( A => n13089, Z => n13082);
   U315 : BUF_X1 port map( A => n13082, Z => n13081);
   U316 : BUF_X1 port map( A => n13086, Z => n13080);
   U317 : BUF_X1 port map( A => n13085, Z => n13079);
   U318 : BUF_X1 port map( A => n13084, Z => n13078);
   U319 : BUF_X1 port map( A => n13083, Z => n13077);
   U320 : BUF_X1 port map( A => n13082, Z => n13076);
   U321 : BUF_X1 port map( A => n13055, Z => n13062);
   U322 : BUF_X1 port map( A => n13069, Z => n13061);
   U323 : BUF_X1 port map( A => n13069, Z => n13060);
   U324 : BUF_X1 port map( A => n13069, Z => n13059);
   U325 : BUF_X1 port map( A => n13069, Z => n13058);
   U326 : BUF_X1 port map( A => n13069, Z => n13057);
   U327 : BUF_X1 port map( A => n13069, Z => n13056);
   U328 : BUF_X1 port map( A => n12861, Z => n12864);
   U329 : BUF_X1 port map( A => n12860, Z => n12863);
   U330 : BUF_X1 port map( A => n12849, Z => n12846);
   U331 : BUF_X1 port map( A => n12849, Z => n12845);
   U332 : BUF_X1 port map( A => n12849, Z => n12844);
   U333 : BUF_X1 port map( A => n12849, Z => n12843);
   U334 : BUF_X1 port map( A => n12809, Z => n12802);
   U335 : BUF_X1 port map( A => n12802, Z => n12801);
   U336 : BUF_X1 port map( A => n12806, Z => n12800);
   U337 : BUF_X1 port map( A => n12805, Z => n12799);
   U338 : BUF_X1 port map( A => n12789, Z => n12786);
   U339 : BUF_X1 port map( A => n12789, Z => n12785);
   U340 : BUF_X1 port map( A => n12789, Z => n12784);
   U341 : BUF_X1 port map( A => n12789, Z => n12783);
   U342 : BUF_X1 port map( A => n12769, Z => n12766);
   U343 : BUF_X1 port map( A => n12769, Z => n12765);
   U344 : BUF_X1 port map( A => n12769, Z => n12764);
   U345 : BUF_X1 port map( A => n12769, Z => n12763);
   U346 : BUF_X1 port map( A => n12722, Z => n12721);
   U347 : BUF_X1 port map( A => n12726, Z => n12720);
   U348 : BUF_X1 port map( A => n12725, Z => n12719);
   U349 : BUF_X1 port map( A => n12724, Z => n12718);
   U350 : BUF_X1 port map( A => n12729, Z => n12726);
   U351 : BUF_X1 port map( A => n12729, Z => n12725);
   U352 : BUF_X1 port map( A => n12855, Z => n12862);
   U353 : BUF_X1 port map( A => n12869, Z => n12861);
   U354 : BUF_X1 port map( A => n12869, Z => n12860);
   U355 : BUF_X1 port map( A => n12869, Z => n12859);
   U356 : BUF_X1 port map( A => n12869, Z => n12858);
   U357 : BUF_X1 port map( A => n12869, Z => n12857);
   U358 : BUF_X1 port map( A => n12869, Z => n12856);
   U359 : BUF_X1 port map( A => n12849, Z => n12842);
   U360 : BUF_X1 port map( A => n12842, Z => n12841);
   U361 : BUF_X1 port map( A => n12846, Z => n12840);
   U362 : BUF_X1 port map( A => n12845, Z => n12839);
   U363 : BUF_X1 port map( A => n12844, Z => n12838);
   U364 : BUF_X1 port map( A => n12843, Z => n12837);
   U365 : BUF_X1 port map( A => n12845, Z => n12836);
   U366 : BUF_X1 port map( A => n12809, Z => n12806);
   U367 : BUF_X1 port map( A => n12809, Z => n12805);
   U368 : BUF_X1 port map( A => n12809, Z => n12804);
   U369 : BUF_X1 port map( A => n12809, Z => n12803);
   U370 : BUF_X1 port map( A => n12789, Z => n12782);
   U371 : BUF_X1 port map( A => n12782, Z => n12781);
   U372 : BUF_X1 port map( A => n12786, Z => n12780);
   U373 : BUF_X1 port map( A => n12785, Z => n12779);
   U374 : BUF_X1 port map( A => n12784, Z => n12778);
   U375 : BUF_X1 port map( A => n12783, Z => n12777);
   U376 : BUF_X1 port map( A => n12785, Z => n12776);
   U377 : BUF_X1 port map( A => n12769, Z => n12762);
   U378 : BUF_X1 port map( A => n12762, Z => n12761);
   U379 : BUF_X1 port map( A => n12766, Z => n12760);
   U380 : BUF_X1 port map( A => n12765, Z => n12759);
   U381 : BUF_X1 port map( A => n12764, Z => n12758);
   U382 : BUF_X1 port map( A => n12763, Z => n12757);
   U383 : BUF_X1 port map( A => n12765, Z => n12756);
   U384 : BUF_X1 port map( A => n12729, Z => n12724);
   U385 : BUF_X1 port map( A => n12729, Z => n12723);
   U386 : BUF_X1 port map( A => n12729, Z => n12722);
   U387 : BUF_X1 port map( A => n12595, Z => n12592);
   U388 : BUF_X1 port map( A => n12595, Z => n12591);
   U389 : BUF_X1 port map( A => n12595, Z => n12590);
   U390 : BUF_X1 port map( A => n12595, Z => n12589);
   U391 : BUF_X1 port map( A => n12652, Z => n12649);
   U392 : BUF_X1 port map( A => n12652, Z => n12648);
   U393 : BUF_X1 port map( A => n12652, Z => n12647);
   U394 : BUF_X1 port map( A => n12652, Z => n12646);
   U395 : BUF_X1 port map( A => n12611, Z => n12603);
   U396 : BUF_X1 port map( A => n12610, Z => n12602);
   U397 : BUF_X1 port map( A => n12609, Z => n12601);
   U398 : BUF_X1 port map( A => n12608, Z => n12600);
   U399 : BUF_X1 port map( A => n12671, Z => n12668);
   U400 : BUF_X1 port map( A => n12671, Z => n12667);
   U401 : BUF_X1 port map( A => n12671, Z => n12666);
   U402 : BUF_X1 port map( A => n12671, Z => n12665);
   U403 : BUF_X1 port map( A => n12687, Z => n12682);
   U404 : BUF_X1 port map( A => n12686, Z => n12681);
   U405 : BUF_X1 port map( A => n12685, Z => n12680);
   U406 : BUF_X1 port map( A => n12684, Z => n12679);
   U407 : BUF_X1 port map( A => n12614, Z => n12610);
   U408 : BUF_X1 port map( A => n12595, Z => n12588);
   U409 : BUF_X1 port map( A => n12588, Z => n12587);
   U410 : BUF_X1 port map( A => n12592, Z => n12586);
   U411 : BUF_X1 port map( A => n12590, Z => n12585);
   U412 : BUF_X1 port map( A => n12589, Z => n12584);
   U413 : BUF_X1 port map( A => n12590, Z => n12583);
   U414 : BUF_X1 port map( A => n12589, Z => n12582);
   U415 : BUF_X1 port map( A => n12652, Z => n12645);
   U416 : BUF_X1 port map( A => n12645, Z => n12644);
   U417 : BUF_X1 port map( A => n12649, Z => n12643);
   U418 : BUF_X1 port map( A => n12647, Z => n12642);
   U419 : BUF_X1 port map( A => n12646, Z => n12641);
   U420 : BUF_X1 port map( A => n12647, Z => n12640);
   U421 : BUF_X1 port map( A => n12646, Z => n12639);
   U422 : BUF_X1 port map( A => n12614, Z => n12609);
   U423 : BUF_X1 port map( A => n12614, Z => n12608);
   U424 : BUF_X1 port map( A => n12614, Z => n12607);
   U425 : BUF_X1 port map( A => n12607, Z => n12606);
   U426 : BUF_X1 port map( A => n12607, Z => n12605);
   U427 : BUF_X1 port map( A => n12611, Z => n12604);
   U428 : BUF_X1 port map( A => n12671, Z => n12664);
   U429 : BUF_X1 port map( A => n12664, Z => n12663);
   U430 : BUF_X1 port map( A => n12668, Z => n12662);
   U431 : BUF_X1 port map( A => n12666, Z => n12661);
   U432 : BUF_X1 port map( A => n12665, Z => n12660);
   U433 : BUF_X1 port map( A => n12666, Z => n12659);
   U434 : BUF_X1 port map( A => n12665, Z => n12658);
   U435 : BUF_X1 port map( A => n12690, Z => n12687);
   U436 : BUF_X1 port map( A => n12690, Z => n12686);
   U437 : BUF_X1 port map( A => n12690, Z => n12685);
   U438 : BUF_X1 port map( A => n12690, Z => n12684);
   U439 : BUF_X1 port map( A => n12690, Z => n12683);
   U440 : BUF_X1 port map( A => n12926, Z => n12915);
   U441 : BUF_X1 port map( A => n12949, Z => n12935);
   U442 : BUF_X1 port map( A => n13006, Z => n12995);
   U443 : BUF_X1 port map( A => n13146, Z => n13135);
   U444 : BUF_X1 port map( A => n13129, Z => n13115);
   U445 : BUF_X1 port map( A => n13106, Z => n13095);
   U446 : BUF_X1 port map( A => n13086, Z => n13075);
   U447 : BUF_X1 port map( A => n13069, Z => n13055);
   U448 : BUF_X1 port map( A => n12869, Z => n12855);
   U449 : BUF_X1 port map( A => n12842, Z => n12835);
   U450 : BUF_X1 port map( A => n12782, Z => n12775);
   U451 : BUF_X1 port map( A => n12762, Z => n12755);
   U452 : BUF_X1 port map( A => n12591, Z => n12581);
   U453 : BUF_X1 port map( A => n12648, Z => n12638);
   U454 : BUF_X1 port map( A => n12667, Z => n12657);
   U455 : BUF_X1 port map( A => n12614, Z => n12611);
   U456 : BUF_X1 port map( A => n12633, Z => n12630);
   U457 : BUF_X1 port map( A => n12633, Z => n12629);
   U458 : BUF_X1 port map( A => n12633, Z => n12628);
   U459 : BUF_X1 port map( A => n12633, Z => n12627);
   U460 : BUF_X1 port map( A => n12633, Z => n12626);
   U461 : BUF_X1 port map( A => n12630, Z => n12625);
   U462 : BUF_X1 port map( A => n12629, Z => n12624);
   U463 : BUF_X1 port map( A => n12628, Z => n12623);
   U464 : BUF_X1 port map( A => n12627, Z => n12622);
   U465 : BUF_X1 port map( A => n12626, Z => n12621);
   U466 : BUF_X1 port map( A => n12628, Z => n12620);
   U467 : BUF_X1 port map( A => n12630, Z => n12619);
   U468 : BUF_X1 port map( A => n12683, Z => n12678);
   U469 : BUF_X1 port map( A => n12687, Z => n12677);
   U470 : BUF_X1 port map( A => n12686, Z => n12676);
   U471 : BUF_X1 port map( A => n12709, Z => n12706);
   U472 : BUF_X1 port map( A => n12709, Z => n12705);
   U473 : BUF_X1 port map( A => n12709, Z => n12704);
   U474 : BUF_X1 port map( A => n12709, Z => n12703);
   U475 : BUF_X1 port map( A => n12709, Z => n12702);
   U476 : BUF_X1 port map( A => n12706, Z => n12701);
   U477 : BUF_X1 port map( A => n12705, Z => n12700);
   U478 : BUF_X1 port map( A => n12704, Z => n12699);
   U479 : BUF_X1 port map( A => n12703, Z => n12698);
   U480 : BUF_X1 port map( A => n12702, Z => n12697);
   U481 : BUF_X1 port map( A => n12704, Z => n12696);
   U482 : BUF_X1 port map( A => n12706, Z => n12695);
   U483 : BUF_X1 port map( A => n12723, Z => n12717);
   U484 : BUF_X1 port map( A => n12722, Z => n12716);
   U485 : BUF_X1 port map( A => n12726, Z => n12715);
   U486 : BUF_X1 port map( A => n12749, Z => n12746);
   U487 : BUF_X1 port map( A => n12749, Z => n12745);
   U488 : BUF_X1 port map( A => n12749, Z => n12744);
   U489 : BUF_X1 port map( A => n12749, Z => n12743);
   U490 : BUF_X1 port map( A => n12749, Z => n12742);
   U491 : BUF_X1 port map( A => n12742, Z => n12741);
   U492 : BUF_X1 port map( A => n12746, Z => n12740);
   U493 : BUF_X1 port map( A => n12745, Z => n12739);
   U494 : BUF_X1 port map( A => n12744, Z => n12738);
   U495 : BUF_X1 port map( A => n12743, Z => n12737);
   U496 : BUF_X1 port map( A => n12745, Z => n12736);
   U497 : BUF_X1 port map( A => n12742, Z => n12735);
   U498 : BUF_X1 port map( A => n12804, Z => n12798);
   U499 : BUF_X1 port map( A => n12803, Z => n12797);
   U500 : BUF_X1 port map( A => n12805, Z => n12796);
   U501 : BUF_X1 port map( A => n12802, Z => n12795);
   U502 : BUF_X1 port map( A => n12829, Z => n12826);
   U503 : BUF_X1 port map( A => n12829, Z => n12825);
   U504 : BUF_X1 port map( A => n12829, Z => n12824);
   U505 : BUF_X1 port map( A => n12829, Z => n12823);
   U506 : BUF_X1 port map( A => n12829, Z => n12822);
   U507 : BUF_X1 port map( A => n12822, Z => n12821);
   U508 : BUF_X1 port map( A => n12826, Z => n12820);
   U509 : BUF_X1 port map( A => n12825, Z => n12819);
   U510 : BUF_X1 port map( A => n12824, Z => n12818);
   U511 : BUF_X1 port map( A => n12823, Z => n12817);
   U512 : BUF_X1 port map( A => n12825, Z => n12816);
   U513 : BUF_X1 port map( A => n12822, Z => n12815);
   U514 : BUF_X1 port map( A => n12889, Z => n12884);
   U515 : BUF_X1 port map( A => n12889, Z => n12883);
   U516 : BUF_X1 port map( A => n12889, Z => n12882);
   U517 : BUF_X1 port map( A => n12882, Z => n12881);
   U518 : BUF_X1 port map( A => n12886, Z => n12880);
   U519 : BUF_X1 port map( A => n12885, Z => n12879);
   U520 : BUF_X1 port map( A => n12884, Z => n12878);
   U521 : BUF_X1 port map( A => n12883, Z => n12877);
   U522 : BUF_X1 port map( A => n12882, Z => n12876);
   U523 : BUF_X1 port map( A => n12886, Z => n12875);
   U524 : BUF_X1 port map( A => n12909, Z => n12906);
   U525 : BUF_X1 port map( A => n12909, Z => n12905);
   U526 : BUF_X1 port map( A => n12909, Z => n12904);
   U527 : BUF_X1 port map( A => n12909, Z => n12903);
   U528 : BUF_X1 port map( A => n12909, Z => n12902);
   U529 : BUF_X1 port map( A => n12902, Z => n12901);
   U530 : BUF_X1 port map( A => n12906, Z => n12900);
   U531 : BUF_X1 port map( A => n12905, Z => n12899);
   U532 : BUF_X1 port map( A => n12904, Z => n12898);
   U533 : BUF_X1 port map( A => n12903, Z => n12897);
   U534 : BUF_X1 port map( A => n12902, Z => n12896);
   U535 : BUF_X1 port map( A => n12906, Z => n12895);
   U536 : BUF_X1 port map( A => n12969, Z => n12964);
   U537 : BUF_X1 port map( A => n12969, Z => n12963);
   U538 : BUF_X1 port map( A => n12969, Z => n12962);
   U539 : BUF_X1 port map( A => n12962, Z => n12961);
   U540 : BUF_X1 port map( A => n12966, Z => n12960);
   U541 : BUF_X1 port map( A => n12965, Z => n12959);
   U542 : BUF_X1 port map( A => n12964, Z => n12958);
   U543 : BUF_X1 port map( A => n12963, Z => n12957);
   U544 : BUF_X1 port map( A => n12962, Z => n12956);
   U545 : BUF_X1 port map( A => n12966, Z => n12955);
   U546 : BUF_X1 port map( A => n12989, Z => n12986);
   U547 : BUF_X1 port map( A => n12989, Z => n12985);
   U548 : BUF_X1 port map( A => n12989, Z => n12984);
   U549 : BUF_X1 port map( A => n12989, Z => n12983);
   U550 : BUF_X1 port map( A => n12989, Z => n12982);
   U551 : BUF_X1 port map( A => n12982, Z => n12981);
   U552 : BUF_X1 port map( A => n12986, Z => n12980);
   U553 : BUF_X1 port map( A => n12985, Z => n12979);
   U554 : BUF_X1 port map( A => n12984, Z => n12978);
   U555 : BUF_X1 port map( A => n12983, Z => n12977);
   U556 : BUF_X1 port map( A => n12982, Z => n12976);
   U557 : BUF_X1 port map( A => n12986, Z => n12975);
   U558 : BUF_X1 port map( A => n13169, Z => n13166);
   U559 : BUF_X1 port map( A => n13169, Z => n13165);
   U560 : BUF_X1 port map( A => n13169, Z => n13164);
   U561 : BUF_X1 port map( A => n13169, Z => n13163);
   U562 : BUF_X1 port map( A => n13169, Z => n13162);
   U563 : BUF_X1 port map( A => n13373, Z => n13367);
   U564 : BUF_X1 port map( A => n13372, Z => n13366);
   U565 : BUF_X1 port map( A => n13371, Z => n13365);
   U566 : BUF_X1 port map( A => n13375, Z => n13364);
   U567 : BUF_X1 port map( A => n13029, Z => n13027);
   U568 : BUF_X1 port map( A => n13049, Z => n13047);
   U569 : BUF_X1 port map( A => n13129, Z => n13127);
   U570 : BUF_X1 port map( A => n13069, Z => n13067);
   U571 : BUF_X1 port map( A => n12869, Z => n12867);
   U572 : BUF_X1 port map( A => n13019, Z => n13025);
   U573 : BUF_X1 port map( A => n13039, Z => n13045);
   U574 : BUF_X1 port map( A => n12935, Z => n12946);
   U575 : BUF_X1 port map( A => n13118, Z => n13125);
   U576 : BUF_X1 port map( A => n13059, Z => n13065);
   U577 : BUF_X1 port map( A => n12859, Z => n12865);
   U578 : BUF_X1 port map( A => n13029, Z => n13028);
   U579 : BUF_X1 port map( A => n13049, Z => n13048);
   U580 : BUF_X1 port map( A => n12614, Z => n12613);
   U581 : BUF_X1 port map( A => n12929, Z => n12928);
   U582 : BUF_X1 port map( A => n12949, Z => n12948);
   U583 : BUF_X1 port map( A => n13009, Z => n13008);
   U584 : BUF_X1 port map( A => n13149, Z => n13148);
   U585 : BUF_X1 port map( A => n13129, Z => n13128);
   U586 : BUF_X1 port map( A => n13109, Z => n13108);
   U587 : BUF_X1 port map( A => n13089, Z => n13088);
   U588 : BUF_X1 port map( A => n13069, Z => n13068);
   U589 : BUF_X1 port map( A => n12869, Z => n12868);
   U590 : BUF_X1 port map( A => n12849, Z => n12848);
   U591 : BUF_X1 port map( A => n12789, Z => n12788);
   U592 : BUF_X1 port map( A => n12769, Z => n12768);
   U593 : BUF_X1 port map( A => n12595, Z => n12594);
   U594 : BUF_X1 port map( A => n12652, Z => n12651);
   U595 : BUF_X1 port map( A => n12671, Z => n12670);
   U596 : BUF_X1 port map( A => n12633, Z => n12632);
   U597 : BUF_X1 port map( A => n12690, Z => n12689);
   U598 : BUF_X1 port map( A => n12709, Z => n12708);
   U599 : BUF_X1 port map( A => n12729, Z => n12728);
   U600 : BUF_X1 port map( A => n12749, Z => n12748);
   U601 : BUF_X1 port map( A => n12809, Z => n12808);
   U602 : BUF_X1 port map( A => n12829, Z => n12828);
   U603 : BUF_X1 port map( A => n12889, Z => n12888);
   U604 : BUF_X1 port map( A => n12909, Z => n12908);
   U605 : BUF_X1 port map( A => n12969, Z => n12968);
   U606 : BUF_X1 port map( A => n12989, Z => n12988);
   U607 : BUF_X1 port map( A => n13169, Z => n13168);
   U608 : BUF_X1 port map( A => n13378, Z => n13377);
   U609 : BUF_X1 port map( A => n12939, Z => n12945);
   U610 : BUF_X1 port map( A => n13018, Z => n13026);
   U611 : BUF_X1 port map( A => n13038, Z => n13046);
   U612 : BUF_X1 port map( A => n12938, Z => n12943);
   U613 : BUF_X1 port map( A => n13117, Z => n13126);
   U614 : BUF_X1 port map( A => n13058, Z => n13066);
   U615 : BUF_X1 port map( A => n12858, Z => n12866);
   U616 : INV_X1 port map( A => n12550, ZN => n12574);
   U617 : INV_X1 port map( A => n12550, ZN => n12575);
   U618 : INV_X1 port map( A => n12550, ZN => n12576);
   U619 : BUF_X1 port map( A => n1982, Z => n12435);
   U620 : BUF_X1 port map( A => n1987, Z => n12411);
   U621 : BUF_X1 port map( A => n1982, Z => n12436);
   U622 : BUF_X1 port map( A => n1987, Z => n12412);
   U623 : BUF_X1 port map( A => n1982, Z => n12437);
   U624 : BUF_X1 port map( A => n1987, Z => n12413);
   U625 : BUF_X1 port map( A => n1982, Z => n12438);
   U626 : BUF_X1 port map( A => n1987, Z => n12414);
   U627 : BUF_X1 port map( A => n1982, Z => n12439);
   U628 : BUF_X1 port map( A => n1987, Z => n12415);
   U629 : BUF_X1 port map( A => n1992, Z => n12387);
   U630 : BUF_X1 port map( A => n1997, Z => n12363);
   U631 : BUF_X1 port map( A => n1958, Z => n12531);
   U632 : BUF_X1 port map( A => n1963, Z => n12507);
   U633 : BUF_X1 port map( A => n1968, Z => n12483);
   U634 : BUF_X1 port map( A => n1973, Z => n12459);
   U635 : BUF_X1 port map( A => n1992, Z => n12388);
   U636 : BUF_X1 port map( A => n1997, Z => n12364);
   U637 : BUF_X1 port map( A => n1958, Z => n12532);
   U638 : BUF_X1 port map( A => n1963, Z => n12508);
   U639 : BUF_X1 port map( A => n1968, Z => n12484);
   U640 : BUF_X1 port map( A => n1973, Z => n12460);
   U641 : BUF_X1 port map( A => n1992, Z => n12389);
   U642 : BUF_X1 port map( A => n1997, Z => n12365);
   U643 : BUF_X1 port map( A => n1958, Z => n12533);
   U644 : BUF_X1 port map( A => n1963, Z => n12509);
   U645 : BUF_X1 port map( A => n1968, Z => n12485);
   U646 : BUF_X1 port map( A => n1973, Z => n12461);
   U647 : BUF_X1 port map( A => n1992, Z => n12390);
   U648 : BUF_X1 port map( A => n1997, Z => n12366);
   U649 : BUF_X1 port map( A => n1958, Z => n12534);
   U650 : BUF_X1 port map( A => n1963, Z => n12510);
   U651 : BUF_X1 port map( A => n1968, Z => n12486);
   U652 : BUF_X1 port map( A => n1973, Z => n12462);
   U653 : BUF_X1 port map( A => n1992, Z => n12391);
   U654 : BUF_X1 port map( A => n1997, Z => n12367);
   U655 : BUF_X1 port map( A => n1958, Z => n12535);
   U656 : BUF_X1 port map( A => n1963, Z => n12511);
   U657 : BUF_X1 port map( A => n1968, Z => n12487);
   U658 : BUF_X1 port map( A => n1973, Z => n12463);
   U659 : BUF_X1 port map( A => n1983, Z => n12429);
   U660 : BUF_X1 port map( A => n1988, Z => n12405);
   U661 : BUF_X1 port map( A => n1993, Z => n12381);
   U662 : BUF_X1 port map( A => n1959, Z => n12525);
   U663 : BUF_X1 port map( A => n1964, Z => n12501);
   U664 : BUF_X1 port map( A => n1969, Z => n12477);
   U665 : BUF_X1 port map( A => n1974, Z => n12453);
   U666 : BUF_X1 port map( A => n1983, Z => n12430);
   U667 : BUF_X1 port map( A => n1988, Z => n12406);
   U668 : BUF_X1 port map( A => n1993, Z => n12382);
   U669 : BUF_X1 port map( A => n1959, Z => n12526);
   U670 : BUF_X1 port map( A => n1964, Z => n12502);
   U671 : BUF_X1 port map( A => n1969, Z => n12478);
   U672 : BUF_X1 port map( A => n1974, Z => n12454);
   U673 : BUF_X1 port map( A => n1983, Z => n12431);
   U674 : BUF_X1 port map( A => n1988, Z => n12407);
   U675 : BUF_X1 port map( A => n1993, Z => n12383);
   U676 : BUF_X1 port map( A => n1959, Z => n12527);
   U677 : BUF_X1 port map( A => n1964, Z => n12503);
   U678 : BUF_X1 port map( A => n1969, Z => n12479);
   U679 : BUF_X1 port map( A => n1974, Z => n12455);
   U680 : BUF_X1 port map( A => n1983, Z => n12432);
   U681 : BUF_X1 port map( A => n1988, Z => n12408);
   U682 : BUF_X1 port map( A => n1993, Z => n12384);
   U683 : BUF_X1 port map( A => n1959, Z => n12528);
   U684 : BUF_X1 port map( A => n1964, Z => n12504);
   U685 : BUF_X1 port map( A => n1969, Z => n12480);
   U686 : BUF_X1 port map( A => n1974, Z => n12456);
   U687 : BUF_X1 port map( A => n1983, Z => n12433);
   U688 : BUF_X1 port map( A => n1988, Z => n12409);
   U689 : BUF_X1 port map( A => n1993, Z => n12385);
   U690 : BUF_X1 port map( A => n1959, Z => n12529);
   U691 : BUF_X1 port map( A => n1964, Z => n12505);
   U692 : BUF_X1 port map( A => n1969, Z => n12481);
   U693 : BUF_X1 port map( A => n1974, Z => n12457);
   U694 : BUF_X1 port map( A => n1995, Z => n12375);
   U695 : BUF_X1 port map( A => n2000, Z => n12351);
   U696 : BUF_X1 port map( A => n1961, Z => n12519);
   U697 : BUF_X1 port map( A => n1966, Z => n12495);
   U698 : BUF_X1 port map( A => n1995, Z => n12376);
   U699 : BUF_X1 port map( A => n2000, Z => n12352);
   U700 : BUF_X1 port map( A => n1961, Z => n12520);
   U701 : BUF_X1 port map( A => n1966, Z => n12496);
   U702 : BUF_X1 port map( A => n1995, Z => n12377);
   U703 : BUF_X1 port map( A => n2000, Z => n12353);
   U704 : BUF_X1 port map( A => n1961, Z => n12521);
   U705 : BUF_X1 port map( A => n1966, Z => n12497);
   U706 : BUF_X1 port map( A => n1995, Z => n12378);
   U707 : BUF_X1 port map( A => n2000, Z => n12354);
   U708 : BUF_X1 port map( A => n1961, Z => n12522);
   U709 : BUF_X1 port map( A => n1966, Z => n12498);
   U710 : BUF_X1 port map( A => n1995, Z => n12379);
   U711 : BUF_X1 port map( A => n2000, Z => n12355);
   U712 : BUF_X1 port map( A => n1961, Z => n12523);
   U713 : BUF_X1 port map( A => n1966, Z => n12499);
   U714 : BUF_X1 port map( A => n1985, Z => n12423);
   U715 : BUF_X1 port map( A => n1990, Z => n12399);
   U716 : BUF_X1 port map( A => n1971, Z => n12471);
   U717 : BUF_X1 port map( A => n1976, Z => n12447);
   U718 : BUF_X1 port map( A => n1985, Z => n12424);
   U719 : BUF_X1 port map( A => n1990, Z => n12400);
   U720 : BUF_X1 port map( A => n1971, Z => n12472);
   U721 : BUF_X1 port map( A => n1976, Z => n12448);
   U722 : BUF_X1 port map( A => n1985, Z => n12425);
   U723 : BUF_X1 port map( A => n1990, Z => n12401);
   U724 : BUF_X1 port map( A => n1971, Z => n12473);
   U725 : BUF_X1 port map( A => n1976, Z => n12449);
   U726 : BUF_X1 port map( A => n1985, Z => n12426);
   U727 : BUF_X1 port map( A => n1990, Z => n12402);
   U728 : BUF_X1 port map( A => n1971, Z => n12474);
   U729 : BUF_X1 port map( A => n1976, Z => n12450);
   U730 : BUF_X1 port map( A => n1985, Z => n12427);
   U731 : BUF_X1 port map( A => n1990, Z => n12403);
   U732 : BUF_X1 port map( A => n1971, Z => n12475);
   U733 : BUF_X1 port map( A => n1976, Z => n12451);
   U734 : BUF_X1 port map( A => n1986, Z => n12417);
   U735 : BUF_X1 port map( A => n1991, Z => n12393);
   U736 : BUF_X1 port map( A => n1986, Z => n12418);
   U737 : BUF_X1 port map( A => n1991, Z => n12394);
   U738 : BUF_X1 port map( A => n1986, Z => n12419);
   U739 : BUF_X1 port map( A => n1991, Z => n12395);
   U740 : BUF_X1 port map( A => n1986, Z => n12420);
   U741 : BUF_X1 port map( A => n1991, Z => n12396);
   U742 : BUF_X1 port map( A => n1986, Z => n12421);
   U743 : BUF_X1 port map( A => n1991, Z => n12397);
   U744 : BUF_X1 port map( A => n1996, Z => n12369);
   U745 : BUF_X1 port map( A => n2001, Z => n12345);
   U746 : BUF_X1 port map( A => n1962, Z => n12513);
   U747 : BUF_X1 port map( A => n1967, Z => n12489);
   U748 : BUF_X1 port map( A => n1996, Z => n12370);
   U749 : BUF_X1 port map( A => n2001, Z => n12346);
   U750 : BUF_X1 port map( A => n1962, Z => n12514);
   U751 : BUF_X1 port map( A => n1967, Z => n12490);
   U752 : BUF_X1 port map( A => n1996, Z => n12371);
   U753 : BUF_X1 port map( A => n2001, Z => n12347);
   U754 : BUF_X1 port map( A => n1962, Z => n12515);
   U755 : BUF_X1 port map( A => n1967, Z => n12491);
   U756 : BUF_X1 port map( A => n1996, Z => n12372);
   U757 : BUF_X1 port map( A => n2001, Z => n12348);
   U758 : BUF_X1 port map( A => n1962, Z => n12516);
   U759 : BUF_X1 port map( A => n1967, Z => n12492);
   U760 : BUF_X1 port map( A => n1996, Z => n12373);
   U761 : BUF_X1 port map( A => n2001, Z => n12349);
   U762 : BUF_X1 port map( A => n1962, Z => n12517);
   U763 : BUF_X1 port map( A => n1967, Z => n12493);
   U764 : BUF_X1 port map( A => n1972, Z => n12465);
   U765 : BUF_X1 port map( A => n1977, Z => n12441);
   U766 : BUF_X1 port map( A => n1972, Z => n12466);
   U767 : BUF_X1 port map( A => n1977, Z => n12442);
   U768 : BUF_X1 port map( A => n1972, Z => n12467);
   U769 : BUF_X1 port map( A => n1977, Z => n12443);
   U770 : BUF_X1 port map( A => n1972, Z => n12468);
   U771 : BUF_X1 port map( A => n1977, Z => n12444);
   U772 : BUF_X1 port map( A => n1972, Z => n12469);
   U773 : BUF_X1 port map( A => n1977, Z => n12445);
   U774 : AND2_X1 port map( A1 => n3209, A2 => n3194, ZN => n1998);
   U775 : BUF_X1 port map( A => n1949, Z => n12550);
   U776 : INV_X1 port map( A => n13030, ZN => n13049);
   U777 : INV_X1 port map( A => n13010, ZN => n13029);
   U778 : INV_X1 port map( A => n12577, ZN => n12595);
   U779 : INV_X1 port map( A => n12910, ZN => n12929);
   U780 : INV_X1 port map( A => n12830, ZN => n12849);
   U781 : INV_X1 port map( A => n12790, ZN => n12809);
   U782 : INV_X1 port map( A => n12770, ZN => n12789);
   U783 : INV_X1 port map( A => n12750, ZN => n12769);
   U784 : INV_X1 port map( A => n12710, ZN => n12729);
   U785 : INV_X1 port map( A => n12730, ZN => n12749);
   U786 : INV_X1 port map( A => n12810, ZN => n12829);
   U787 : INV_X1 port map( A => n12850, ZN => n12869);
   U788 : INV_X1 port map( A => n13359, ZN => n13378);
   U789 : INV_X1 port map( A => n13130, ZN => n13149);
   U790 : INV_X1 port map( A => n13090, ZN => n13109);
   U791 : INV_X1 port map( A => n13070, ZN => n13089);
   U792 : INV_X1 port map( A => n13150, ZN => n13169);
   U793 : INV_X1 port map( A => n13110, ZN => n13129);
   U794 : INV_X1 port map( A => n13050, ZN => n13069);
   U795 : INV_X1 port map( A => n12990, ZN => n13009);
   U796 : INV_X1 port map( A => n12930, ZN => n12949);
   U797 : INV_X1 port map( A => n12634, ZN => n12652);
   U798 : INV_X1 port map( A => n12653, ZN => n12671);
   U799 : INV_X1 port map( A => n12672, ZN => n12690);
   U800 : INV_X1 port map( A => n12596, ZN => n12614);
   U801 : INV_X1 port map( A => n12615, ZN => n12633);
   U802 : INV_X1 port map( A => n12691, ZN => n12709);
   U803 : INV_X1 port map( A => n12870, ZN => n12889);
   U804 : INV_X1 port map( A => n12890, ZN => n12909);
   U805 : INV_X1 port map( A => n12950, ZN => n12969);
   U806 : INV_X1 port map( A => n12970, ZN => n12989);
   U807 : BUF_X1 port map( A => n3259, Z => n12152);
   U808 : BUF_X1 port map( A => n3259, Z => n12153);
   U809 : BUF_X1 port map( A => n3259, Z => n12154);
   U810 : BUF_X1 port map( A => n3259, Z => n12155);
   U811 : BUF_X1 port map( A => n3259, Z => n12156);
   U812 : NOR2_X1 port map( A1 => n14463, A2 => n14464, ZN => n3194);
   U813 : NOR3_X1 port map( A1 => n14465, A2 => n14461, A3 => n14462, ZN => 
                           n3209);
   U814 : NAND2_X1 port map( A1 => n3189, A2 => n3205, ZN => n1985);
   U815 : NAND2_X1 port map( A1 => n3193, A2 => n3205, ZN => n1990);
   U816 : NAND2_X1 port map( A1 => n3208, A2 => n3189, ZN => n1996);
   U817 : NAND2_X1 port map( A1 => n3190, A2 => n3189, ZN => n1961);
   U818 : NAND2_X1 port map( A1 => n3188, A2 => n3189, ZN => n1962);
   U819 : NAND2_X1 port map( A1 => n3209, A2 => n3193, ZN => n2000);
   U820 : NAND2_X1 port map( A1 => n3208, A2 => n3193, ZN => n2001);
   U821 : NAND2_X1 port map( A1 => n3190, A2 => n3193, ZN => n1966);
   U822 : NAND2_X1 port map( A1 => n3188, A2 => n3193, ZN => n1967);
   U823 : NAND2_X1 port map( A1 => n3197, A2 => n3194, ZN => n1976);
   U824 : NAND2_X1 port map( A1 => n3196, A2 => n3194, ZN => n1977);
   U825 : NAND2_X1 port map( A1 => n3197, A2 => n3191, ZN => n1971);
   U826 : NAND2_X1 port map( A1 => n3196, A2 => n3191, ZN => n1972);
   U827 : OAI21_X1 port map( B1 => n1921, B2 => n1942, A => n12137, ZN => n1949
                           );
   U828 : AND2_X1 port map( A1 => n3205, A2 => n3191, ZN => n1983);
   U829 : AND2_X1 port map( A1 => n3194, A2 => n3205, ZN => n1988);
   U830 : AND2_X1 port map( A1 => n3208, A2 => n3191, ZN => n1992);
   U831 : AND2_X1 port map( A1 => n3208, A2 => n3194, ZN => n1997);
   U832 : AND2_X1 port map( A1 => n3188, A2 => n3191, ZN => n1958);
   U833 : AND2_X1 port map( A1 => n3190, A2 => n3191, ZN => n1959);
   U834 : AND2_X1 port map( A1 => n3188, A2 => n3194, ZN => n1963);
   U835 : AND2_X1 port map( A1 => n3190, A2 => n3194, ZN => n1964);
   U836 : AND2_X1 port map( A1 => n3196, A2 => n3189, ZN => n1968);
   U837 : AND2_X1 port map( A1 => n3197, A2 => n3189, ZN => n1969);
   U838 : AND2_X1 port map( A1 => n3196, A2 => n3193, ZN => n1973);
   U839 : AND2_X1 port map( A1 => n3197, A2 => n3193, ZN => n1974);
   U840 : AND2_X1 port map( A1 => n3209, A2 => n3191, ZN => n1993);
   U841 : OAI21_X1 port map( B1 => n1919, B2 => n1942, A => n12137, ZN => n1948
                           );
   U842 : OAI21_X1 port map( B1 => n1913, B2 => n1942, A => n12137, ZN => n1945
                           );
   U843 : OAI21_X1 port map( B1 => n1911, B2 => n1942, A => n12137, ZN => n1944
                           );
   U844 : OAI21_X1 port map( B1 => n1917, B2 => n1942, A => n12137, ZN => n1947
                           );
   U845 : OAI21_X1 port map( B1 => n1915, B2 => n1942, A => n12137, ZN => n1946
                           );
   U846 : OAI21_X1 port map( B1 => n1909, B2 => n1942, A => n12137, ZN => n1943
                           );
   U847 : OAI21_X1 port map( B1 => n1907, B2 => n1942, A => n12137, ZN => n1941
                           );
   U848 : OAI21_X1 port map( B1 => n1917, B2 => n1924, A => n12138, ZN => n1929
                           );
   U849 : OAI21_X1 port map( B1 => n1921, B2 => n1924, A => n12138, ZN => n1931
                           );
   U850 : OAI21_X1 port map( B1 => n1919, B2 => n1924, A => n12138, ZN => n1930
                           );
   U851 : OAI21_X1 port map( B1 => n1913, B2 => n1924, A => n12138, ZN => n1927
                           );
   U852 : OAI21_X1 port map( B1 => n1911, B2 => n1924, A => n12139, ZN => n1926
                           );
   U853 : BUF_X1 port map( A => n3219, Z => n12326);
   U854 : BUF_X1 port map( A => n3224, Z => n12302);
   U855 : BUF_X1 port map( A => n3229, Z => n12278);
   U856 : BUF_X1 port map( A => n3234, Z => n12254);
   U857 : BUF_X1 port map( A => n3243, Z => n12230);
   U858 : BUF_X1 port map( A => n3248, Z => n12206);
   U859 : BUF_X1 port map( A => n3253, Z => n12182);
   U860 : BUF_X1 port map( A => n3258, Z => n12158);
   U861 : BUF_X1 port map( A => n3219, Z => n12327);
   U862 : BUF_X1 port map( A => n3224, Z => n12303);
   U863 : BUF_X1 port map( A => n3229, Z => n12279);
   U864 : BUF_X1 port map( A => n3234, Z => n12255);
   U865 : BUF_X1 port map( A => n3243, Z => n12231);
   U866 : BUF_X1 port map( A => n3248, Z => n12207);
   U867 : BUF_X1 port map( A => n3253, Z => n12183);
   U868 : BUF_X1 port map( A => n3258, Z => n12159);
   U869 : BUF_X1 port map( A => n3219, Z => n12328);
   U870 : BUF_X1 port map( A => n3224, Z => n12304);
   U871 : BUF_X1 port map( A => n3229, Z => n12280);
   U872 : BUF_X1 port map( A => n3234, Z => n12256);
   U873 : BUF_X1 port map( A => n3243, Z => n12232);
   U874 : BUF_X1 port map( A => n3248, Z => n12208);
   U875 : BUF_X1 port map( A => n3253, Z => n12184);
   U876 : BUF_X1 port map( A => n3258, Z => n12160);
   U877 : BUF_X1 port map( A => n3219, Z => n12329);
   U878 : BUF_X1 port map( A => n3224, Z => n12305);
   U879 : BUF_X1 port map( A => n3229, Z => n12281);
   U880 : BUF_X1 port map( A => n3234, Z => n12257);
   U881 : BUF_X1 port map( A => n3243, Z => n12233);
   U882 : BUF_X1 port map( A => n3248, Z => n12209);
   U883 : BUF_X1 port map( A => n3253, Z => n12185);
   U884 : BUF_X1 port map( A => n3258, Z => n12161);
   U885 : BUF_X1 port map( A => n3219, Z => n12330);
   U886 : BUF_X1 port map( A => n3224, Z => n12306);
   U887 : BUF_X1 port map( A => n3229, Z => n12282);
   U888 : BUF_X1 port map( A => n3234, Z => n12258);
   U889 : BUF_X1 port map( A => n3243, Z => n12234);
   U890 : BUF_X1 port map( A => n3248, Z => n12210);
   U891 : BUF_X1 port map( A => n3253, Z => n12186);
   U892 : BUF_X1 port map( A => n3258, Z => n12162);
   U893 : BUF_X1 port map( A => n3220, Z => n12320);
   U894 : BUF_X1 port map( A => n3225, Z => n12296);
   U895 : BUF_X1 port map( A => n3230, Z => n12272);
   U896 : BUF_X1 port map( A => n3235, Z => n12248);
   U897 : BUF_X1 port map( A => n3244, Z => n12224);
   U898 : BUF_X1 port map( A => n3249, Z => n12200);
   U899 : BUF_X1 port map( A => n3254, Z => n12176);
   U900 : BUF_X1 port map( A => n3220, Z => n12321);
   U901 : BUF_X1 port map( A => n3225, Z => n12297);
   U902 : BUF_X1 port map( A => n3230, Z => n12273);
   U903 : BUF_X1 port map( A => n3235, Z => n12249);
   U904 : BUF_X1 port map( A => n3244, Z => n12225);
   U905 : BUF_X1 port map( A => n3249, Z => n12201);
   U906 : BUF_X1 port map( A => n3254, Z => n12177);
   U907 : BUF_X1 port map( A => n3220, Z => n12322);
   U908 : BUF_X1 port map( A => n3225, Z => n12298);
   U909 : BUF_X1 port map( A => n3230, Z => n12274);
   U910 : BUF_X1 port map( A => n3235, Z => n12250);
   U911 : BUF_X1 port map( A => n3244, Z => n12226);
   U912 : BUF_X1 port map( A => n3249, Z => n12202);
   U913 : BUF_X1 port map( A => n3254, Z => n12178);
   U914 : BUF_X1 port map( A => n3220, Z => n12323);
   U915 : BUF_X1 port map( A => n3225, Z => n12299);
   U916 : BUF_X1 port map( A => n3230, Z => n12275);
   U917 : BUF_X1 port map( A => n3235, Z => n12251);
   U918 : BUF_X1 port map( A => n3244, Z => n12227);
   U919 : BUF_X1 port map( A => n3249, Z => n12203);
   U920 : BUF_X1 port map( A => n3254, Z => n12179);
   U921 : BUF_X1 port map( A => n3220, Z => n12324);
   U922 : BUF_X1 port map( A => n3225, Z => n12300);
   U923 : BUF_X1 port map( A => n3230, Z => n12276);
   U924 : BUF_X1 port map( A => n3235, Z => n12252);
   U925 : BUF_X1 port map( A => n3244, Z => n12228);
   U926 : BUF_X1 port map( A => n3249, Z => n12204);
   U927 : BUF_X1 port map( A => n3254, Z => n12180);
   U928 : BUF_X1 port map( A => n3222, Z => n12314);
   U929 : BUF_X1 port map( A => n3227, Z => n12290);
   U930 : BUF_X1 port map( A => n3256, Z => n12170);
   U931 : BUF_X1 port map( A => n3261, Z => n12146);
   U932 : BUF_X1 port map( A => n3222, Z => n12315);
   U933 : BUF_X1 port map( A => n3227, Z => n12291);
   U934 : BUF_X1 port map( A => n3256, Z => n12171);
   U935 : BUF_X1 port map( A => n3261, Z => n12147);
   U936 : BUF_X1 port map( A => n3222, Z => n12316);
   U937 : BUF_X1 port map( A => n3227, Z => n12292);
   U938 : BUF_X1 port map( A => n3256, Z => n12172);
   U939 : BUF_X1 port map( A => n3261, Z => n12148);
   U940 : BUF_X1 port map( A => n3222, Z => n12317);
   U941 : BUF_X1 port map( A => n3227, Z => n12293);
   U942 : BUF_X1 port map( A => n3256, Z => n12173);
   U943 : BUF_X1 port map( A => n3261, Z => n12149);
   U944 : BUF_X1 port map( A => n3222, Z => n12318);
   U945 : BUF_X1 port map( A => n3227, Z => n12294);
   U946 : BUF_X1 port map( A => n3256, Z => n12174);
   U947 : BUF_X1 port map( A => n3261, Z => n12150);
   U948 : BUF_X1 port map( A => n3232, Z => n12266);
   U949 : BUF_X1 port map( A => n3246, Z => n12218);
   U950 : BUF_X1 port map( A => n3251, Z => n12194);
   U951 : BUF_X1 port map( A => n3232, Z => n12267);
   U952 : BUF_X1 port map( A => n3246, Z => n12219);
   U953 : BUF_X1 port map( A => n3251, Z => n12195);
   U954 : BUF_X1 port map( A => n3232, Z => n12268);
   U955 : BUF_X1 port map( A => n3246, Z => n12220);
   U956 : BUF_X1 port map( A => n3251, Z => n12196);
   U957 : BUF_X1 port map( A => n3232, Z => n12269);
   U958 : BUF_X1 port map( A => n3246, Z => n12221);
   U959 : BUF_X1 port map( A => n3251, Z => n12197);
   U960 : BUF_X1 port map( A => n3232, Z => n12270);
   U961 : BUF_X1 port map( A => n3246, Z => n12222);
   U962 : BUF_X1 port map( A => n3251, Z => n12198);
   U963 : BUF_X1 port map( A => n3237, Z => n12242);
   U964 : BUF_X1 port map( A => n3237, Z => n12243);
   U965 : BUF_X1 port map( A => n3237, Z => n12244);
   U966 : BUF_X1 port map( A => n3237, Z => n12245);
   U967 : BUF_X1 port map( A => n3237, Z => n12246);
   U968 : BUF_X1 port map( A => n3223, Z => n12308);
   U969 : BUF_X1 port map( A => n3228, Z => n12284);
   U970 : BUF_X1 port map( A => n3257, Z => n12164);
   U971 : BUF_X1 port map( A => n3262, Z => n12140);
   U972 : BUF_X1 port map( A => n3223, Z => n12309);
   U973 : BUF_X1 port map( A => n3228, Z => n12285);
   U974 : BUF_X1 port map( A => n3257, Z => n12165);
   U975 : BUF_X1 port map( A => n3262, Z => n12141);
   U976 : BUF_X1 port map( A => n3223, Z => n12310);
   U977 : BUF_X1 port map( A => n3228, Z => n12286);
   U978 : BUF_X1 port map( A => n3257, Z => n12166);
   U979 : BUF_X1 port map( A => n3262, Z => n12142);
   U980 : BUF_X1 port map( A => n3223, Z => n12311);
   U981 : BUF_X1 port map( A => n3228, Z => n12287);
   U982 : BUF_X1 port map( A => n3257, Z => n12167);
   U983 : BUF_X1 port map( A => n3262, Z => n12143);
   U984 : BUF_X1 port map( A => n3223, Z => n12312);
   U985 : BUF_X1 port map( A => n3228, Z => n12288);
   U986 : BUF_X1 port map( A => n3257, Z => n12168);
   U987 : BUF_X1 port map( A => n3262, Z => n12144);
   U988 : BUF_X1 port map( A => n3233, Z => n12260);
   U989 : BUF_X1 port map( A => n3247, Z => n12212);
   U990 : BUF_X1 port map( A => n3252, Z => n12188);
   U991 : BUF_X1 port map( A => n3233, Z => n12261);
   U992 : BUF_X1 port map( A => n3247, Z => n12213);
   U993 : BUF_X1 port map( A => n3252, Z => n12189);
   U994 : BUF_X1 port map( A => n3233, Z => n12262);
   U995 : BUF_X1 port map( A => n3247, Z => n12214);
   U996 : BUF_X1 port map( A => n3252, Z => n12190);
   U997 : BUF_X1 port map( A => n3233, Z => n12263);
   U998 : BUF_X1 port map( A => n3247, Z => n12215);
   U999 : BUF_X1 port map( A => n3252, Z => n12191);
   U1000 : BUF_X1 port map( A => n3233, Z => n12264);
   U1001 : BUF_X1 port map( A => n3247, Z => n12216);
   U1002 : BUF_X1 port map( A => n3252, Z => n12192);
   U1003 : BUF_X1 port map( A => n3238, Z => n12236);
   U1004 : BUF_X1 port map( A => n3238, Z => n12237);
   U1005 : BUF_X1 port map( A => n3238, Z => n12238);
   U1006 : BUF_X1 port map( A => n3238, Z => n12239);
   U1007 : BUF_X1 port map( A => n3238, Z => n12240);
   U1008 : BUF_X1 port map( A => n12332, Z => n12338);
   U1009 : BUF_X1 port map( A => n12332, Z => n12337);
   U1010 : BUF_X1 port map( A => n12332, Z => n12335);
   U1011 : BUF_X1 port map( A => n12332, Z => n12334);
   U1012 : BUF_X1 port map( A => n12332, Z => n12336);
   U1013 : BUF_X1 port map( A => n12332, Z => n12339);
   U1014 : BUF_X1 port map( A => n12333, Z => n12340);
   U1015 : BUF_X1 port map( A => n12333, Z => n12341);
   U1016 : BUF_X1 port map( A => n12333, Z => n12342);
   U1017 : BUF_X1 port map( A => n12333, Z => n12343);
   U1018 : AND2_X1 port map( A1 => n4470, A2 => n4455, ZN => n3259);
   U1019 : BUF_X1 port map( A => n12130, Z => n12137);
   U1020 : BUF_X1 port map( A => n12130, Z => n12136);
   U1021 : BUF_X1 port map( A => n12129, Z => n12134);
   U1022 : BUF_X1 port map( A => n12130, Z => n12135);
   U1023 : BUF_X1 port map( A => n12129, Z => n12133);
   U1024 : BUF_X1 port map( A => n12129, Z => n12132);
   U1025 : BUF_X1 port map( A => n12537, Z => n12543);
   U1026 : BUF_X1 port map( A => n12537, Z => n12542);
   U1027 : BUF_X1 port map( A => n12537, Z => n12540);
   U1028 : BUF_X1 port map( A => n12537, Z => n12539);
   U1029 : BUF_X1 port map( A => n12537, Z => n12541);
   U1030 : BUF_X1 port map( A => n12537, Z => n12544);
   U1031 : BUF_X1 port map( A => n12538, Z => n12545);
   U1032 : BUF_X1 port map( A => n12538, Z => n12546);
   U1033 : BUF_X1 port map( A => n12538, Z => n12547);
   U1034 : BUF_X1 port map( A => n12538, Z => n12548);
   U1035 : BUF_X1 port map( A => n12131, Z => n12138);
   U1036 : BUF_X1 port map( A => n12131, Z => n12139);
   U1037 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n3189);
   U1038 : NOR2_X1 port map( A1 => n14463, A2 => ADD_RD1(1), ZN => n3193);
   U1039 : NOR3_X1 port map( A1 => n14461, A2 => ADD_RD1(3), A3 => n14465, ZN 
                           => n3205);
   U1040 : NOR2_X1 port map( A1 => n14464, A2 => ADD_RD1(2), ZN => n3191);
   U1041 : NOR3_X1 port map( A1 => n14461, A2 => ADD_RD1(0), A3 => n14462, ZN 
                           => n3208);
   U1042 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n14465, 
                           ZN => n3188);
   U1043 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n3190);
   U1044 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n14462, 
                           ZN => n3196);
   U1045 : NOR3_X1 port map( A1 => n14465, A2 => ADD_RD1(4), A3 => n14462, ZN 
                           => n3197);
   U1046 : AOI221_X1 port map( B1 => n12507, B2 => n11586, C1 => n12501, C2 => 
                           n11406, A => n3192, ZN => n3185);
   U1047 : OAI22_X1 port map( A1 => n14362, A2 => n12495, B1 => n14361, B2 => 
                           n12489, ZN => n3192);
   U1048 : AOI221_X1 port map( B1 => n12507, B2 => n11762, C1 => n12501, C2 => 
                           n11582, A => n3169, ZN => n3166);
   U1049 : OAI22_X1 port map( A1 => n14408, A2 => n12495, B1 => n14385, B2 => 
                           n12489, ZN => n3169);
   U1050 : AOI221_X1 port map( B1 => n12507, B2 => n11587, C1 => n12501, C2 => 
                           n11407, A => n3150, ZN => n3147);
   U1051 : OAI22_X1 port map( A1 => n14407, A2 => n12495, B1 => n14384, B2 => 
                           n12489, ZN => n3150);
   U1052 : AOI221_X1 port map( B1 => n12507, B2 => n11588, C1 => n12501, C2 => 
                           n11408, A => n3131, ZN => n3128);
   U1053 : OAI22_X1 port map( A1 => n14406, A2 => n12495, B1 => n14383, B2 => 
                           n12489, ZN => n3131);
   U1054 : AOI221_X1 port map( B1 => n12507, B2 => n11589, C1 => n12501, C2 => 
                           n11409, A => n3112, ZN => n3109);
   U1055 : OAI22_X1 port map( A1 => n14405, A2 => n12495, B1 => n14382, B2 => 
                           n12489, ZN => n3112);
   U1056 : AOI221_X1 port map( B1 => n12507, B2 => n11763, C1 => n12501, C2 => 
                           n11583, A => n3093, ZN => n3090);
   U1057 : OAI22_X1 port map( A1 => n14404, A2 => n12495, B1 => n14381, B2 => 
                           n12489, ZN => n3093);
   U1058 : AOI221_X1 port map( B1 => n12507, B2 => n11764, C1 => n12501, C2 => 
                           n11584, A => n3074, ZN => n3071);
   U1059 : OAI22_X1 port map( A1 => n14403, A2 => n12495, B1 => n14380, B2 => 
                           n12489, ZN => n3074);
   U1060 : AOI221_X1 port map( B1 => n12507, B2 => n11590, C1 => n12501, C2 => 
                           n11410, A => n3055, ZN => n3052);
   U1061 : OAI22_X1 port map( A1 => n14402, A2 => n12495, B1 => n14379, B2 => 
                           n12489, ZN => n3055);
   U1062 : AOI221_X1 port map( B1 => n12507, B2 => n11591, C1 => n12501, C2 => 
                           n11411, A => n3036, ZN => n3033);
   U1063 : OAI22_X1 port map( A1 => n14401, A2 => n12495, B1 => n14378, B2 => 
                           n12489, ZN => n3036);
   U1064 : AOI221_X1 port map( B1 => n12507, B2 => n11592, C1 => n12501, C2 => 
                           n11412, A => n3017, ZN => n3014);
   U1065 : OAI22_X1 port map( A1 => n14400, A2 => n12495, B1 => n14377, B2 => 
                           n12489, ZN => n3017);
   U1066 : AOI221_X1 port map( B1 => n12507, B2 => n11593, C1 => n12501, C2 => 
                           n11413, A => n2998, ZN => n2995);
   U1067 : OAI22_X1 port map( A1 => n14399, A2 => n12495, B1 => n14376, B2 => 
                           n12489, ZN => n2998);
   U1068 : AOI221_X1 port map( B1 => n12507, B2 => n11594, C1 => n12501, C2 => 
                           n11414, A => n2979, ZN => n2976);
   U1069 : OAI22_X1 port map( A1 => n14398, A2 => n12495, B1 => n14375, B2 => 
                           n12489, ZN => n2979);
   U1070 : AOI221_X1 port map( B1 => n12508, B2 => n11595, C1 => n12502, C2 => 
                           n11415, A => n2960, ZN => n2957);
   U1071 : OAI22_X1 port map( A1 => n14397, A2 => n12496, B1 => n14374, B2 => 
                           n12490, ZN => n2960);
   U1072 : AOI221_X1 port map( B1 => n12508, B2 => n11596, C1 => n12502, C2 => 
                           n11416, A => n2941, ZN => n2938);
   U1073 : OAI22_X1 port map( A1 => n14396, A2 => n12496, B1 => n14373, B2 => 
                           n12490, ZN => n2941);
   U1074 : AOI221_X1 port map( B1 => n12508, B2 => n11597, C1 => n12502, C2 => 
                           n11417, A => n2922, ZN => n2919);
   U1075 : OAI22_X1 port map( A1 => n14395, A2 => n12496, B1 => n14372, B2 => 
                           n12490, ZN => n2922);
   U1076 : AOI221_X1 port map( B1 => n12508, B2 => n11598, C1 => n12502, C2 => 
                           n11418, A => n2903, ZN => n2900);
   U1077 : OAI22_X1 port map( A1 => n14394, A2 => n12496, B1 => n14371, B2 => 
                           n12490, ZN => n2903);
   U1078 : AOI221_X1 port map( B1 => n12508, B2 => n11599, C1 => n12502, C2 => 
                           n11419, A => n2884, ZN => n2881);
   U1079 : OAI22_X1 port map( A1 => n14393, A2 => n12496, B1 => n14370, B2 => 
                           n12490, ZN => n2884);
   U1080 : AOI221_X1 port map( B1 => n12508, B2 => n11600, C1 => n12502, C2 => 
                           n11420, A => n2865, ZN => n2862);
   U1081 : OAI22_X1 port map( A1 => n14392, A2 => n12496, B1 => n14369, B2 => 
                           n12490, ZN => n2865);
   U1082 : AOI221_X1 port map( B1 => n12508, B2 => n11601, C1 => n12502, C2 => 
                           n11421, A => n2846, ZN => n2843);
   U1083 : OAI22_X1 port map( A1 => n14391, A2 => n12496, B1 => n14368, B2 => 
                           n12490, ZN => n2846);
   U1084 : AOI221_X1 port map( B1 => n12508, B2 => n11602, C1 => n12502, C2 => 
                           n11422, A => n2827, ZN => n2824);
   U1085 : OAI22_X1 port map( A1 => n14390, A2 => n12496, B1 => n14367, B2 => 
                           n12490, ZN => n2827);
   U1086 : AOI221_X1 port map( B1 => n12508, B2 => n11603, C1 => n12502, C2 => 
                           n11423, A => n2808, ZN => n2805);
   U1087 : OAI22_X1 port map( A1 => n14389, A2 => n12496, B1 => n14366, B2 => 
                           n12490, ZN => n2808);
   U1088 : AOI221_X1 port map( B1 => n12508, B2 => n11604, C1 => n12502, C2 => 
                           n11424, A => n2789, ZN => n2786);
   U1089 : OAI22_X1 port map( A1 => n14388, A2 => n12496, B1 => n14365, B2 => 
                           n12490, ZN => n2789);
   U1090 : AOI221_X1 port map( B1 => n12508, B2 => n11605, C1 => n12502, C2 => 
                           n11425, A => n2770, ZN => n2767);
   U1091 : OAI22_X1 port map( A1 => n14387, A2 => n12496, B1 => n14364, B2 => 
                           n12490, ZN => n2770);
   U1092 : AOI221_X1 port map( B1 => n12508, B2 => n11606, C1 => n12502, C2 => 
                           n11426, A => n2751, ZN => n2748);
   U1093 : OAI22_X1 port map( A1 => n14386, A2 => n12496, B1 => n14363, B2 => 
                           n12490, ZN => n2751);
   U1094 : AOI221_X1 port map( B1 => n12509, B2 => n11607, C1 => n12503, C2 => 
                           n11427, A => n2732, ZN => n2729);
   U1095 : OAI22_X1 port map( A1 => n14288, A2 => n12497, B1 => n14252, B2 => 
                           n12491, ZN => n2732);
   U1096 : AOI221_X1 port map( B1 => n12509, B2 => n11608, C1 => n12503, C2 => 
                           n11428, A => n2713, ZN => n2710);
   U1097 : OAI22_X1 port map( A1 => n14287, A2 => n12497, B1 => n14251, B2 => 
                           n12491, ZN => n2713);
   U1098 : AOI221_X1 port map( B1 => n12509, B2 => n11609, C1 => n12503, C2 => 
                           n11429, A => n2694, ZN => n2691);
   U1099 : OAI22_X1 port map( A1 => n14286, A2 => n12497, B1 => n14250, B2 => 
                           n12491, ZN => n2694);
   U1100 : AOI221_X1 port map( B1 => n12509, B2 => n11610, C1 => n12503, C2 => 
                           n11430, A => n2675, ZN => n2672);
   U1101 : OAI22_X1 port map( A1 => n14285, A2 => n12497, B1 => n14249, B2 => 
                           n12491, ZN => n2675);
   U1102 : AOI221_X1 port map( B1 => n12509, B2 => n11611, C1 => n12503, C2 => 
                           n11431, A => n2656, ZN => n2653);
   U1103 : OAI22_X1 port map( A1 => n14284, A2 => n12497, B1 => n14248, B2 => 
                           n12491, ZN => n2656);
   U1104 : AOI221_X1 port map( B1 => n12509, B2 => n11612, C1 => n12503, C2 => 
                           n11432, A => n2637, ZN => n2634);
   U1105 : OAI22_X1 port map( A1 => n14283, A2 => n12497, B1 => n14247, B2 => 
                           n12491, ZN => n2637);
   U1106 : AOI221_X1 port map( B1 => n12509, B2 => n11613, C1 => n12503, C2 => 
                           n11433, A => n2618, ZN => n2615);
   U1107 : OAI22_X1 port map( A1 => n14282, A2 => n12497, B1 => n14246, B2 => 
                           n12491, ZN => n2618);
   U1108 : AOI221_X1 port map( B1 => n12509, B2 => n11614, C1 => n12503, C2 => 
                           n11434, A => n2599, ZN => n2596);
   U1109 : OAI22_X1 port map( A1 => n14281, A2 => n12497, B1 => n14245, B2 => 
                           n12491, ZN => n2599);
   U1110 : AOI221_X1 port map( B1 => n12509, B2 => n11615, C1 => n12503, C2 => 
                           n11435, A => n2580, ZN => n2577);
   U1111 : OAI22_X1 port map( A1 => n14280, A2 => n12497, B1 => n14244, B2 => 
                           n12491, ZN => n2580);
   U1112 : AOI221_X1 port map( B1 => n12509, B2 => n11616, C1 => n12503, C2 => 
                           n11436, A => n2561, ZN => n2558);
   U1113 : OAI22_X1 port map( A1 => n14279, A2 => n12497, B1 => n14243, B2 => 
                           n12491, ZN => n2561);
   U1114 : AOI221_X1 port map( B1 => n12509, B2 => n11617, C1 => n12503, C2 => 
                           n11437, A => n2542, ZN => n2539);
   U1115 : OAI22_X1 port map( A1 => n14278, A2 => n12497, B1 => n14242, B2 => 
                           n12491, ZN => n2542);
   U1116 : AOI221_X1 port map( B1 => n12509, B2 => n11618, C1 => n12503, C2 => 
                           n11438, A => n2523, ZN => n2520);
   U1117 : OAI22_X1 port map( A1 => n14277, A2 => n12497, B1 => n14241, B2 => 
                           n12491, ZN => n2523);
   U1118 : AOI221_X1 port map( B1 => n12510, B2 => n11619, C1 => n12504, C2 => 
                           n11439, A => n2504, ZN => n2501);
   U1119 : OAI22_X1 port map( A1 => n14276, A2 => n12498, B1 => n14240, B2 => 
                           n12492, ZN => n2504);
   U1120 : AOI221_X1 port map( B1 => n12510, B2 => n11620, C1 => n12504, C2 => 
                           n11440, A => n2485, ZN => n2482);
   U1121 : OAI22_X1 port map( A1 => n14275, A2 => n12498, B1 => n14239, B2 => 
                           n12492, ZN => n2485);
   U1122 : AOI221_X1 port map( B1 => n12510, B2 => n11621, C1 => n12504, C2 => 
                           n11441, A => n2466, ZN => n2463);
   U1123 : OAI22_X1 port map( A1 => n14274, A2 => n12498, B1 => n14238, B2 => 
                           n12492, ZN => n2466);
   U1124 : AOI221_X1 port map( B1 => n12510, B2 => n11622, C1 => n12504, C2 => 
                           n11442, A => n2447, ZN => n2444);
   U1125 : OAI22_X1 port map( A1 => n14273, A2 => n12498, B1 => n14237, B2 => 
                           n12492, ZN => n2447);
   U1126 : AOI221_X1 port map( B1 => n12510, B2 => n11623, C1 => n12504, C2 => 
                           n11443, A => n2428, ZN => n2425);
   U1127 : OAI22_X1 port map( A1 => n14272, A2 => n12498, B1 => n14236, B2 => 
                           n12492, ZN => n2428);
   U1128 : AOI221_X1 port map( B1 => n12510, B2 => n11624, C1 => n12504, C2 => 
                           n11444, A => n2409, ZN => n2406);
   U1129 : OAI22_X1 port map( A1 => n14271, A2 => n12498, B1 => n14235, B2 => 
                           n12492, ZN => n2409);
   U1130 : AOI221_X1 port map( B1 => n12510, B2 => n11625, C1 => n12504, C2 => 
                           n11445, A => n2390, ZN => n2387);
   U1131 : OAI22_X1 port map( A1 => n14270, A2 => n12498, B1 => n14234, B2 => 
                           n12492, ZN => n2390);
   U1132 : AOI221_X1 port map( B1 => n12510, B2 => n11626, C1 => n12504, C2 => 
                           n11446, A => n2371, ZN => n2368);
   U1133 : OAI22_X1 port map( A1 => n14269, A2 => n12498, B1 => n14233, B2 => 
                           n12492, ZN => n2371);
   U1134 : AOI221_X1 port map( B1 => n12510, B2 => n11627, C1 => n12504, C2 => 
                           n11447, A => n2352, ZN => n2349);
   U1135 : OAI22_X1 port map( A1 => n14268, A2 => n12498, B1 => n14232, B2 => 
                           n12492, ZN => n2352);
   U1136 : AOI221_X1 port map( B1 => n12510, B2 => n11628, C1 => n12504, C2 => 
                           n11448, A => n2333, ZN => n2330);
   U1137 : OAI22_X1 port map( A1 => n14267, A2 => n12498, B1 => n14231, B2 => 
                           n12492, ZN => n2333);
   U1138 : AOI221_X1 port map( B1 => n12510, B2 => n11629, C1 => n12504, C2 => 
                           n11449, A => n2314, ZN => n2311);
   U1139 : OAI22_X1 port map( A1 => n14266, A2 => n12498, B1 => n14230, B2 => 
                           n12492, ZN => n2314);
   U1140 : AOI221_X1 port map( B1 => n12510, B2 => n11630, C1 => n12504, C2 => 
                           n11450, A => n2295, ZN => n2292);
   U1141 : OAI22_X1 port map( A1 => n14265, A2 => n12498, B1 => n14229, B2 => 
                           n12492, ZN => n2295);
   U1142 : AOI221_X1 port map( B1 => n12511, B2 => n11631, C1 => n12505, C2 => 
                           n11451, A => n2276, ZN => n2273);
   U1143 : OAI22_X1 port map( A1 => n14264, A2 => n12499, B1 => n14228, B2 => 
                           n12493, ZN => n2276);
   U1144 : AOI221_X1 port map( B1 => n12511, B2 => n11632, C1 => n12505, C2 => 
                           n11452, A => n2257, ZN => n2254);
   U1145 : OAI22_X1 port map( A1 => n14263, A2 => n12499, B1 => n14227, B2 => 
                           n12493, ZN => n2257);
   U1146 : AOI221_X1 port map( B1 => n12511, B2 => n11633, C1 => n12505, C2 => 
                           n11453, A => n2238, ZN => n2235);
   U1147 : OAI22_X1 port map( A1 => n14262, A2 => n12499, B1 => n14226, B2 => 
                           n12493, ZN => n2238);
   U1148 : AOI221_X1 port map( B1 => n12511, B2 => n11634, C1 => n12505, C2 => 
                           n11454, A => n2219, ZN => n2216);
   U1149 : OAI22_X1 port map( A1 => n14261, A2 => n12499, B1 => n14225, B2 => 
                           n12493, ZN => n2219);
   U1150 : AOI221_X1 port map( B1 => n12511, B2 => n11635, C1 => n12505, C2 => 
                           n11455, A => n2200, ZN => n2197);
   U1151 : OAI22_X1 port map( A1 => n14260, A2 => n12499, B1 => n14224, B2 => 
                           n12493, ZN => n2200);
   U1152 : AOI221_X1 port map( B1 => n12511, B2 => n11636, C1 => n12505, C2 => 
                           n11456, A => n2181, ZN => n2178);
   U1153 : OAI22_X1 port map( A1 => n14259, A2 => n12499, B1 => n14223, B2 => 
                           n12493, ZN => n2181);
   U1154 : AOI221_X1 port map( B1 => n12511, B2 => n11637, C1 => n12505, C2 => 
                           n11457, A => n2162, ZN => n2159);
   U1155 : OAI22_X1 port map( A1 => n14258, A2 => n12499, B1 => n14222, B2 => 
                           n12493, ZN => n2162);
   U1156 : AOI221_X1 port map( B1 => n12511, B2 => n11638, C1 => n12505, C2 => 
                           n11458, A => n2143, ZN => n2140);
   U1157 : OAI22_X1 port map( A1 => n14257, A2 => n12499, B1 => n14221, B2 => 
                           n12493, ZN => n2143);
   U1158 : AOI221_X1 port map( B1 => n12511, B2 => n11639, C1 => n12505, C2 => 
                           n11459, A => n2124, ZN => n2121);
   U1159 : OAI22_X1 port map( A1 => n14256, A2 => n12499, B1 => n14220, B2 => 
                           n12493, ZN => n2124);
   U1160 : AOI221_X1 port map( B1 => n12511, B2 => n11640, C1 => n12505, C2 => 
                           n11460, A => n2105, ZN => n2102);
   U1161 : OAI22_X1 port map( A1 => n14255, A2 => n12499, B1 => n14219, B2 => 
                           n12493, ZN => n2105);
   U1162 : AOI221_X1 port map( B1 => n12511, B2 => n11641, C1 => n12505, C2 => 
                           n11461, A => n2086, ZN => n2083);
   U1163 : OAI22_X1 port map( A1 => n14254, A2 => n12499, B1 => n14218, B2 => 
                           n12493, ZN => n2086);
   U1164 : AOI221_X1 port map( B1 => n12511, B2 => n11765, C1 => n12505, C2 => 
                           n11585, A => n2067, ZN => n2064);
   U1165 : OAI22_X1 port map( A1 => n14253, A2 => n12499, B1 => n14217, B2 => 
                           n12493, ZN => n2067);
   U1166 : AOI221_X1 port map( B1 => n12512, B2 => n13835, C1 => n12506, C2 => 
                           n13839, A => n2048, ZN => n2045);
   U1167 : OAI22_X1 port map( A1 => n13847, A2 => n12500, B1 => n13843, B2 => 
                           n12494, ZN => n2048);
   U1168 : AOI221_X1 port map( B1 => n12512, B2 => n13834, C1 => n12506, C2 => 
                           n13838, A => n2029, ZN => n2026);
   U1169 : OAI22_X1 port map( A1 => n13846, A2 => n12500, B1 => n13842, B2 => 
                           n12494, ZN => n2029);
   U1170 : AOI221_X1 port map( B1 => n12512, B2 => n13833, C1 => n12506, C2 => 
                           n13837, A => n2010, ZN => n2007);
   U1171 : OAI22_X1 port map( A1 => n13845, A2 => n12500, B1 => n13841, B2 => 
                           n12494, ZN => n2010);
   U1172 : AOI221_X1 port map( B1 => n12512, B2 => n13832, C1 => n12506, C2 => 
                           n13836, A => n1965, ZN => n1956);
   U1173 : OAI22_X1 port map( A1 => n13844, A2 => n12500, B1 => n13840, B2 => 
                           n12494, ZN => n1965);
   U1174 : AOI221_X1 port map( B1 => n12387, B2 => n14153, C1 => n12381, C2 => 
                           n14154, A => n3207, ZN => n3200);
   U1175 : OAI22_X1 port map( A1 => n13746, A2 => n12375, B1 => n13730, B2 => 
                           n12369, ZN => n3207);
   U1176 : AOI221_X1 port map( B1 => n12483, B2 => n11642, C1 => n12477, C2 => 
                           n11462, A => n3195, ZN => n3184);
   U1177 : OAI22_X1 port map( A1 => n13539, A2 => n12471, B1 => n13494, B2 => 
                           n12465, ZN => n3195);
   U1178 : AOI221_X1 port map( B1 => n12387, B2 => n14082, C1 => n12381, C2 => 
                           n14129, A => n3178, ZN => n3173);
   U1179 : OAI22_X1 port map( A1 => n13745, A2 => n12375, B1 => n13729, B2 => 
                           n12369, ZN => n3178);
   U1180 : AOI221_X1 port map( B1 => n12483, B2 => n11643, C1 => n12477, C2 => 
                           n11463, A => n3170, ZN => n3165);
   U1181 : OAI22_X1 port map( A1 => n13538, A2 => n12471, B1 => n13493, B2 => 
                           n12465, ZN => n3170);
   U1182 : AOI221_X1 port map( B1 => n12387, B2 => n14081, C1 => n12381, C2 => 
                           n14128, A => n3159, ZN => n3154);
   U1183 : OAI22_X1 port map( A1 => n13744, A2 => n12375, B1 => n13728, B2 => 
                           n12369, ZN => n3159);
   U1184 : AOI221_X1 port map( B1 => n12483, B2 => n11644, C1 => n12477, C2 => 
                           n11464, A => n3151, ZN => n3146);
   U1185 : OAI22_X1 port map( A1 => n13537, A2 => n12471, B1 => n13492, B2 => 
                           n12465, ZN => n3151);
   U1186 : AOI221_X1 port map( B1 => n12483, B2 => n11645, C1 => n12477, C2 => 
                           n11465, A => n3132, ZN => n3127);
   U1187 : OAI22_X1 port map( A1 => n13536, A2 => n12471, B1 => n13491, B2 => 
                           n12465, ZN => n3132);
   U1188 : AOI221_X1 port map( B1 => n12483, B2 => n11646, C1 => n12477, C2 => 
                           n11466, A => n3113, ZN => n3108);
   U1189 : OAI22_X1 port map( A1 => n14360, A2 => n12471, B1 => n13490, B2 => 
                           n12465, ZN => n3113);
   U1190 : AOI221_X1 port map( B1 => n12387, B2 => n14078, C1 => n12381, C2 => 
                           n14125, A => n3102, ZN => n3097);
   U1191 : OAI22_X1 port map( A1 => n13891, A2 => n12375, B1 => n13725, B2 => 
                           n12369, ZN => n3102);
   U1192 : AOI221_X1 port map( B1 => n12483, B2 => n11647, C1 => n12477, C2 => 
                           n11467, A => n3094, ZN => n3089);
   U1193 : OAI22_X1 port map( A1 => n14359, A2 => n12471, B1 => n13489, B2 => 
                           n12465, ZN => n3094);
   U1194 : AOI221_X1 port map( B1 => n12387, B2 => n14077, C1 => n12381, C2 => 
                           n14124, A => n3083, ZN => n3078);
   U1195 : OAI22_X1 port map( A1 => n13890, A2 => n12375, B1 => n13724, B2 => 
                           n12369, ZN => n3083);
   U1196 : AOI221_X1 port map( B1 => n12483, B2 => n11648, C1 => n12477, C2 => 
                           n11468, A => n3075, ZN => n3070);
   U1197 : OAI22_X1 port map( A1 => n14358, A2 => n12471, B1 => n13488, B2 => 
                           n12465, ZN => n3075);
   U1198 : AOI221_X1 port map( B1 => n12483, B2 => n11649, C1 => n12477, C2 => 
                           n11469, A => n3056, ZN => n3051);
   U1199 : OAI22_X1 port map( A1 => n14340, A2 => n12471, B1 => n13487, B2 => 
                           n12465, ZN => n3056);
   U1200 : AOI221_X1 port map( B1 => n12483, B2 => n11650, C1 => n12477, C2 => 
                           n11470, A => n3037, ZN => n3032);
   U1201 : OAI22_X1 port map( A1 => n14339, A2 => n12471, B1 => n13486, B2 => 
                           n12465, ZN => n3037);
   U1202 : AOI221_X1 port map( B1 => n12483, B2 => n11651, C1 => n12477, C2 => 
                           n11471, A => n3018, ZN => n3013);
   U1203 : OAI22_X1 port map( A1 => n14338, A2 => n12471, B1 => n13485, B2 => 
                           n12465, ZN => n3018);
   U1204 : AOI221_X1 port map( B1 => n12483, B2 => n11652, C1 => n12477, C2 => 
                           n11472, A => n2999, ZN => n2994);
   U1205 : OAI22_X1 port map( A1 => n14337, A2 => n12471, B1 => n13484, B2 => 
                           n12465, ZN => n2999);
   U1206 : AOI221_X1 port map( B1 => n12483, B2 => n11653, C1 => n12477, C2 => 
                           n11473, A => n2980, ZN => n2975);
   U1207 : OAI22_X1 port map( A1 => n14336, A2 => n12471, B1 => n13483, B2 => 
                           n12465, ZN => n2980);
   U1208 : AOI221_X1 port map( B1 => n12484, B2 => n11654, C1 => n12478, C2 => 
                           n11474, A => n2961, ZN => n2956);
   U1209 : OAI22_X1 port map( A1 => n14335, A2 => n12472, B1 => n13482, B2 => 
                           n12466, ZN => n2961);
   U1210 : AOI221_X1 port map( B1 => n12484, B2 => n11655, C1 => n12478, C2 => 
                           n11475, A => n2942, ZN => n2937);
   U1211 : OAI22_X1 port map( A1 => n14334, A2 => n12472, B1 => n13481, B2 => 
                           n12466, ZN => n2942);
   U1212 : AOI221_X1 port map( B1 => n12484, B2 => n11656, C1 => n12478, C2 => 
                           n11476, A => n2923, ZN => n2918);
   U1213 : OAI22_X1 port map( A1 => n14333, A2 => n12472, B1 => n13480, B2 => 
                           n12466, ZN => n2923);
   U1214 : AOI221_X1 port map( B1 => n12484, B2 => n11657, C1 => n12478, C2 => 
                           n11477, A => n2904, ZN => n2899);
   U1215 : OAI22_X1 port map( A1 => n14332, A2 => n12472, B1 => n13479, B2 => 
                           n12466, ZN => n2904);
   U1216 : AOI221_X1 port map( B1 => n12484, B2 => n11658, C1 => n12478, C2 => 
                           n11478, A => n2885, ZN => n2880);
   U1217 : OAI22_X1 port map( A1 => n13535, A2 => n12472, B1 => n13478, B2 => 
                           n12466, ZN => n2885);
   U1218 : AOI221_X1 port map( B1 => n12484, B2 => n11659, C1 => n12478, C2 => 
                           n11479, A => n2866, ZN => n2861);
   U1219 : OAI22_X1 port map( A1 => n14331, A2 => n12472, B1 => n13477, B2 => 
                           n12466, ZN => n2866);
   U1220 : AOI221_X1 port map( B1 => n12484, B2 => n11660, C1 => n12478, C2 => 
                           n11480, A => n2847, ZN => n2842);
   U1221 : OAI22_X1 port map( A1 => n14330, A2 => n12472, B1 => n13476, B2 => 
                           n12466, ZN => n2847);
   U1222 : AOI221_X1 port map( B1 => n12484, B2 => n11661, C1 => n12478, C2 => 
                           n11481, A => n2828, ZN => n2823);
   U1223 : OAI22_X1 port map( A1 => n14329, A2 => n12472, B1 => n13475, B2 => 
                           n12466, ZN => n2828);
   U1224 : AOI221_X1 port map( B1 => n12484, B2 => n11662, C1 => n12478, C2 => 
                           n11482, A => n2809, ZN => n2804);
   U1225 : OAI22_X1 port map( A1 => n13534, A2 => n12472, B1 => n13474, B2 => 
                           n12466, ZN => n2809);
   U1226 : AOI221_X1 port map( B1 => n12484, B2 => n11663, C1 => n12478, C2 => 
                           n11483, A => n2790, ZN => n2785);
   U1227 : OAI22_X1 port map( A1 => n13533, A2 => n12472, B1 => n13473, B2 => 
                           n12466, ZN => n2790);
   U1228 : AOI221_X1 port map( B1 => n12484, B2 => n11664, C1 => n12478, C2 => 
                           n11484, A => n2771, ZN => n2766);
   U1229 : OAI22_X1 port map( A1 => n13532, A2 => n12472, B1 => n13472, B2 => 
                           n12466, ZN => n2771);
   U1230 : AOI221_X1 port map( B1 => n12484, B2 => n11665, C1 => n12478, C2 => 
                           n11485, A => n2752, ZN => n2747);
   U1231 : OAI22_X1 port map( A1 => n13531, A2 => n12472, B1 => n13471, B2 => 
                           n12466, ZN => n2752);
   U1232 : AOI221_X1 port map( B1 => n12485, B2 => n11666, C1 => n12479, C2 => 
                           n11486, A => n2733, ZN => n2728);
   U1233 : OAI22_X1 port map( A1 => n13530, A2 => n12473, B1 => n13470, B2 => 
                           n12467, ZN => n2733);
   U1234 : AOI221_X1 port map( B1 => n12485, B2 => n11667, C1 => n12479, C2 => 
                           n11487, A => n2714, ZN => n2709);
   U1235 : OAI22_X1 port map( A1 => n13529, A2 => n12473, B1 => n13469, B2 => 
                           n12467, ZN => n2714);
   U1236 : AOI221_X1 port map( B1 => n12485, B2 => n11668, C1 => n12479, C2 => 
                           n11488, A => n2695, ZN => n2690);
   U1237 : OAI22_X1 port map( A1 => n13528, A2 => n12473, B1 => n13468, B2 => 
                           n12467, ZN => n2695);
   U1238 : AOI221_X1 port map( B1 => n12485, B2 => n11669, C1 => n12479, C2 => 
                           n11489, A => n2676, ZN => n2671);
   U1239 : OAI22_X1 port map( A1 => n13527, A2 => n12473, B1 => n13467, B2 => 
                           n12467, ZN => n2676);
   U1240 : AOI221_X1 port map( B1 => n12485, B2 => n11670, C1 => n12479, C2 => 
                           n11490, A => n2657, ZN => n2652);
   U1241 : OAI22_X1 port map( A1 => n13526, A2 => n12473, B1 => n13466, B2 => 
                           n12467, ZN => n2657);
   U1242 : AOI221_X1 port map( B1 => n12485, B2 => n11671, C1 => n12479, C2 => 
                           n11491, A => n2638, ZN => n2633);
   U1243 : OAI22_X1 port map( A1 => n13525, A2 => n12473, B1 => n13465, B2 => 
                           n12467, ZN => n2638);
   U1244 : AOI221_X1 port map( B1 => n12485, B2 => n11672, C1 => n12479, C2 => 
                           n11492, A => n2619, ZN => n2614);
   U1245 : OAI22_X1 port map( A1 => n13524, A2 => n12473, B1 => n13464, B2 => 
                           n12467, ZN => n2619);
   U1246 : AOI221_X1 port map( B1 => n12485, B2 => n11673, C1 => n12479, C2 => 
                           n11493, A => n2600, ZN => n2595);
   U1247 : OAI22_X1 port map( A1 => n13523, A2 => n12473, B1 => n13463, B2 => 
                           n12467, ZN => n2600);
   U1248 : AOI221_X1 port map( B1 => n12485, B2 => n11674, C1 => n12479, C2 => 
                           n11494, A => n2581, ZN => n2576);
   U1249 : OAI22_X1 port map( A1 => n13522, A2 => n12473, B1 => n13462, B2 => 
                           n12467, ZN => n2581);
   U1250 : AOI221_X1 port map( B1 => n12485, B2 => n11675, C1 => n12479, C2 => 
                           n11495, A => n2562, ZN => n2557);
   U1251 : OAI22_X1 port map( A1 => n13521, A2 => n12473, B1 => n13461, B2 => 
                           n12467, ZN => n2562);
   U1252 : AOI221_X1 port map( B1 => n12485, B2 => n11676, C1 => n12479, C2 => 
                           n11496, A => n2543, ZN => n2538);
   U1253 : OAI22_X1 port map( A1 => n13520, A2 => n12473, B1 => n13460, B2 => 
                           n12467, ZN => n2543);
   U1254 : AOI221_X1 port map( B1 => n12485, B2 => n11677, C1 => n12479, C2 => 
                           n11497, A => n2524, ZN => n2519);
   U1255 : OAI22_X1 port map( A1 => n13519, A2 => n12473, B1 => n13459, B2 => 
                           n12467, ZN => n2524);
   U1256 : AOI221_X1 port map( B1 => n12486, B2 => n11678, C1 => n12480, C2 => 
                           n11498, A => n2505, ZN => n2500);
   U1257 : OAI22_X1 port map( A1 => n13518, A2 => n12474, B1 => n13458, B2 => 
                           n12468, ZN => n2505);
   U1258 : AOI221_X1 port map( B1 => n12486, B2 => n11679, C1 => n12480, C2 => 
                           n11499, A => n2486, ZN => n2481);
   U1259 : OAI22_X1 port map( A1 => n13517, A2 => n12474, B1 => n13457, B2 => 
                           n12468, ZN => n2486);
   U1260 : AOI221_X1 port map( B1 => n12486, B2 => n11680, C1 => n12480, C2 => 
                           n11500, A => n2467, ZN => n2462);
   U1261 : OAI22_X1 port map( A1 => n13516, A2 => n12474, B1 => n13456, B2 => 
                           n12468, ZN => n2467);
   U1262 : AOI221_X1 port map( B1 => n12486, B2 => n11681, C1 => n12480, C2 => 
                           n11501, A => n2448, ZN => n2443);
   U1263 : OAI22_X1 port map( A1 => n14460, A2 => n12474, B1 => n13455, B2 => 
                           n12468, ZN => n2448);
   U1264 : AOI221_X1 port map( B1 => n12486, B2 => n11682, C1 => n12480, C2 => 
                           n11502, A => n2429, ZN => n2424);
   U1265 : OAI22_X1 port map( A1 => n14459, A2 => n12474, B1 => n13454, B2 => 
                           n12468, ZN => n2429);
   U1266 : AOI221_X1 port map( B1 => n12486, B2 => n11683, C1 => n12480, C2 => 
                           n11503, A => n2410, ZN => n2405);
   U1267 : OAI22_X1 port map( A1 => n14458, A2 => n12474, B1 => n13453, B2 => 
                           n12468, ZN => n2410);
   U1268 : AOI221_X1 port map( B1 => n12486, B2 => n11684, C1 => n12480, C2 => 
                           n11504, A => n2391, ZN => n2386);
   U1269 : OAI22_X1 port map( A1 => n14457, A2 => n12474, B1 => n13452, B2 => 
                           n12468, ZN => n2391);
   U1270 : AOI221_X1 port map( B1 => n12486, B2 => n11685, C1 => n12480, C2 => 
                           n11505, A => n2372, ZN => n2367);
   U1271 : OAI22_X1 port map( A1 => n13515, A2 => n12474, B1 => n13451, B2 => 
                           n12468, ZN => n2372);
   U1272 : AOI221_X1 port map( B1 => n12486, B2 => n11686, C1 => n12480, C2 => 
                           n11506, A => n2353, ZN => n2348);
   U1273 : OAI22_X1 port map( A1 => n13514, A2 => n12474, B1 => n13450, B2 => 
                           n12468, ZN => n2353);
   U1274 : AOI221_X1 port map( B1 => n12486, B2 => n11687, C1 => n12480, C2 => 
                           n11507, A => n2334, ZN => n2329);
   U1275 : OAI22_X1 port map( A1 => n13513, A2 => n12474, B1 => n13449, B2 => 
                           n12468, ZN => n2334);
   U1276 : AOI221_X1 port map( B1 => n12486, B2 => n11688, C1 => n12480, C2 => 
                           n11508, A => n2315, ZN => n2310);
   U1277 : OAI22_X1 port map( A1 => n13512, A2 => n12474, B1 => n13448, B2 => 
                           n12468, ZN => n2315);
   U1278 : AOI221_X1 port map( B1 => n12486, B2 => n11689, C1 => n12480, C2 => 
                           n11509, A => n2296, ZN => n2291);
   U1279 : OAI22_X1 port map( A1 => n13511, A2 => n12474, B1 => n13447, B2 => 
                           n12468, ZN => n2296);
   U1280 : AOI221_X1 port map( B1 => n12487, B2 => n11690, C1 => n12481, C2 => 
                           n11510, A => n2277, ZN => n2272);
   U1281 : OAI22_X1 port map( A1 => n13510, A2 => n12475, B1 => n13446, B2 => 
                           n12469, ZN => n2277);
   U1282 : AOI221_X1 port map( B1 => n12487, B2 => n11691, C1 => n12481, C2 => 
                           n11511, A => n2258, ZN => n2253);
   U1283 : OAI22_X1 port map( A1 => n13509, A2 => n12475, B1 => n13445, B2 => 
                           n12469, ZN => n2258);
   U1284 : AOI221_X1 port map( B1 => n12487, B2 => n11692, C1 => n12481, C2 => 
                           n11512, A => n2239, ZN => n2234);
   U1285 : OAI22_X1 port map( A1 => n13508, A2 => n12475, B1 => n13444, B2 => 
                           n12469, ZN => n2239);
   U1286 : AOI221_X1 port map( B1 => n12487, B2 => n11693, C1 => n12481, C2 => 
                           n11513, A => n2220, ZN => n2215);
   U1287 : OAI22_X1 port map( A1 => n13507, A2 => n12475, B1 => n13443, B2 => 
                           n12469, ZN => n2220);
   U1288 : AOI221_X1 port map( B1 => n12487, B2 => n11694, C1 => n12481, C2 => 
                           n11514, A => n2201, ZN => n2196);
   U1289 : OAI22_X1 port map( A1 => n13506, A2 => n12475, B1 => n13442, B2 => 
                           n12469, ZN => n2201);
   U1290 : AOI221_X1 port map( B1 => n12487, B2 => n11695, C1 => n12481, C2 => 
                           n11515, A => n2182, ZN => n2177);
   U1291 : OAI22_X1 port map( A1 => n13505, A2 => n12475, B1 => n13441, B2 => 
                           n12469, ZN => n2182);
   U1292 : AOI221_X1 port map( B1 => n12487, B2 => n11696, C1 => n12481, C2 => 
                           n11516, A => n2163, ZN => n2158);
   U1293 : OAI22_X1 port map( A1 => n13504, A2 => n12475, B1 => n13440, B2 => 
                           n12469, ZN => n2163);
   U1294 : AOI221_X1 port map( B1 => n12487, B2 => n11697, C1 => n12481, C2 => 
                           n11517, A => n2144, ZN => n2139);
   U1295 : OAI22_X1 port map( A1 => n13503, A2 => n12475, B1 => n13439, B2 => 
                           n12469, ZN => n2144);
   U1296 : AOI221_X1 port map( B1 => n12487, B2 => n11698, C1 => n12481, C2 => 
                           n11518, A => n2125, ZN => n2120);
   U1297 : OAI22_X1 port map( A1 => n13502, A2 => n12475, B1 => n13438, B2 => 
                           n12469, ZN => n2125);
   U1298 : AOI221_X1 port map( B1 => n12487, B2 => n11699, C1 => n12481, C2 => 
                           n11519, A => n2106, ZN => n2101);
   U1299 : OAI22_X1 port map( A1 => n13501, A2 => n12475, B1 => n13437, B2 => 
                           n12469, ZN => n2106);
   U1300 : AOI221_X1 port map( B1 => n12487, B2 => n11700, C1 => n12481, C2 => 
                           n11520, A => n2087, ZN => n2082);
   U1301 : OAI22_X1 port map( A1 => n13500, A2 => n12475, B1 => n13436, B2 => 
                           n12469, ZN => n2087);
   U1302 : AOI221_X1 port map( B1 => n12391, B2 => n13893, C1 => n12385, C2 => 
                           n13953, A => n2076, ZN => n2071);
   U1303 : OAI22_X1 port map( A1 => n13735, A2 => n12379, B1 => n13671, B2 => 
                           n12373, ZN => n2076);
   U1304 : AOI221_X1 port map( B1 => n12487, B2 => n11701, C1 => n12481, C2 => 
                           n11521, A => n2068, ZN => n2063);
   U1305 : OAI22_X1 port map( A1 => n13499, A2 => n12475, B1 => n13435, B2 => 
                           n12469, ZN => n2068);
   U1306 : AOI221_X1 port map( B1 => n12392, B2 => n13819, C1 => n12386, C2 => 
                           n13823, A => n2057, ZN => n2052);
   U1307 : OAI22_X1 port map( A1 => n13734, A2 => n12380, B1 => n13670, B2 => 
                           n12374, ZN => n2057);
   U1308 : AOI221_X1 port map( B1 => n12488, B2 => n13860, C1 => n12482, C2 => 
                           n13856, A => n2049, ZN => n2044);
   U1309 : OAI22_X1 port map( A1 => n13498, A2 => n12476, B1 => n13434, B2 => 
                           n12470, ZN => n2049);
   U1310 : AOI221_X1 port map( B1 => n12392, B2 => n13818, C1 => n12386, C2 => 
                           n13822, A => n2038, ZN => n2033);
   U1311 : OAI22_X1 port map( A1 => n13733, A2 => n12380, B1 => n13669, B2 => 
                           n12374, ZN => n2038);
   U1312 : AOI221_X1 port map( B1 => n12488, B2 => n13859, C1 => n12482, C2 => 
                           n13855, A => n2030, ZN => n2025);
   U1313 : OAI22_X1 port map( A1 => n13497, A2 => n12476, B1 => n13433, B2 => 
                           n12470, ZN => n2030);
   U1314 : AOI221_X1 port map( B1 => n12392, B2 => n13817, C1 => n12386, C2 => 
                           n13821, A => n2019, ZN => n2014);
   U1315 : OAI22_X1 port map( A1 => n13732, A2 => n12380, B1 => n13668, B2 => 
                           n12374, ZN => n2019);
   U1316 : AOI221_X1 port map( B1 => n12488, B2 => n13858, C1 => n12482, C2 => 
                           n13854, A => n2011, ZN => n2006);
   U1317 : OAI22_X1 port map( A1 => n13496, A2 => n12476, B1 => n13432, B2 => 
                           n12470, ZN => n2011);
   U1318 : AOI221_X1 port map( B1 => n12392, B2 => n13816, C1 => n12386, C2 => 
                           n13820, A => n1994, ZN => n1979);
   U1319 : OAI22_X1 port map( A1 => n13731, A2 => n12380, B1 => n13667, B2 => 
                           n12374, ZN => n1994);
   U1320 : AOI221_X1 port map( B1 => n12488, B2 => n13857, C1 => n12482, C2 => 
                           n13853, A => n1970, ZN => n1955);
   U1321 : OAI22_X1 port map( A1 => n13495, A2 => n12476, B1 => n13431, B2 => 
                           n12470, ZN => n1970);
   U1322 : AOI221_X1 port map( B1 => n12363, B2 => n14155, C1 => n12357, C2 => 
                           n13831, A => n3210, ZN => n3199);
   U1323 : OAI22_X1 port map( A1 => n13815, A2 => n12351, B1 => n13810, B2 => 
                           n12345, ZN => n3210);
   U1324 : AOI221_X1 port map( B1 => n12459, B2 => n11702, C1 => n12453, C2 => 
                           n11522, A => n3198, ZN => n3183);
   U1325 : OAI22_X1 port map( A1 => n13650, A2 => n12447, B1 => n13603, B2 => 
                           n12441, ZN => n3198);
   U1326 : AOI221_X1 port map( B1 => n12363, B2 => n14152, C1 => n12357, C2 => 
                           n13830, A => n3179, ZN => n3172);
   U1327 : OAI22_X1 port map( A1 => n13814, A2 => n12351, B1 => n13809, B2 => 
                           n12345, ZN => n3179);
   U1328 : AOI221_X1 port map( B1 => n12459, B2 => n11703, C1 => n12453, C2 => 
                           n11523, A => n3171, ZN => n3164);
   U1329 : OAI22_X1 port map( A1 => n13649, A2 => n12447, B1 => n13602, B2 => 
                           n12441, ZN => n3171);
   U1330 : AOI221_X1 port map( B1 => n12363, B2 => n14151, C1 => n12357, C2 => 
                           n13829, A => n3160, ZN => n3153);
   U1331 : OAI22_X1 port map( A1 => n13813, A2 => n12351, B1 => n13808, B2 => 
                           n12345, ZN => n3160);
   U1332 : AOI221_X1 port map( B1 => n12459, B2 => n11704, C1 => n12453, C2 => 
                           n11524, A => n3152, ZN => n3145);
   U1333 : OAI22_X1 port map( A1 => n13648, A2 => n12447, B1 => n13601, B2 => 
                           n12441, ZN => n3152);
   U1334 : AOI221_X1 port map( B1 => n12363, B2 => n14149, C1 => n12357, C2 => 
                           n13828, A => n3141, ZN => n3134);
   U1335 : OAI22_X1 port map( A1 => n13812, A2 => n12351, B1 => n13807, B2 => 
                           n12345, ZN => n3141);
   U1336 : AOI221_X1 port map( B1 => n12459, B2 => n11705, C1 => n12453, C2 => 
                           n11525, A => n3133, ZN => n3126);
   U1337 : OAI22_X1 port map( A1 => n13647, A2 => n12447, B1 => n13600, B2 => 
                           n12441, ZN => n3133);
   U1338 : AOI221_X1 port map( B1 => n12363, B2 => n14150, C1 => n12357, C2 => 
                           n14215, A => n3122, ZN => n3115);
   U1339 : OAI22_X1 port map( A1 => n13811, A2 => n12351, B1 => n13806, B2 => 
                           n12345, ZN => n3122);
   U1340 : AOI221_X1 port map( B1 => n12459, B2 => n11706, C1 => n12453, C2 => 
                           n11526, A => n3114, ZN => n3107);
   U1341 : OAI22_X1 port map( A1 => n14357, A2 => n12447, B1 => n13599, B2 => 
                           n12441, ZN => n3114);
   U1342 : AOI221_X1 port map( B1 => n12363, B2 => n14148, C1 => n12357, C2 => 
                           n14214, A => n3103, ZN => n3096);
   U1343 : OAI22_X1 port map( A1 => n14035, A2 => n12351, B1 => n13805, B2 => 
                           n12345, ZN => n3103);
   U1344 : AOI221_X1 port map( B1 => n12459, B2 => n11707, C1 => n12453, C2 => 
                           n11527, A => n3095, ZN => n3088);
   U1345 : OAI22_X1 port map( A1 => n14356, A2 => n12447, B1 => n13598, B2 => 
                           n12441, ZN => n3095);
   U1346 : AOI221_X1 port map( B1 => n12363, B2 => n14147, C1 => n12357, C2 => 
                           n14213, A => n3084, ZN => n3077);
   U1347 : OAI22_X1 port map( A1 => n14034, A2 => n12351, B1 => n13804, B2 => 
                           n12345, ZN => n3084);
   U1348 : AOI221_X1 port map( B1 => n12459, B2 => n11708, C1 => n12453, C2 => 
                           n11528, A => n3076, ZN => n3069);
   U1349 : OAI22_X1 port map( A1 => n14355, A2 => n12447, B1 => n13597, B2 => 
                           n12441, ZN => n3076);
   U1350 : AOI221_X1 port map( B1 => n12363, B2 => n14146, C1 => n12357, C2 => 
                           n14212, A => n3065, ZN => n3058);
   U1351 : OAI22_X1 port map( A1 => n14033, A2 => n12351, B1 => n13803, B2 => 
                           n12345, ZN => n3065);
   U1352 : AOI221_X1 port map( B1 => n12459, B2 => n11709, C1 => n12453, C2 => 
                           n11529, A => n3057, ZN => n3050);
   U1353 : OAI22_X1 port map( A1 => n14354, A2 => n12447, B1 => n13596, B2 => 
                           n12441, ZN => n3057);
   U1354 : AOI221_X1 port map( B1 => n12363, B2 => n14145, C1 => n12357, C2 => 
                           n14211, A => n3046, ZN => n3039);
   U1355 : OAI22_X1 port map( A1 => n14032, A2 => n12351, B1 => n13802, B2 => 
                           n12345, ZN => n3046);
   U1356 : AOI221_X1 port map( B1 => n12459, B2 => n11710, C1 => n12453, C2 => 
                           n11530, A => n3038, ZN => n3031);
   U1357 : OAI22_X1 port map( A1 => n14353, A2 => n12447, B1 => n13595, B2 => 
                           n12441, ZN => n3038);
   U1358 : AOI221_X1 port map( B1 => n12363, B2 => n14144, C1 => n12357, C2 => 
                           n14210, A => n3027, ZN => n3020);
   U1359 : OAI22_X1 port map( A1 => n14031, A2 => n12351, B1 => n13801, B2 => 
                           n12345, ZN => n3027);
   U1360 : AOI221_X1 port map( B1 => n12459, B2 => n11711, C1 => n12453, C2 => 
                           n11531, A => n3019, ZN => n3012);
   U1361 : OAI22_X1 port map( A1 => n14352, A2 => n12447, B1 => n13594, B2 => 
                           n12441, ZN => n3019);
   U1362 : AOI221_X1 port map( B1 => n12363, B2 => n14143, C1 => n12357, C2 => 
                           n14209, A => n3008, ZN => n3001);
   U1363 : OAI22_X1 port map( A1 => n14030, A2 => n12351, B1 => n13800, B2 => 
                           n12345, ZN => n3008);
   U1364 : AOI221_X1 port map( B1 => n12459, B2 => n11712, C1 => n12453, C2 => 
                           n11532, A => n3000, ZN => n2993);
   U1365 : OAI22_X1 port map( A1 => n14351, A2 => n12447, B1 => n13593, B2 => 
                           n12441, ZN => n3000);
   U1366 : AOI221_X1 port map( B1 => n12363, B2 => n14142, C1 => n12357, C2 => 
                           n14208, A => n2989, ZN => n2982);
   U1367 : OAI22_X1 port map( A1 => n14029, A2 => n12351, B1 => n13799, B2 => 
                           n12345, ZN => n2989);
   U1368 : AOI221_X1 port map( B1 => n12459, B2 => n11713, C1 => n12453, C2 => 
                           n11533, A => n2981, ZN => n2974);
   U1369 : OAI22_X1 port map( A1 => n14350, A2 => n12447, B1 => n13592, B2 => 
                           n12441, ZN => n2981);
   U1370 : AOI221_X1 port map( B1 => n12364, B2 => n14141, C1 => n12358, C2 => 
                           n14207, A => n2970, ZN => n2963);
   U1371 : OAI22_X1 port map( A1 => n14028, A2 => n12352, B1 => n13798, B2 => 
                           n12346, ZN => n2970);
   U1372 : AOI221_X1 port map( B1 => n12460, B2 => n11714, C1 => n12454, C2 => 
                           n11534, A => n2962, ZN => n2955);
   U1373 : OAI22_X1 port map( A1 => n14349, A2 => n12448, B1 => n13591, B2 => 
                           n12442, ZN => n2962);
   U1374 : AOI221_X1 port map( B1 => n12364, B2 => n14140, C1 => n12358, C2 => 
                           n14206, A => n2951, ZN => n2944);
   U1375 : OAI22_X1 port map( A1 => n14027, A2 => n12352, B1 => n13797, B2 => 
                           n12346, ZN => n2951);
   U1376 : AOI221_X1 port map( B1 => n12460, B2 => n11715, C1 => n12454, C2 => 
                           n11535, A => n2943, ZN => n2936);
   U1377 : OAI22_X1 port map( A1 => n14348, A2 => n12448, B1 => n13590, B2 => 
                           n12442, ZN => n2943);
   U1378 : AOI221_X1 port map( B1 => n12364, B2 => n14139, C1 => n12358, C2 => 
                           n14205, A => n2932, ZN => n2925);
   U1379 : OAI22_X1 port map( A1 => n14026, A2 => n12352, B1 => n13796, B2 => 
                           n12346, ZN => n2932);
   U1380 : AOI221_X1 port map( B1 => n12460, B2 => n11716, C1 => n12454, C2 => 
                           n11536, A => n2924, ZN => n2917);
   U1381 : OAI22_X1 port map( A1 => n14347, A2 => n12448, B1 => n13589, B2 => 
                           n12442, ZN => n2924);
   U1382 : AOI221_X1 port map( B1 => n12364, B2 => n14138, C1 => n12358, C2 => 
                           n14204, A => n2913, ZN => n2906);
   U1383 : OAI22_X1 port map( A1 => n14025, A2 => n12352, B1 => n13795, B2 => 
                           n12346, ZN => n2913);
   U1384 : AOI221_X1 port map( B1 => n12460, B2 => n11717, C1 => n12454, C2 => 
                           n11537, A => n2905, ZN => n2898);
   U1385 : OAI22_X1 port map( A1 => n14346, A2 => n12448, B1 => n13588, B2 => 
                           n12442, ZN => n2905);
   U1386 : AOI221_X1 port map( B1 => n12364, B2 => n14137, C1 => n12358, C2 => 
                           n14203, A => n2894, ZN => n2887);
   U1387 : OAI22_X1 port map( A1 => n13952, A2 => n12352, B1 => n13794, B2 => 
                           n12346, ZN => n2894);
   U1388 : AOI221_X1 port map( B1 => n12460, B2 => n11718, C1 => n12454, C2 => 
                           n11538, A => n2886, ZN => n2879);
   U1389 : OAI22_X1 port map( A1 => n13646, A2 => n12448, B1 => n13587, B2 => 
                           n12442, ZN => n2886);
   U1390 : AOI221_X1 port map( B1 => n12364, B2 => n14136, C1 => n12358, C2 => 
                           n14202, A => n2875, ZN => n2868);
   U1391 : OAI22_X1 port map( A1 => n13951, A2 => n12352, B1 => n13793, B2 => 
                           n12346, ZN => n2875);
   U1392 : AOI221_X1 port map( B1 => n12460, B2 => n11719, C1 => n12454, C2 => 
                           n11539, A => n2867, ZN => n2860);
   U1393 : OAI22_X1 port map( A1 => n14345, A2 => n12448, B1 => n13586, B2 => 
                           n12442, ZN => n2867);
   U1394 : AOI221_X1 port map( B1 => n12364, B2 => n14135, C1 => n12358, C2 => 
                           n14201, A => n2856, ZN => n2849);
   U1395 : OAI22_X1 port map( A1 => n13950, A2 => n12352, B1 => n13792, B2 => 
                           n12346, ZN => n2856);
   U1396 : AOI221_X1 port map( B1 => n12460, B2 => n11720, C1 => n12454, C2 => 
                           n11540, A => n2848, ZN => n2841);
   U1397 : OAI22_X1 port map( A1 => n14344, A2 => n12448, B1 => n13585, B2 => 
                           n12442, ZN => n2848);
   U1398 : AOI221_X1 port map( B1 => n12364, B2 => n14134, C1 => n12358, C2 => 
                           n14200, A => n2837, ZN => n2830);
   U1399 : OAI22_X1 port map( A1 => n13949, A2 => n12352, B1 => n13791, B2 => 
                           n12346, ZN => n2837);
   U1400 : AOI221_X1 port map( B1 => n12460, B2 => n11721, C1 => n12454, C2 => 
                           n11541, A => n2829, ZN => n2822);
   U1401 : OAI22_X1 port map( A1 => n14343, A2 => n12448, B1 => n13584, B2 => 
                           n12442, ZN => n2829);
   U1402 : AOI221_X1 port map( B1 => n12364, B2 => n14133, C1 => n12358, C2 => 
                           n14199, A => n2818, ZN => n2811);
   U1403 : OAI22_X1 port map( A1 => n13948, A2 => n12352, B1 => n13790, B2 => 
                           n12346, ZN => n2818);
   U1404 : AOI221_X1 port map( B1 => n12460, B2 => n11722, C1 => n12454, C2 => 
                           n11542, A => n2810, ZN => n2803);
   U1405 : OAI22_X1 port map( A1 => n14342, A2 => n12448, B1 => n13583, B2 => 
                           n12442, ZN => n2810);
   U1406 : AOI221_X1 port map( B1 => n12364, B2 => n14132, C1 => n12358, C2 => 
                           n14198, A => n2799, ZN => n2792);
   U1407 : OAI22_X1 port map( A1 => n13947, A2 => n12352, B1 => n13789, B2 => 
                           n12346, ZN => n2799);
   U1408 : AOI221_X1 port map( B1 => n12460, B2 => n11723, C1 => n12454, C2 => 
                           n11543, A => n2791, ZN => n2784);
   U1409 : OAI22_X1 port map( A1 => n14341, A2 => n12448, B1 => n13582, B2 => 
                           n12442, ZN => n2791);
   U1410 : AOI221_X1 port map( B1 => n12364, B2 => n14131, C1 => n12358, C2 => 
                           n14197, A => n2780, ZN => n2773);
   U1411 : OAI22_X1 port map( A1 => n13946, A2 => n12352, B1 => n13788, B2 => 
                           n12346, ZN => n2780);
   U1412 : AOI221_X1 port map( B1 => n12460, B2 => n11724, C1 => n12454, C2 => 
                           n11544, A => n2772, ZN => n2765);
   U1413 : OAI22_X1 port map( A1 => n13645, A2 => n12448, B1 => n13581, B2 => 
                           n12442, ZN => n2772);
   U1414 : AOI221_X1 port map( B1 => n12364, B2 => n14130, C1 => n12358, C2 => 
                           n14196, A => n2761, ZN => n2754);
   U1415 : OAI22_X1 port map( A1 => n13945, A2 => n12352, B1 => n13787, B2 => 
                           n12346, ZN => n2761);
   U1416 : AOI221_X1 port map( B1 => n12460, B2 => n11725, C1 => n12454, C2 => 
                           n11545, A => n2753, ZN => n2746);
   U1417 : OAI22_X1 port map( A1 => n13644, A2 => n12448, B1 => n13580, B2 => 
                           n12442, ZN => n2753);
   U1418 : AOI221_X1 port map( B1 => n12365, B2 => n14024, C1 => n12359, C2 => 
                           n14195, A => n2742, ZN => n2735);
   U1419 : OAI22_X1 port map( A1 => n13944, A2 => n12353, B1 => n13786, B2 => 
                           n12347, ZN => n2742);
   U1420 : AOI221_X1 port map( B1 => n12461, B2 => n11726, C1 => n12455, C2 => 
                           n11546, A => n2734, ZN => n2727);
   U1421 : OAI22_X1 port map( A1 => n13643, A2 => n12449, B1 => n13579, B2 => 
                           n12443, ZN => n2734);
   U1422 : AOI221_X1 port map( B1 => n12365, B2 => n14023, C1 => n12359, C2 => 
                           n14194, A => n2723, ZN => n2716);
   U1423 : OAI22_X1 port map( A1 => n13943, A2 => n12353, B1 => n13785, B2 => 
                           n12347, ZN => n2723);
   U1424 : AOI221_X1 port map( B1 => n12461, B2 => n11727, C1 => n12455, C2 => 
                           n11547, A => n2715, ZN => n2708);
   U1425 : OAI22_X1 port map( A1 => n13642, A2 => n12449, B1 => n13578, B2 => 
                           n12443, ZN => n2715);
   U1426 : AOI221_X1 port map( B1 => n12365, B2 => n14022, C1 => n12359, C2 => 
                           n14193, A => n2704, ZN => n2697);
   U1427 : OAI22_X1 port map( A1 => n13942, A2 => n12353, B1 => n13784, B2 => 
                           n12347, ZN => n2704);
   U1428 : AOI221_X1 port map( B1 => n12461, B2 => n11728, C1 => n12455, C2 => 
                           n11548, A => n2696, ZN => n2689);
   U1429 : OAI22_X1 port map( A1 => n13641, A2 => n12449, B1 => n13577, B2 => 
                           n12443, ZN => n2696);
   U1430 : AOI221_X1 port map( B1 => n12365, B2 => n14021, C1 => n12359, C2 => 
                           n14192, A => n2685, ZN => n2678);
   U1431 : OAI22_X1 port map( A1 => n13941, A2 => n12353, B1 => n13783, B2 => 
                           n12347, ZN => n2685);
   U1432 : AOI221_X1 port map( B1 => n12461, B2 => n11729, C1 => n12455, C2 => 
                           n11549, A => n2677, ZN => n2670);
   U1433 : OAI22_X1 port map( A1 => n13640, A2 => n12449, B1 => n13576, B2 => 
                           n12443, ZN => n2677);
   U1434 : AOI221_X1 port map( B1 => n12365, B2 => n14020, C1 => n12359, C2 => 
                           n14191, A => n2666, ZN => n2659);
   U1435 : OAI22_X1 port map( A1 => n13940, A2 => n12353, B1 => n13782, B2 => 
                           n12347, ZN => n2666);
   U1436 : AOI221_X1 port map( B1 => n12461, B2 => n11730, C1 => n12455, C2 => 
                           n11550, A => n2658, ZN => n2651);
   U1437 : OAI22_X1 port map( A1 => n13639, A2 => n12449, B1 => n13575, B2 => 
                           n12443, ZN => n2658);
   U1438 : AOI221_X1 port map( B1 => n12365, B2 => n14019, C1 => n12359, C2 => 
                           n14190, A => n2647, ZN => n2640);
   U1439 : OAI22_X1 port map( A1 => n13939, A2 => n12353, B1 => n13781, B2 => 
                           n12347, ZN => n2647);
   U1440 : AOI221_X1 port map( B1 => n12461, B2 => n11731, C1 => n12455, C2 => 
                           n11551, A => n2639, ZN => n2632);
   U1441 : OAI22_X1 port map( A1 => n13638, A2 => n12449, B1 => n13574, B2 => 
                           n12443, ZN => n2639);
   U1442 : AOI221_X1 port map( B1 => n12365, B2 => n14018, C1 => n12359, C2 => 
                           n14189, A => n2628, ZN => n2621);
   U1443 : OAI22_X1 port map( A1 => n13938, A2 => n12353, B1 => n13780, B2 => 
                           n12347, ZN => n2628);
   U1444 : AOI221_X1 port map( B1 => n12461, B2 => n11732, C1 => n12455, C2 => 
                           n11552, A => n2620, ZN => n2613);
   U1445 : OAI22_X1 port map( A1 => n13637, A2 => n12449, B1 => n13573, B2 => 
                           n12443, ZN => n2620);
   U1446 : AOI221_X1 port map( B1 => n12365, B2 => n14017, C1 => n12359, C2 => 
                           n14188, A => n2609, ZN => n2602);
   U1447 : OAI22_X1 port map( A1 => n13937, A2 => n12353, B1 => n13779, B2 => 
                           n12347, ZN => n2609);
   U1448 : AOI221_X1 port map( B1 => n12461, B2 => n11733, C1 => n12455, C2 => 
                           n11553, A => n2601, ZN => n2594);
   U1449 : OAI22_X1 port map( A1 => n13636, A2 => n12449, B1 => n13572, B2 => 
                           n12443, ZN => n2601);
   U1450 : AOI221_X1 port map( B1 => n12365, B2 => n14016, C1 => n12359, C2 => 
                           n14187, A => n2590, ZN => n2583);
   U1451 : OAI22_X1 port map( A1 => n13936, A2 => n12353, B1 => n13778, B2 => 
                           n12347, ZN => n2590);
   U1452 : AOI221_X1 port map( B1 => n12461, B2 => n11734, C1 => n12455, C2 => 
                           n11554, A => n2582, ZN => n2575);
   U1453 : OAI22_X1 port map( A1 => n13635, A2 => n12449, B1 => n13571, B2 => 
                           n12443, ZN => n2582);
   U1454 : AOI221_X1 port map( B1 => n12365, B2 => n14015, C1 => n12359, C2 => 
                           n14186, A => n2571, ZN => n2564);
   U1455 : OAI22_X1 port map( A1 => n13935, A2 => n12353, B1 => n13777, B2 => 
                           n12347, ZN => n2571);
   U1456 : AOI221_X1 port map( B1 => n12461, B2 => n11735, C1 => n12455, C2 => 
                           n11555, A => n2563, ZN => n2556);
   U1457 : OAI22_X1 port map( A1 => n13634, A2 => n12449, B1 => n13570, B2 => 
                           n12443, ZN => n2563);
   U1458 : AOI221_X1 port map( B1 => n12365, B2 => n14014, C1 => n12359, C2 => 
                           n14185, A => n2552, ZN => n2545);
   U1459 : OAI22_X1 port map( A1 => n13934, A2 => n12353, B1 => n13776, B2 => 
                           n12347, ZN => n2552);
   U1460 : AOI221_X1 port map( B1 => n12461, B2 => n11736, C1 => n12455, C2 => 
                           n11556, A => n2544, ZN => n2537);
   U1461 : OAI22_X1 port map( A1 => n13633, A2 => n12449, B1 => n13569, B2 => 
                           n12443, ZN => n2544);
   U1462 : AOI221_X1 port map( B1 => n12365, B2 => n14013, C1 => n12359, C2 => 
                           n14184, A => n2533, ZN => n2526);
   U1463 : OAI22_X1 port map( A1 => n13933, A2 => n12353, B1 => n13775, B2 => 
                           n12347, ZN => n2533);
   U1464 : AOI221_X1 port map( B1 => n12461, B2 => n11737, C1 => n12455, C2 => 
                           n11557, A => n2525, ZN => n2518);
   U1465 : OAI22_X1 port map( A1 => n13632, A2 => n12449, B1 => n13568, B2 => 
                           n12443, ZN => n2525);
   U1466 : AOI221_X1 port map( B1 => n12366, B2 => n14012, C1 => n12360, C2 => 
                           n14183, A => n2514, ZN => n2507);
   U1467 : OAI22_X1 port map( A1 => n13932, A2 => n12354, B1 => n13774, B2 => 
                           n12348, ZN => n2514);
   U1468 : AOI221_X1 port map( B1 => n12462, B2 => n11738, C1 => n12456, C2 => 
                           n11558, A => n2506, ZN => n2499);
   U1469 : OAI22_X1 port map( A1 => n13631, A2 => n12450, B1 => n13567, B2 => 
                           n12444, ZN => n2506);
   U1470 : AOI221_X1 port map( B1 => n12366, B2 => n14011, C1 => n12360, C2 => 
                           n14182, A => n2495, ZN => n2488);
   U1471 : OAI22_X1 port map( A1 => n13931, A2 => n12354, B1 => n13773, B2 => 
                           n12348, ZN => n2495);
   U1472 : AOI221_X1 port map( B1 => n12462, B2 => n11739, C1 => n12456, C2 => 
                           n11559, A => n2487, ZN => n2480);
   U1473 : OAI22_X1 port map( A1 => n13630, A2 => n12450, B1 => n13566, B2 => 
                           n12444, ZN => n2487);
   U1474 : AOI221_X1 port map( B1 => n12366, B2 => n14010, C1 => n12360, C2 => 
                           n14181, A => n2476, ZN => n2469);
   U1475 : OAI22_X1 port map( A1 => n13930, A2 => n12354, B1 => n13772, B2 => 
                           n12348, ZN => n2476);
   U1476 : AOI221_X1 port map( B1 => n12462, B2 => n11740, C1 => n12456, C2 => 
                           n11560, A => n2468, ZN => n2461);
   U1477 : OAI22_X1 port map( A1 => n13629, A2 => n12450, B1 => n13565, B2 => 
                           n12444, ZN => n2468);
   U1478 : AOI221_X1 port map( B1 => n12366, B2 => n14009, C1 => n12360, C2 => 
                           n14180, A => n2457, ZN => n2450);
   U1479 : OAI22_X1 port map( A1 => n13929, A2 => n12354, B1 => n13771, B2 => 
                           n12348, ZN => n2457);
   U1480 : AOI221_X1 port map( B1 => n12462, B2 => n11741, C1 => n12456, C2 => 
                           n11561, A => n2449, ZN => n2442);
   U1481 : OAI22_X1 port map( A1 => n13628, A2 => n12450, B1 => n13564, B2 => 
                           n12444, ZN => n2449);
   U1482 : AOI221_X1 port map( B1 => n12366, B2 => n14008, C1 => n12360, C2 => 
                           n14179, A => n2438, ZN => n2431);
   U1483 : OAI22_X1 port map( A1 => n14106, A2 => n12354, B1 => n13770, B2 => 
                           n12348, ZN => n2438);
   U1484 : AOI221_X1 port map( B1 => n12462, B2 => n11742, C1 => n12456, C2 => 
                           n11562, A => n2430, ZN => n2423);
   U1485 : OAI22_X1 port map( A1 => n13627, A2 => n12450, B1 => n13563, B2 => 
                           n12444, ZN => n2430);
   U1486 : AOI221_X1 port map( B1 => n12366, B2 => n14007, C1 => n12360, C2 => 
                           n14178, A => n2419, ZN => n2412);
   U1487 : OAI22_X1 port map( A1 => n14105, A2 => n12354, B1 => n13769, B2 => 
                           n12348, ZN => n2419);
   U1488 : AOI221_X1 port map( B1 => n12462, B2 => n11743, C1 => n12456, C2 => 
                           n11563, A => n2411, ZN => n2404);
   U1489 : OAI22_X1 port map( A1 => n13626, A2 => n12450, B1 => n13562, B2 => 
                           n12444, ZN => n2411);
   U1490 : AOI221_X1 port map( B1 => n12366, B2 => n14006, C1 => n12360, C2 => 
                           n14177, A => n2400, ZN => n2393);
   U1491 : OAI22_X1 port map( A1 => n14104, A2 => n12354, B1 => n13768, B2 => 
                           n12348, ZN => n2400);
   U1492 : AOI221_X1 port map( B1 => n12462, B2 => n11744, C1 => n12456, C2 => 
                           n11564, A => n2392, ZN => n2385);
   U1493 : OAI22_X1 port map( A1 => n13625, A2 => n12450, B1 => n13561, B2 => 
                           n12444, ZN => n2392);
   U1494 : AOI221_X1 port map( B1 => n12366, B2 => n14005, C1 => n12360, C2 => 
                           n14176, A => n2381, ZN => n2374);
   U1495 : OAI22_X1 port map( A1 => n14103, A2 => n12354, B1 => n13767, B2 => 
                           n12348, ZN => n2381);
   U1496 : AOI221_X1 port map( B1 => n12462, B2 => n11745, C1 => n12456, C2 => 
                           n11565, A => n2373, ZN => n2366);
   U1497 : OAI22_X1 port map( A1 => n13624, A2 => n12450, B1 => n13560, B2 => 
                           n12444, ZN => n2373);
   U1498 : AOI221_X1 port map( B1 => n12366, B2 => n14004, C1 => n12360, C2 => 
                           n14175, A => n2362, ZN => n2355);
   U1499 : OAI22_X1 port map( A1 => n14102, A2 => n12354, B1 => n13766, B2 => 
                           n12348, ZN => n2362);
   U1500 : AOI221_X1 port map( B1 => n12462, B2 => n11746, C1 => n12456, C2 => 
                           n11566, A => n2354, ZN => n2347);
   U1501 : OAI22_X1 port map( A1 => n13623, A2 => n12450, B1 => n13559, B2 => 
                           n12444, ZN => n2354);
   U1502 : AOI221_X1 port map( B1 => n12366, B2 => n14003, C1 => n12360, C2 => 
                           n14174, A => n2343, ZN => n2336);
   U1503 : OAI22_X1 port map( A1 => n14101, A2 => n12354, B1 => n13765, B2 => 
                           n12348, ZN => n2343);
   U1504 : AOI221_X1 port map( B1 => n12462, B2 => n11747, C1 => n12456, C2 => 
                           n11567, A => n2335, ZN => n2328);
   U1505 : OAI22_X1 port map( A1 => n13622, A2 => n12450, B1 => n13558, B2 => 
                           n12444, ZN => n2335);
   U1506 : AOI221_X1 port map( B1 => n12366, B2 => n14002, C1 => n12360, C2 => 
                           n14173, A => n2324, ZN => n2317);
   U1507 : OAI22_X1 port map( A1 => n14100, A2 => n12354, B1 => n13764, B2 => 
                           n12348, ZN => n2324);
   U1508 : AOI221_X1 port map( B1 => n12462, B2 => n11748, C1 => n12456, C2 => 
                           n11568, A => n2316, ZN => n2309);
   U1509 : OAI22_X1 port map( A1 => n13621, A2 => n12450, B1 => n13557, B2 => 
                           n12444, ZN => n2316);
   U1510 : AOI221_X1 port map( B1 => n12366, B2 => n14001, C1 => n12360, C2 => 
                           n14172, A => n2305, ZN => n2298);
   U1511 : OAI22_X1 port map( A1 => n14099, A2 => n12354, B1 => n13763, B2 => 
                           n12348, ZN => n2305);
   U1512 : AOI221_X1 port map( B1 => n12462, B2 => n11749, C1 => n12456, C2 => 
                           n11569, A => n2297, ZN => n2290);
   U1513 : OAI22_X1 port map( A1 => n13620, A2 => n12450, B1 => n13556, B2 => 
                           n12444, ZN => n2297);
   U1514 : AOI221_X1 port map( B1 => n12367, B2 => n14000, C1 => n12361, C2 => 
                           n14171, A => n2286, ZN => n2279);
   U1515 : OAI22_X1 port map( A1 => n14098, A2 => n12355, B1 => n13762, B2 => 
                           n12349, ZN => n2286);
   U1516 : AOI221_X1 port map( B1 => n12463, B2 => n11750, C1 => n12457, C2 => 
                           n11570, A => n2278, ZN => n2271);
   U1517 : OAI22_X1 port map( A1 => n13619, A2 => n12451, B1 => n13555, B2 => 
                           n12445, ZN => n2278);
   U1518 : AOI221_X1 port map( B1 => n12367, B2 => n13999, C1 => n12361, C2 => 
                           n14170, A => n2267, ZN => n2260);
   U1519 : OAI22_X1 port map( A1 => n14097, A2 => n12355, B1 => n13761, B2 => 
                           n12349, ZN => n2267);
   U1520 : AOI221_X1 port map( B1 => n12463, B2 => n11751, C1 => n12457, C2 => 
                           n11571, A => n2259, ZN => n2252);
   U1521 : OAI22_X1 port map( A1 => n13618, A2 => n12451, B1 => n13554, B2 => 
                           n12445, ZN => n2259);
   U1522 : AOI221_X1 port map( B1 => n12367, B2 => n13998, C1 => n12361, C2 => 
                           n14169, A => n2248, ZN => n2241);
   U1523 : OAI22_X1 port map( A1 => n14096, A2 => n12355, B1 => n13760, B2 => 
                           n12349, ZN => n2248);
   U1524 : AOI221_X1 port map( B1 => n12463, B2 => n11752, C1 => n12457, C2 => 
                           n11572, A => n2240, ZN => n2233);
   U1525 : OAI22_X1 port map( A1 => n13617, A2 => n12451, B1 => n13553, B2 => 
                           n12445, ZN => n2240);
   U1526 : AOI221_X1 port map( B1 => n12367, B2 => n13997, C1 => n12361, C2 => 
                           n14168, A => n2229, ZN => n2222);
   U1527 : OAI22_X1 port map( A1 => n14095, A2 => n12355, B1 => n13759, B2 => 
                           n12349, ZN => n2229);
   U1528 : AOI221_X1 port map( B1 => n12463, B2 => n11753, C1 => n12457, C2 => 
                           n11573, A => n2221, ZN => n2214);
   U1529 : OAI22_X1 port map( A1 => n13616, A2 => n12451, B1 => n13552, B2 => 
                           n12445, ZN => n2221);
   U1530 : AOI221_X1 port map( B1 => n12367, B2 => n13996, C1 => n12361, C2 => 
                           n14167, A => n2210, ZN => n2203);
   U1531 : OAI22_X1 port map( A1 => n14094, A2 => n12355, B1 => n13758, B2 => 
                           n12349, ZN => n2210);
   U1532 : AOI221_X1 port map( B1 => n12463, B2 => n11754, C1 => n12457, C2 => 
                           n11574, A => n2202, ZN => n2195);
   U1533 : OAI22_X1 port map( A1 => n13615, A2 => n12451, B1 => n13551, B2 => 
                           n12445, ZN => n2202);
   U1534 : AOI221_X1 port map( B1 => n12367, B2 => n13995, C1 => n12361, C2 => 
                           n14166, A => n2191, ZN => n2184);
   U1535 : OAI22_X1 port map( A1 => n14093, A2 => n12355, B1 => n13757, B2 => 
                           n12349, ZN => n2191);
   U1536 : AOI221_X1 port map( B1 => n12463, B2 => n11755, C1 => n12457, C2 => 
                           n11575, A => n2183, ZN => n2176);
   U1537 : OAI22_X1 port map( A1 => n13614, A2 => n12451, B1 => n13550, B2 => 
                           n12445, ZN => n2183);
   U1538 : AOI221_X1 port map( B1 => n12367, B2 => n13994, C1 => n12361, C2 => 
                           n14165, A => n2172, ZN => n2165);
   U1539 : OAI22_X1 port map( A1 => n14092, A2 => n12355, B1 => n13756, B2 => 
                           n12349, ZN => n2172);
   U1540 : AOI221_X1 port map( B1 => n12463, B2 => n11756, C1 => n12457, C2 => 
                           n11576, A => n2164, ZN => n2157);
   U1541 : OAI22_X1 port map( A1 => n13613, A2 => n12451, B1 => n13549, B2 => 
                           n12445, ZN => n2164);
   U1542 : AOI221_X1 port map( B1 => n12367, B2 => n13993, C1 => n12361, C2 => 
                           n14164, A => n2153, ZN => n2146);
   U1543 : OAI22_X1 port map( A1 => n14091, A2 => n12355, B1 => n13755, B2 => 
                           n12349, ZN => n2153);
   U1544 : AOI221_X1 port map( B1 => n12463, B2 => n11757, C1 => n12457, C2 => 
                           n11577, A => n2145, ZN => n2138);
   U1545 : OAI22_X1 port map( A1 => n13612, A2 => n12451, B1 => n13548, B2 => 
                           n12445, ZN => n2145);
   U1546 : AOI221_X1 port map( B1 => n12367, B2 => n13992, C1 => n12361, C2 => 
                           n14163, A => n2134, ZN => n2127);
   U1547 : OAI22_X1 port map( A1 => n14090, A2 => n12355, B1 => n13754, B2 => 
                           n12349, ZN => n2134);
   U1548 : AOI221_X1 port map( B1 => n12463, B2 => n11758, C1 => n12457, C2 => 
                           n11578, A => n2126, ZN => n2119);
   U1549 : OAI22_X1 port map( A1 => n13611, A2 => n12451, B1 => n13547, B2 => 
                           n12445, ZN => n2126);
   U1550 : AOI221_X1 port map( B1 => n12367, B2 => n13991, C1 => n12361, C2 => 
                           n14162, A => n2115, ZN => n2108);
   U1551 : OAI22_X1 port map( A1 => n14089, A2 => n12355, B1 => n13753, B2 => 
                           n12349, ZN => n2115);
   U1552 : AOI221_X1 port map( B1 => n12463, B2 => n11759, C1 => n12457, C2 => 
                           n11579, A => n2107, ZN => n2100);
   U1553 : OAI22_X1 port map( A1 => n13610, A2 => n12451, B1 => n13546, B2 => 
                           n12445, ZN => n2107);
   U1554 : AOI221_X1 port map( B1 => n12367, B2 => n13990, C1 => n12361, C2 => 
                           n14161, A => n2096, ZN => n2089);
   U1555 : OAI22_X1 port map( A1 => n14088, A2 => n12355, B1 => n13752, B2 => 
                           n12349, ZN => n2096);
   U1556 : AOI221_X1 port map( B1 => n12463, B2 => n11760, C1 => n12457, C2 => 
                           n11580, A => n2088, ZN => n2081);
   U1557 : OAI22_X1 port map( A1 => n13609, A2 => n12451, B1 => n13545, B2 => 
                           n12445, ZN => n2088);
   U1558 : AOI221_X1 port map( B1 => n12367, B2 => n13989, C1 => n12361, C2 => 
                           n14160, A => n2077, ZN => n2070);
   U1559 : OAI22_X1 port map( A1 => n14087, A2 => n12355, B1 => n13751, B2 => 
                           n12349, ZN => n2077);
   U1560 : AOI221_X1 port map( B1 => n12463, B2 => n11761, C1 => n12457, C2 => 
                           n11581, A => n2069, ZN => n2062);
   U1561 : OAI22_X1 port map( A1 => n13608, A2 => n12451, B1 => n13544, B2 => 
                           n12445, ZN => n2069);
   U1562 : AOI221_X1 port map( B1 => n12368, B2 => n13827, C1 => n12362, C2 => 
                           n14159, A => n2058, ZN => n2051);
   U1563 : OAI22_X1 port map( A1 => n14086, A2 => n12356, B1 => n13750, B2 => 
                           n12350, ZN => n2058);
   U1564 : AOI221_X1 port map( B1 => n12464, B2 => n13864, C1 => n12458, C2 => 
                           n13868, A => n2050, ZN => n2043);
   U1565 : OAI22_X1 port map( A1 => n13607, A2 => n12452, B1 => n13543, B2 => 
                           n12446, ZN => n2050);
   U1566 : AOI221_X1 port map( B1 => n12368, B2 => n13826, C1 => n12362, C2 => 
                           n14158, A => n2039, ZN => n2032);
   U1567 : OAI22_X1 port map( A1 => n14085, A2 => n12356, B1 => n13749, B2 => 
                           n12350, ZN => n2039);
   U1568 : AOI221_X1 port map( B1 => n12464, B2 => n13863, C1 => n12458, C2 => 
                           n13867, A => n2031, ZN => n2024);
   U1569 : OAI22_X1 port map( A1 => n13606, A2 => n12452, B1 => n13542, B2 => 
                           n12446, ZN => n2031);
   U1570 : AOI221_X1 port map( B1 => n12368, B2 => n13825, C1 => n12362, C2 => 
                           n14157, A => n2020, ZN => n2013);
   U1571 : OAI22_X1 port map( A1 => n14084, A2 => n12356, B1 => n13748, B2 => 
                           n12350, ZN => n2020);
   U1572 : AOI221_X1 port map( B1 => n12464, B2 => n13862, C1 => n12458, C2 => 
                           n13866, A => n2012, ZN => n2005);
   U1573 : OAI22_X1 port map( A1 => n13605, A2 => n12452, B1 => n13541, B2 => 
                           n12446, ZN => n2012);
   U1574 : AOI221_X1 port map( B1 => n12368, B2 => n13824, C1 => n12362, C2 => 
                           n14156, A => n1999, ZN => n1978);
   U1575 : OAI22_X1 port map( A1 => n14083, A2 => n12356, B1 => n13747, B2 => 
                           n12350, ZN => n1999);
   U1576 : AOI221_X1 port map( B1 => n12464, B2 => n13861, C1 => n12458, C2 => 
                           n13865, A => n1975, ZN => n1954);
   U1577 : OAI22_X1 port map( A1 => n13604, A2 => n12452, B1 => n13540, B2 => 
                           n12446, ZN => n1975);
   U1578 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(3), A3 => n14461, 
                           ZN => n3204);
   U1579 : AOI221_X1 port map( B1 => n12387, B2 => n14079, C1 => n12381, C2 => 
                           n14126, A => n3140, ZN => n3135);
   U1580 : OAI22_X1 port map( A1 => n13743, A2 => n12375, B1 => n13727, B2 => 
                           n12369, ZN => n3140);
   U1581 : AOI221_X1 port map( B1 => n12387, B2 => n14080, C1 => n12381, C2 => 
                           n14127, A => n3121, ZN => n3116);
   U1582 : OAI22_X1 port map( A1 => n13892, A2 => n12375, B1 => n13726, B2 => 
                           n12369, ZN => n3121);
   U1583 : AOI221_X1 port map( B1 => n12387, B2 => n14076, C1 => n12381, C2 => 
                           n14123, A => n3064, ZN => n3059);
   U1584 : OAI22_X1 port map( A1 => n13889, A2 => n12375, B1 => n13723, B2 => 
                           n12369, ZN => n3064);
   U1585 : AOI221_X1 port map( B1 => n12387, B2 => n14075, C1 => n12381, C2 => 
                           n14122, A => n3045, ZN => n3040);
   U1586 : OAI22_X1 port map( A1 => n13888, A2 => n12375, B1 => n13722, B2 => 
                           n12369, ZN => n3045);
   U1587 : AOI221_X1 port map( B1 => n12387, B2 => n14074, C1 => n12381, C2 => 
                           n14121, A => n3026, ZN => n3021);
   U1588 : OAI22_X1 port map( A1 => n13887, A2 => n12375, B1 => n13721, B2 => 
                           n12369, ZN => n3026);
   U1589 : AOI221_X1 port map( B1 => n12387, B2 => n14073, C1 => n12381, C2 => 
                           n14120, A => n3007, ZN => n3002);
   U1590 : OAI22_X1 port map( A1 => n13886, A2 => n12375, B1 => n13720, B2 => 
                           n12369, ZN => n3007);
   U1591 : AOI221_X1 port map( B1 => n12387, B2 => n14072, C1 => n12381, C2 => 
                           n14119, A => n2988, ZN => n2983);
   U1592 : OAI22_X1 port map( A1 => n13885, A2 => n12375, B1 => n13719, B2 => 
                           n12369, ZN => n2988);
   U1593 : AOI221_X1 port map( B1 => n12388, B2 => n14071, C1 => n12382, C2 => 
                           n14118, A => n2969, ZN => n2964);
   U1594 : OAI22_X1 port map( A1 => n13884, A2 => n12376, B1 => n13718, B2 => 
                           n12370, ZN => n2969);
   U1595 : AOI221_X1 port map( B1 => n12388, B2 => n14070, C1 => n12382, C2 => 
                           n14117, A => n2950, ZN => n2945);
   U1596 : OAI22_X1 port map( A1 => n13883, A2 => n12376, B1 => n13717, B2 => 
                           n12370, ZN => n2950);
   U1597 : AOI221_X1 port map( B1 => n12388, B2 => n14069, C1 => n12382, C2 => 
                           n14116, A => n2931, ZN => n2926);
   U1598 : OAI22_X1 port map( A1 => n13882, A2 => n12376, B1 => n13716, B2 => 
                           n12370, ZN => n2931);
   U1599 : AOI221_X1 port map( B1 => n12388, B2 => n14068, C1 => n12382, C2 => 
                           n14115, A => n2912, ZN => n2907);
   U1600 : OAI22_X1 port map( A1 => n13881, A2 => n12376, B1 => n13715, B2 => 
                           n12370, ZN => n2912);
   U1601 : AOI221_X1 port map( B1 => n12388, B2 => n14067, C1 => n12382, C2 => 
                           n14114, A => n2893, ZN => n2888);
   U1602 : OAI22_X1 port map( A1 => n13880, A2 => n12376, B1 => n13714, B2 => 
                           n12370, ZN => n2893);
   U1603 : AOI221_X1 port map( B1 => n12388, B2 => n14066, C1 => n12382, C2 => 
                           n14113, A => n2874, ZN => n2869);
   U1604 : OAI22_X1 port map( A1 => n13879, A2 => n12376, B1 => n13713, B2 => 
                           n12370, ZN => n2874);
   U1605 : AOI221_X1 port map( B1 => n12388, B2 => n14065, C1 => n12382, C2 => 
                           n14112, A => n2855, ZN => n2850);
   U1606 : OAI22_X1 port map( A1 => n13878, A2 => n12376, B1 => n13712, B2 => 
                           n12370, ZN => n2855);
   U1607 : AOI221_X1 port map( B1 => n12388, B2 => n14064, C1 => n12382, C2 => 
                           n14111, A => n2836, ZN => n2831);
   U1608 : OAI22_X1 port map( A1 => n13877, A2 => n12376, B1 => n13711, B2 => 
                           n12370, ZN => n2836);
   U1609 : AOI221_X1 port map( B1 => n12388, B2 => n14063, C1 => n12382, C2 => 
                           n14110, A => n2817, ZN => n2812);
   U1610 : OAI22_X1 port map( A1 => n13876, A2 => n12376, B1 => n13710, B2 => 
                           n12370, ZN => n2817);
   U1611 : AOI221_X1 port map( B1 => n12388, B2 => n14062, C1 => n12382, C2 => 
                           n14109, A => n2798, ZN => n2793);
   U1612 : OAI22_X1 port map( A1 => n13875, A2 => n12376, B1 => n13709, B2 => 
                           n12370, ZN => n2798);
   U1613 : AOI221_X1 port map( B1 => n12388, B2 => n14061, C1 => n12382, C2 => 
                           n14108, A => n2779, ZN => n2774);
   U1614 : OAI22_X1 port map( A1 => n13874, A2 => n12376, B1 => n13708, B2 => 
                           n12370, ZN => n2779);
   U1615 : AOI221_X1 port map( B1 => n12388, B2 => n14060, C1 => n12382, C2 => 
                           n14107, A => n2760, ZN => n2755);
   U1616 : OAI22_X1 port map( A1 => n13873, A2 => n12376, B1 => n13707, B2 => 
                           n12370, ZN => n2760);
   U1617 : AOI221_X1 port map( B1 => n12389, B2 => n13928, C1 => n12383, C2 => 
                           n13988, A => n2741, ZN => n2736);
   U1618 : OAI22_X1 port map( A1 => n13872, A2 => n12377, B1 => n13706, B2 => 
                           n12371, ZN => n2741);
   U1619 : AOI221_X1 port map( B1 => n12389, B2 => n13927, C1 => n12383, C2 => 
                           n13987, A => n2722, ZN => n2717);
   U1620 : OAI22_X1 port map( A1 => n13871, A2 => n12377, B1 => n13705, B2 => 
                           n12371, ZN => n2722);
   U1621 : AOI221_X1 port map( B1 => n12389, B2 => n13926, C1 => n12383, C2 => 
                           n13986, A => n2703, ZN => n2698);
   U1622 : OAI22_X1 port map( A1 => n13870, A2 => n12377, B1 => n13704, B2 => 
                           n12371, ZN => n2703);
   U1623 : AOI221_X1 port map( B1 => n12389, B2 => n13925, C1 => n12383, C2 => 
                           n13985, A => n2684, ZN => n2679);
   U1624 : OAI22_X1 port map( A1 => n13869, A2 => n12377, B1 => n13703, B2 => 
                           n12371, ZN => n2684);
   U1625 : AOI221_X1 port map( B1 => n12389, B2 => n13924, C1 => n12383, C2 => 
                           n13984, A => n2665, ZN => n2660);
   U1626 : OAI22_X1 port map( A1 => n14059, A2 => n12377, B1 => n13702, B2 => 
                           n12371, ZN => n2665);
   U1627 : AOI221_X1 port map( B1 => n12389, B2 => n13923, C1 => n12383, C2 => 
                           n13983, A => n2646, ZN => n2641);
   U1628 : OAI22_X1 port map( A1 => n14058, A2 => n12377, B1 => n13701, B2 => 
                           n12371, ZN => n2646);
   U1629 : AOI221_X1 port map( B1 => n12389, B2 => n13922, C1 => n12383, C2 => 
                           n13982, A => n2627, ZN => n2622);
   U1630 : OAI22_X1 port map( A1 => n14057, A2 => n12377, B1 => n13700, B2 => 
                           n12371, ZN => n2627);
   U1631 : AOI221_X1 port map( B1 => n12389, B2 => n13921, C1 => n12383, C2 => 
                           n13981, A => n2608, ZN => n2603);
   U1632 : OAI22_X1 port map( A1 => n14056, A2 => n12377, B1 => n13699, B2 => 
                           n12371, ZN => n2608);
   U1633 : AOI221_X1 port map( B1 => n12389, B2 => n13920, C1 => n12383, C2 => 
                           n13980, A => n2589, ZN => n2584);
   U1634 : OAI22_X1 port map( A1 => n14055, A2 => n12377, B1 => n13698, B2 => 
                           n12371, ZN => n2589);
   U1635 : AOI221_X1 port map( B1 => n12389, B2 => n13919, C1 => n12383, C2 => 
                           n13979, A => n2570, ZN => n2565);
   U1636 : OAI22_X1 port map( A1 => n14054, A2 => n12377, B1 => n13697, B2 => 
                           n12371, ZN => n2570);
   U1637 : AOI221_X1 port map( B1 => n12389, B2 => n13918, C1 => n12383, C2 => 
                           n13978, A => n2551, ZN => n2546);
   U1638 : OAI22_X1 port map( A1 => n14053, A2 => n12377, B1 => n13696, B2 => 
                           n12371, ZN => n2551);
   U1639 : AOI221_X1 port map( B1 => n12389, B2 => n13917, C1 => n12383, C2 => 
                           n13977, A => n2532, ZN => n2527);
   U1640 : OAI22_X1 port map( A1 => n14052, A2 => n12377, B1 => n13695, B2 => 
                           n12371, ZN => n2532);
   U1641 : AOI221_X1 port map( B1 => n12390, B2 => n13916, C1 => n12384, C2 => 
                           n13976, A => n2513, ZN => n2508);
   U1642 : OAI22_X1 port map( A1 => n14051, A2 => n12378, B1 => n13694, B2 => 
                           n12372, ZN => n2513);
   U1643 : AOI221_X1 port map( B1 => n12390, B2 => n13915, C1 => n12384, C2 => 
                           n13975, A => n2494, ZN => n2489);
   U1644 : OAI22_X1 port map( A1 => n14050, A2 => n12378, B1 => n13693, B2 => 
                           n12372, ZN => n2494);
   U1645 : AOI221_X1 port map( B1 => n12390, B2 => n13914, C1 => n12384, C2 => 
                           n13974, A => n2475, ZN => n2470);
   U1646 : OAI22_X1 port map( A1 => n14049, A2 => n12378, B1 => n13692, B2 => 
                           n12372, ZN => n2475);
   U1647 : AOI221_X1 port map( B1 => n12390, B2 => n13913, C1 => n12384, C2 => 
                           n13973, A => n2456, ZN => n2451);
   U1648 : OAI22_X1 port map( A1 => n14048, A2 => n12378, B1 => n13691, B2 => 
                           n12372, ZN => n2456);
   U1649 : AOI221_X1 port map( B1 => n12390, B2 => n13912, C1 => n12384, C2 => 
                           n13972, A => n2437, ZN => n2432);
   U1650 : OAI22_X1 port map( A1 => n14047, A2 => n12378, B1 => n13690, B2 => 
                           n12372, ZN => n2437);
   U1651 : AOI221_X1 port map( B1 => n12390, B2 => n13911, C1 => n12384, C2 => 
                           n13971, A => n2418, ZN => n2413);
   U1652 : OAI22_X1 port map( A1 => n14046, A2 => n12378, B1 => n13689, B2 => 
                           n12372, ZN => n2418);
   U1653 : AOI221_X1 port map( B1 => n12390, B2 => n13910, C1 => n12384, C2 => 
                           n13970, A => n2399, ZN => n2394);
   U1654 : OAI22_X1 port map( A1 => n14045, A2 => n12378, B1 => n13688, B2 => 
                           n12372, ZN => n2399);
   U1655 : AOI221_X1 port map( B1 => n12390, B2 => n13909, C1 => n12384, C2 => 
                           n13969, A => n2380, ZN => n2375);
   U1656 : OAI22_X1 port map( A1 => n14044, A2 => n12378, B1 => n13687, B2 => 
                           n12372, ZN => n2380);
   U1657 : AOI221_X1 port map( B1 => n12390, B2 => n13908, C1 => n12384, C2 => 
                           n13968, A => n2361, ZN => n2356);
   U1658 : OAI22_X1 port map( A1 => n14043, A2 => n12378, B1 => n13686, B2 => 
                           n12372, ZN => n2361);
   U1659 : AOI221_X1 port map( B1 => n12390, B2 => n13907, C1 => n12384, C2 => 
                           n13967, A => n2342, ZN => n2337);
   U1660 : OAI22_X1 port map( A1 => n14042, A2 => n12378, B1 => n13685, B2 => 
                           n12372, ZN => n2342);
   U1661 : AOI221_X1 port map( B1 => n12390, B2 => n13906, C1 => n12384, C2 => 
                           n13966, A => n2323, ZN => n2318);
   U1662 : OAI22_X1 port map( A1 => n14041, A2 => n12378, B1 => n13684, B2 => 
                           n12372, ZN => n2323);
   U1663 : AOI221_X1 port map( B1 => n12390, B2 => n13905, C1 => n12384, C2 => 
                           n13965, A => n2304, ZN => n2299);
   U1664 : OAI22_X1 port map( A1 => n14040, A2 => n12378, B1 => n13683, B2 => 
                           n12372, ZN => n2304);
   U1665 : AOI221_X1 port map( B1 => n12391, B2 => n13904, C1 => n12385, C2 => 
                           n13964, A => n2285, ZN => n2280);
   U1666 : OAI22_X1 port map( A1 => n14039, A2 => n12379, B1 => n13682, B2 => 
                           n12373, ZN => n2285);
   U1667 : AOI221_X1 port map( B1 => n12391, B2 => n13903, C1 => n12385, C2 => 
                           n13963, A => n2266, ZN => n2261);
   U1668 : OAI22_X1 port map( A1 => n14038, A2 => n12379, B1 => n13681, B2 => 
                           n12373, ZN => n2266);
   U1669 : AOI221_X1 port map( B1 => n12391, B2 => n13902, C1 => n12385, C2 => 
                           n13962, A => n2247, ZN => n2242);
   U1670 : OAI22_X1 port map( A1 => n14037, A2 => n12379, B1 => n13680, B2 => 
                           n12373, ZN => n2247);
   U1671 : AOI221_X1 port map( B1 => n12391, B2 => n13901, C1 => n12385, C2 => 
                           n13961, A => n2228, ZN => n2223);
   U1672 : OAI22_X1 port map( A1 => n14036, A2 => n12379, B1 => n13679, B2 => 
                           n12373, ZN => n2228);
   U1673 : AOI221_X1 port map( B1 => n12391, B2 => n13900, C1 => n12385, C2 => 
                           n13960, A => n2209, ZN => n2204);
   U1674 : OAI22_X1 port map( A1 => n13742, A2 => n12379, B1 => n13678, B2 => 
                           n12373, ZN => n2209);
   U1675 : AOI221_X1 port map( B1 => n12391, B2 => n13899, C1 => n12385, C2 => 
                           n13959, A => n2190, ZN => n2185);
   U1676 : OAI22_X1 port map( A1 => n13741, A2 => n12379, B1 => n13677, B2 => 
                           n12373, ZN => n2190);
   U1677 : AOI221_X1 port map( B1 => n12391, B2 => n13898, C1 => n12385, C2 => 
                           n13958, A => n2171, ZN => n2166);
   U1678 : OAI22_X1 port map( A1 => n13740, A2 => n12379, B1 => n13676, B2 => 
                           n12373, ZN => n2171);
   U1679 : AOI221_X1 port map( B1 => n12391, B2 => n13897, C1 => n12385, C2 => 
                           n13957, A => n2152, ZN => n2147);
   U1680 : OAI22_X1 port map( A1 => n13739, A2 => n12379, B1 => n13675, B2 => 
                           n12373, ZN => n2152);
   U1681 : AOI221_X1 port map( B1 => n12391, B2 => n13896, C1 => n12385, C2 => 
                           n13956, A => n2133, ZN => n2128);
   U1682 : OAI22_X1 port map( A1 => n13738, A2 => n12379, B1 => n13674, B2 => 
                           n12373, ZN => n2133);
   U1683 : AOI221_X1 port map( B1 => n12391, B2 => n13895, C1 => n12385, C2 => 
                           n13955, A => n2114, ZN => n2109);
   U1684 : OAI22_X1 port map( A1 => n13737, A2 => n12379, B1 => n13673, B2 => 
                           n12373, ZN => n2114);
   U1685 : AOI221_X1 port map( B1 => n12391, B2 => n13894, C1 => n12385, C2 => 
                           n13954, A => n2095, ZN => n2090);
   U1686 : OAI22_X1 port map( A1 => n13736, A2 => n12379, B1 => n13672, B2 => 
                           n12373, ZN => n2095);
   U1687 : OAI22_X1 port map( A1 => n13107, A2 => n13173, B1 => n13093, B2 => 
                           n14408, ZN => n6719);
   U1688 : OAI22_X1 port map( A1 => n13107, A2 => n13176, B1 => n13094, B2 => 
                           n14407, ZN => n6720);
   U1689 : OAI22_X1 port map( A1 => n13107, A2 => n13179, B1 => n13091, B2 => 
                           n14406, ZN => n6721);
   U1690 : OAI22_X1 port map( A1 => n13106, A2 => n13182, B1 => n13093, B2 => 
                           n14405, ZN => n6722);
   U1691 : OAI22_X1 port map( A1 => n13106, A2 => n13185, B1 => n13094, B2 => 
                           n14404, ZN => n6723);
   U1692 : OAI22_X1 port map( A1 => n13106, A2 => n13188, B1 => n13090, B2 => 
                           n14403, ZN => n6724);
   U1693 : OAI22_X1 port map( A1 => n13106, A2 => n13191, B1 => n1914, B2 => 
                           n14402, ZN => n6725);
   U1694 : OAI22_X1 port map( A1 => n13106, A2 => n13194, B1 => n1914, B2 => 
                           n14401, ZN => n6726);
   U1695 : OAI22_X1 port map( A1 => n13105, A2 => n13197, B1 => n1914, B2 => 
                           n14400, ZN => n6727);
   U1696 : OAI22_X1 port map( A1 => n13105, A2 => n13200, B1 => n1914, B2 => 
                           n14399, ZN => n6728);
   U1697 : OAI22_X1 port map( A1 => n13105, A2 => n13203, B1 => n1914, B2 => 
                           n14398, ZN => n6729);
   U1698 : OAI22_X1 port map( A1 => n13105, A2 => n13206, B1 => n13091, B2 => 
                           n14397, ZN => n6730);
   U1699 : OAI22_X1 port map( A1 => n13105, A2 => n13209, B1 => n13091, B2 => 
                           n14396, ZN => n6731);
   U1700 : OAI22_X1 port map( A1 => n13104, A2 => n13212, B1 => n13091, B2 => 
                           n14395, ZN => n6732);
   U1701 : OAI22_X1 port map( A1 => n13104, A2 => n13215, B1 => n13091, B2 => 
                           n14394, ZN => n6733);
   U1702 : OAI22_X1 port map( A1 => n13104, A2 => n13218, B1 => n13091, B2 => 
                           n14393, ZN => n6734);
   U1703 : OAI22_X1 port map( A1 => n13104, A2 => n13221, B1 => n13091, B2 => 
                           n14392, ZN => n6735);
   U1704 : OAI22_X1 port map( A1 => n13104, A2 => n13224, B1 => n13091, B2 => 
                           n14391, ZN => n6736);
   U1705 : OAI22_X1 port map( A1 => n13103, A2 => n13227, B1 => n13091, B2 => 
                           n14390, ZN => n6737);
   U1706 : OAI22_X1 port map( A1 => n13103, A2 => n13230, B1 => n13091, B2 => 
                           n14389, ZN => n6738);
   U1707 : OAI22_X1 port map( A1 => n13103, A2 => n13233, B1 => n13091, B2 => 
                           n14388, ZN => n6739);
   U1708 : OAI22_X1 port map( A1 => n13103, A2 => n13236, B1 => n13091, B2 => 
                           n14387, ZN => n6740);
   U1709 : OAI22_X1 port map( A1 => n13103, A2 => n13239, B1 => n13091, B2 => 
                           n14386, ZN => n6741);
   U1710 : OAI22_X1 port map( A1 => n13087, A2 => n13173, B1 => n13073, B2 => 
                           n14385, ZN => n6655);
   U1711 : OAI22_X1 port map( A1 => n13087, A2 => n13176, B1 => n13074, B2 => 
                           n14384, ZN => n6656);
   U1712 : OAI22_X1 port map( A1 => n13087, A2 => n13179, B1 => n13071, B2 => 
                           n14383, ZN => n6657);
   U1713 : OAI22_X1 port map( A1 => n13086, A2 => n13182, B1 => n13073, B2 => 
                           n14382, ZN => n6658);
   U1714 : OAI22_X1 port map( A1 => n13086, A2 => n13185, B1 => n13074, B2 => 
                           n14381, ZN => n6659);
   U1715 : OAI22_X1 port map( A1 => n13086, A2 => n13188, B1 => n13070, B2 => 
                           n14380, ZN => n6660);
   U1716 : OAI22_X1 port map( A1 => n13086, A2 => n13191, B1 => n1916, B2 => 
                           n14379, ZN => n6661);
   U1717 : OAI22_X1 port map( A1 => n13086, A2 => n13194, B1 => n1916, B2 => 
                           n14378, ZN => n6662);
   U1718 : OAI22_X1 port map( A1 => n13085, A2 => n13197, B1 => n1916, B2 => 
                           n14377, ZN => n6663);
   U1719 : OAI22_X1 port map( A1 => n13085, A2 => n13200, B1 => n1916, B2 => 
                           n14376, ZN => n6664);
   U1720 : OAI22_X1 port map( A1 => n13085, A2 => n13203, B1 => n1916, B2 => 
                           n14375, ZN => n6665);
   U1721 : OAI22_X1 port map( A1 => n13085, A2 => n13206, B1 => n13071, B2 => 
                           n14374, ZN => n6666);
   U1722 : OAI22_X1 port map( A1 => n13085, A2 => n13209, B1 => n13071, B2 => 
                           n14373, ZN => n6667);
   U1723 : OAI22_X1 port map( A1 => n13084, A2 => n13212, B1 => n13071, B2 => 
                           n14372, ZN => n6668);
   U1724 : OAI22_X1 port map( A1 => n13084, A2 => n13215, B1 => n13071, B2 => 
                           n14371, ZN => n6669);
   U1725 : OAI22_X1 port map( A1 => n13084, A2 => n13218, B1 => n13071, B2 => 
                           n14370, ZN => n6670);
   U1726 : OAI22_X1 port map( A1 => n13084, A2 => n13221, B1 => n13071, B2 => 
                           n14369, ZN => n6671);
   U1727 : OAI22_X1 port map( A1 => n13084, A2 => n13224, B1 => n13071, B2 => 
                           n14368, ZN => n6672);
   U1728 : OAI22_X1 port map( A1 => n13083, A2 => n13227, B1 => n13071, B2 => 
                           n14367, ZN => n6673);
   U1729 : OAI22_X1 port map( A1 => n13083, A2 => n13230, B1 => n13071, B2 => 
                           n14366, ZN => n6674);
   U1730 : OAI22_X1 port map( A1 => n13083, A2 => n13233, B1 => n13071, B2 => 
                           n14365, ZN => n6675);
   U1731 : OAI22_X1 port map( A1 => n13083, A2 => n13236, B1 => n13071, B2 => 
                           n14364, ZN => n6676);
   U1732 : OAI22_X1 port map( A1 => n13083, A2 => n13239, B1 => n13071, B2 => 
                           n14363, ZN => n6677);
   U1733 : OAI22_X1 port map( A1 => n13107, A2 => n13170, B1 => n1914, B2 => 
                           n14362, ZN => n6718);
   U1734 : OAI22_X1 port map( A1 => n13087, A2 => n13170, B1 => n1916, B2 => 
                           n14361, ZN => n6654);
   U1735 : OAI22_X1 port map( A1 => n12966, A2 => n13182, B1 => n12951, B2 => 
                           n14360, ZN => n6274);
   U1736 : OAI22_X1 port map( A1 => n12966, A2 => n13185, B1 => n12951, B2 => 
                           n14359, ZN => n6275);
   U1737 : OAI22_X1 port map( A1 => n12966, A2 => n13188, B1 => n12951, B2 => 
                           n14358, ZN => n6276);
   U1738 : OAI22_X1 port map( A1 => n12886, A2 => n13183, B1 => n12871, B2 => 
                           n14357, ZN => n6018);
   U1739 : OAI22_X1 port map( A1 => n12886, A2 => n13186, B1 => n12871, B2 => 
                           n14356, ZN => n6019);
   U1740 : OAI22_X1 port map( A1 => n12886, A2 => n13189, B1 => n12871, B2 => 
                           n14355, ZN => n6020);
   U1741 : OAI22_X1 port map( A1 => n12886, A2 => n13192, B1 => n12871, B2 => 
                           n14354, ZN => n6021);
   U1742 : OAI22_X1 port map( A1 => n12886, A2 => n13195, B1 => n12871, B2 => 
                           n14353, ZN => n6022);
   U1743 : OAI22_X1 port map( A1 => n12885, A2 => n13198, B1 => n12871, B2 => 
                           n14352, ZN => n6023);
   U1744 : OAI22_X1 port map( A1 => n12885, A2 => n13201, B1 => n12871, B2 => 
                           n14351, ZN => n6024);
   U1745 : OAI22_X1 port map( A1 => n12885, A2 => n13204, B1 => n12871, B2 => 
                           n14350, ZN => n6025);
   U1746 : OAI22_X1 port map( A1 => n12885, A2 => n13207, B1 => n12873, B2 => 
                           n14349, ZN => n6026);
   U1747 : OAI22_X1 port map( A1 => n12885, A2 => n13210, B1 => n12874, B2 => 
                           n14348, ZN => n6027);
   U1748 : OAI22_X1 port map( A1 => n12884, A2 => n13213, B1 => n12871, B2 => 
                           n14347, ZN => n6028);
   U1749 : OAI22_X1 port map( A1 => n12884, A2 => n13216, B1 => n12873, B2 => 
                           n14346, ZN => n6029);
   U1750 : OAI22_X1 port map( A1 => n12884, A2 => n13222, B1 => n12874, B2 => 
                           n14345, ZN => n6031);
   U1751 : OAI22_X1 port map( A1 => n12884, A2 => n13225, B1 => n12870, B2 => 
                           n14344, ZN => n6032);
   U1752 : OAI22_X1 port map( A1 => n12883, A2 => n13228, B1 => n1931, B2 => 
                           n14343, ZN => n6033);
   U1753 : OAI22_X1 port map( A1 => n12883, A2 => n13231, B1 => n1931, B2 => 
                           n14342, ZN => n6034);
   U1754 : OAI22_X1 port map( A1 => n12883, A2 => n13234, B1 => n1931, B2 => 
                           n14341, ZN => n6035);
   U1755 : OAI22_X1 port map( A1 => n12966, A2 => n13191, B1 => n12951, B2 => 
                           n14340, ZN => n6277);
   U1756 : OAI22_X1 port map( A1 => n12966, A2 => n13194, B1 => n12951, B2 => 
                           n14339, ZN => n6278);
   U1757 : OAI22_X1 port map( A1 => n12965, A2 => n13197, B1 => n12951, B2 => 
                           n14338, ZN => n6279);
   U1758 : OAI22_X1 port map( A1 => n12965, A2 => n13200, B1 => n12951, B2 => 
                           n14337, ZN => n6280);
   U1759 : OAI22_X1 port map( A1 => n12965, A2 => n13203, B1 => n12951, B2 => 
                           n14336, ZN => n6281);
   U1760 : OAI22_X1 port map( A1 => n12965, A2 => n13206, B1 => n12953, B2 => 
                           n14335, ZN => n6282);
   U1761 : OAI22_X1 port map( A1 => n12965, A2 => n13209, B1 => n12954, B2 => 
                           n14334, ZN => n6283);
   U1762 : OAI22_X1 port map( A1 => n12964, A2 => n13212, B1 => n12951, B2 => 
                           n14333, ZN => n6284);
   U1763 : OAI22_X1 port map( A1 => n12964, A2 => n13215, B1 => n12953, B2 => 
                           n14332, ZN => n6285);
   U1764 : OAI22_X1 port map( A1 => n12964, A2 => n13221, B1 => n12954, B2 => 
                           n14331, ZN => n6287);
   U1765 : OAI22_X1 port map( A1 => n12964, A2 => n13224, B1 => n12950, B2 => 
                           n14330, ZN => n6288);
   U1766 : OAI22_X1 port map( A1 => n12963, A2 => n13227, B1 => n1927, B2 => 
                           n14329, ZN => n6289);
   U1767 : OAI22_X1 port map( A1 => n13376, A2 => n13173, B1 => n13362, B2 => 
                           n14328, ZN => n6975);
   U1768 : OAI22_X1 port map( A1 => n13376, A2 => n13176, B1 => n13363, B2 => 
                           n14327, ZN => n6976);
   U1769 : OAI22_X1 port map( A1 => n13376, A2 => n13179, B1 => n13360, B2 => 
                           n14326, ZN => n6977);
   U1770 : OAI22_X1 port map( A1 => n13375, A2 => n13182, B1 => n13362, B2 => 
                           n14325, ZN => n6978);
   U1771 : OAI22_X1 port map( A1 => n13375, A2 => n13185, B1 => n13363, B2 => 
                           n14324, ZN => n6979);
   U1772 : OAI22_X1 port map( A1 => n13375, A2 => n13194, B1 => n13359, B2 => 
                           n14323, ZN => n6982);
   U1773 : OAI22_X1 port map( A1 => n13375, A2 => n13188, B1 => n1842, B2 => 
                           n14311, ZN => n6980);
   U1774 : OAI22_X1 port map( A1 => n13375, A2 => n13191, B1 => n1842, B2 => 
                           n14310, ZN => n6981);
   U1775 : OAI22_X1 port map( A1 => n13374, A2 => n13197, B1 => n1842, B2 => 
                           n14309, ZN => n6983);
   U1776 : OAI22_X1 port map( A1 => n13374, A2 => n13200, B1 => n1842, B2 => 
                           n14308, ZN => n6984);
   U1777 : OAI22_X1 port map( A1 => n13374, A2 => n13203, B1 => n1842, B2 => 
                           n14307, ZN => n6985);
   U1778 : OAI22_X1 port map( A1 => n13374, A2 => n13206, B1 => n13360, B2 => 
                           n14306, ZN => n6986);
   U1779 : OAI22_X1 port map( A1 => n13374, A2 => n13209, B1 => n13360, B2 => 
                           n14305, ZN => n6987);
   U1780 : OAI22_X1 port map( A1 => n13373, A2 => n13212, B1 => n13360, B2 => 
                           n14304, ZN => n6988);
   U1781 : OAI22_X1 port map( A1 => n13373, A2 => n13215, B1 => n13360, B2 => 
                           n14303, ZN => n6989);
   U1782 : OAI22_X1 port map( A1 => n13373, A2 => n13218, B1 => n13360, B2 => 
                           n14302, ZN => n6990);
   U1783 : OAI22_X1 port map( A1 => n13373, A2 => n13221, B1 => n13360, B2 => 
                           n14301, ZN => n6991);
   U1784 : OAI22_X1 port map( A1 => n13373, A2 => n13224, B1 => n13360, B2 => 
                           n14300, ZN => n6992);
   U1785 : OAI22_X1 port map( A1 => n13372, A2 => n13227, B1 => n13360, B2 => 
                           n14299, ZN => n6993);
   U1786 : OAI22_X1 port map( A1 => n13372, A2 => n13230, B1 => n13360, B2 => 
                           n14298, ZN => n6994);
   U1787 : OAI22_X1 port map( A1 => n13372, A2 => n13233, B1 => n13360, B2 => 
                           n14297, ZN => n6995);
   U1788 : OAI22_X1 port map( A1 => n13372, A2 => n13236, B1 => n13360, B2 => 
                           n14296, ZN => n6996);
   U1789 : OAI22_X1 port map( A1 => n13372, A2 => n13239, B1 => n13360, B2 => 
                           n14295, ZN => n6997);
   U1790 : OAI22_X1 port map( A1 => n13376, A2 => n13170, B1 => n1842, B2 => 
                           n14216, ZN => n6974);
   U1791 : OAI22_X1 port map( A1 => n12611, A2 => n13187, B1 => n12597, B2 => 
                           n14035, ZN => n5123);
   U1792 : OAI22_X1 port map( A1 => n12611, A2 => n13190, B1 => n12598, B2 => 
                           n14034, ZN => n5124);
   U1793 : OAI22_X1 port map( A1 => n12611, A2 => n13193, B1 => n12599, B2 => 
                           n14033, ZN => n5125);
   U1794 : OAI22_X1 port map( A1 => n12611, A2 => n13196, B1 => n12597, B2 => 
                           n14032, ZN => n5126);
   U1795 : OAI22_X1 port map( A1 => n12610, A2 => n13199, B1 => n12598, B2 => 
                           n14031, ZN => n5127);
   U1796 : OAI22_X1 port map( A1 => n12610, A2 => n13202, B1 => n12596, B2 => 
                           n14030, ZN => n5128);
   U1797 : OAI22_X1 port map( A1 => n12610, A2 => n13205, B1 => n1947, B2 => 
                           n14029, ZN => n5129);
   U1798 : OAI22_X1 port map( A1 => n12610, A2 => n13208, B1 => n12599, B2 => 
                           n14028, ZN => n5130);
   U1799 : OAI22_X1 port map( A1 => n12610, A2 => n13211, B1 => n12596, B2 => 
                           n14027, ZN => n5131);
   U1800 : OAI22_X1 port map( A1 => n12609, A2 => n13214, B1 => n12596, B2 => 
                           n14026, ZN => n5132);
   U1801 : OAI22_X1 port map( A1 => n12609, A2 => n13217, B1 => n1947, B2 => 
                           n14025, ZN => n5133);
   U1802 : OAI22_X1 port map( A1 => n12609, A2 => n13220, B1 => n1947, B2 => 
                           n13952, ZN => n5134);
   U1803 : OAI22_X1 port map( A1 => n12609, A2 => n13223, B1 => n1947, B2 => 
                           n13951, ZN => n5135);
   U1804 : OAI22_X1 port map( A1 => n12609, A2 => n13226, B1 => n1947, B2 => 
                           n13950, ZN => n5136);
   U1805 : OAI22_X1 port map( A1 => n12608, A2 => n13229, B1 => n1947, B2 => 
                           n13949, ZN => n5137);
   U1806 : OAI22_X1 port map( A1 => n12608, A2 => n13232, B1 => n12596, B2 => 
                           n13948, ZN => n5138);
   U1807 : OAI22_X1 port map( A1 => n12608, A2 => n13235, B1 => n12596, B2 => 
                           n13947, ZN => n5139);
   U1808 : OAI22_X1 port map( A1 => n12608, A2 => n13238, B1 => n12596, B2 => 
                           n13946, ZN => n5140);
   U1809 : OAI22_X1 port map( A1 => n12608, A2 => n13241, B1 => n12596, B2 => 
                           n13945, ZN => n5141);
   U1810 : OAI22_X1 port map( A1 => n12687, A2 => n13184, B1 => n12673, B2 => 
                           n13892, ZN => n5378);
   U1811 : OAI22_X1 port map( A1 => n12687, A2 => n13187, B1 => n12675, B2 => 
                           n13891, ZN => n5379);
   U1812 : OAI22_X1 port map( A1 => n12687, A2 => n13190, B1 => n12674, B2 => 
                           n13890, ZN => n5380);
   U1813 : OAI22_X1 port map( A1 => n12687, A2 => n13193, B1 => n12673, B2 => 
                           n13889, ZN => n5381);
   U1814 : OAI22_X1 port map( A1 => n12687, A2 => n13196, B1 => n12675, B2 => 
                           n13888, ZN => n5382);
   U1815 : OAI22_X1 port map( A1 => n12686, A2 => n13199, B1 => n12672, B2 => 
                           n13887, ZN => n5383);
   U1816 : OAI22_X1 port map( A1 => n12686, A2 => n13202, B1 => n1943, B2 => 
                           n13886, ZN => n5384);
   U1817 : OAI22_X1 port map( A1 => n12686, A2 => n13205, B1 => n1943, B2 => 
                           n13885, ZN => n5385);
   U1818 : OAI22_X1 port map( A1 => n12686, A2 => n13208, B1 => n12674, B2 => 
                           n13884, ZN => n5386);
   U1819 : OAI22_X1 port map( A1 => n12686, A2 => n13211, B1 => n12672, B2 => 
                           n13883, ZN => n5387);
   U1820 : OAI22_X1 port map( A1 => n12685, A2 => n13214, B1 => n12672, B2 => 
                           n13882, ZN => n5388);
   U1821 : OAI22_X1 port map( A1 => n12685, A2 => n13217, B1 => n1943, B2 => 
                           n13881, ZN => n5389);
   U1822 : OAI22_X1 port map( A1 => n12685, A2 => n13220, B1 => n1943, B2 => 
                           n13880, ZN => n5390);
   U1823 : OAI22_X1 port map( A1 => n12685, A2 => n13223, B1 => n1943, B2 => 
                           n13879, ZN => n5391);
   U1824 : OAI22_X1 port map( A1 => n12685, A2 => n13226, B1 => n1943, B2 => 
                           n13878, ZN => n5392);
   U1825 : OAI22_X1 port map( A1 => n12684, A2 => n13229, B1 => n1943, B2 => 
                           n13877, ZN => n5393);
   U1826 : OAI22_X1 port map( A1 => n12684, A2 => n13232, B1 => n12672, B2 => 
                           n13876, ZN => n5394);
   U1827 : OAI22_X1 port map( A1 => n12684, A2 => n13235, B1 => n12672, B2 => 
                           n13875, ZN => n5395);
   U1828 : OAI22_X1 port map( A1 => n12684, A2 => n13238, B1 => n12672, B2 => 
                           n13874, ZN => n5396);
   U1829 : OAI22_X1 port map( A1 => n12684, A2 => n13241, B1 => n12672, B2 => 
                           n13873, ZN => n5397);
   U1830 : OAI22_X1 port map( A1 => n12612, A2 => n13172, B1 => n1947, B2 => 
                           n13815, ZN => n5118);
   U1831 : OAI22_X1 port map( A1 => n12612, A2 => n13175, B1 => n1947, B2 => 
                           n13814, ZN => n5119);
   U1832 : OAI22_X1 port map( A1 => n12612, A2 => n13178, B1 => n1947, B2 => 
                           n13813, ZN => n5120);
   U1833 : OAI22_X1 port map( A1 => n12612, A2 => n13181, B1 => n1947, B2 => 
                           n13812, ZN => n5121);
   U1834 : OAI22_X1 port map( A1 => n12611, A2 => n13184, B1 => n1947, B2 => 
                           n13811, ZN => n5122);
   U1835 : OAI22_X1 port map( A1 => n12631, A2 => n13172, B1 => n12616, B2 => 
                           n13810, ZN => n5182);
   U1836 : OAI22_X1 port map( A1 => n12631, A2 => n13175, B1 => n12615, B2 => 
                           n13809, ZN => n5183);
   U1837 : OAI22_X1 port map( A1 => n12631, A2 => n13178, B1 => n12615, B2 => 
                           n13808, ZN => n5184);
   U1838 : OAI22_X1 port map( A1 => n12631, A2 => n13181, B1 => n1946, B2 => 
                           n13807, ZN => n5185);
   U1839 : OAI22_X1 port map( A1 => n12630, A2 => n13184, B1 => n1946, B2 => 
                           n13806, ZN => n5186);
   U1840 : OAI22_X1 port map( A1 => n12630, A2 => n13187, B1 => n1946, B2 => 
                           n13805, ZN => n5187);
   U1841 : OAI22_X1 port map( A1 => n12630, A2 => n13190, B1 => n1946, B2 => 
                           n13804, ZN => n5188);
   U1842 : OAI22_X1 port map( A1 => n12630, A2 => n13193, B1 => n1946, B2 => 
                           n13803, ZN => n5189);
   U1843 : OAI22_X1 port map( A1 => n12630, A2 => n13196, B1 => n12615, B2 => 
                           n13802, ZN => n5190);
   U1844 : OAI22_X1 port map( A1 => n12629, A2 => n13199, B1 => n12615, B2 => 
                           n13801, ZN => n5191);
   U1845 : OAI22_X1 port map( A1 => n12629, A2 => n13202, B1 => n12615, B2 => 
                           n13800, ZN => n5192);
   U1846 : OAI22_X1 port map( A1 => n12629, A2 => n13205, B1 => n12615, B2 => 
                           n13799, ZN => n5193);
   U1847 : OAI22_X1 port map( A1 => n12629, A2 => n13208, B1 => n12617, B2 => 
                           n13798, ZN => n5194);
   U1848 : OAI22_X1 port map( A1 => n12629, A2 => n13211, B1 => n12618, B2 => 
                           n13797, ZN => n5195);
   U1849 : OAI22_X1 port map( A1 => n12628, A2 => n13214, B1 => n12616, B2 => 
                           n13796, ZN => n5196);
   U1850 : OAI22_X1 port map( A1 => n12628, A2 => n13217, B1 => n12617, B2 => 
                           n13795, ZN => n5197);
   U1851 : OAI22_X1 port map( A1 => n12628, A2 => n13220, B1 => n12618, B2 => 
                           n13794, ZN => n5198);
   U1852 : OAI22_X1 port map( A1 => n12628, A2 => n13223, B1 => n12615, B2 => 
                           n13793, ZN => n5199);
   U1853 : OAI22_X1 port map( A1 => n12628, A2 => n13226, B1 => n1946, B2 => 
                           n13792, ZN => n5200);
   U1854 : OAI22_X1 port map( A1 => n12627, A2 => n13229, B1 => n1946, B2 => 
                           n13791, ZN => n5201);
   U1855 : OAI22_X1 port map( A1 => n12627, A2 => n13232, B1 => n1946, B2 => 
                           n13790, ZN => n5202);
   U1856 : OAI22_X1 port map( A1 => n12627, A2 => n13235, B1 => n1946, B2 => 
                           n13789, ZN => n5203);
   U1857 : OAI22_X1 port map( A1 => n12627, A2 => n13238, B1 => n1946, B2 => 
                           n13788, ZN => n5204);
   U1858 : OAI22_X1 port map( A1 => n12627, A2 => n13241, B1 => n1946, B2 => 
                           n13787, ZN => n5205);
   U1859 : OAI22_X1 port map( A1 => n12688, A2 => n13172, B1 => n1943, B2 => 
                           n13746, ZN => n5374);
   U1860 : OAI22_X1 port map( A1 => n12688, A2 => n13175, B1 => n1943, B2 => 
                           n13745, ZN => n5375);
   U1861 : OAI22_X1 port map( A1 => n12688, A2 => n13178, B1 => n1943, B2 => 
                           n13744, ZN => n5376);
   U1862 : OAI22_X1 port map( A1 => n12688, A2 => n13181, B1 => n1943, B2 => 
                           n13743, ZN => n5377);
   U1863 : OAI22_X1 port map( A1 => n12707, A2 => n13172, B1 => n12692, B2 => 
                           n13730, ZN => n5438);
   U1864 : OAI22_X1 port map( A1 => n12707, A2 => n13175, B1 => n12691, B2 => 
                           n13729, ZN => n5439);
   U1865 : OAI22_X1 port map( A1 => n12707, A2 => n13178, B1 => n12691, B2 => 
                           n13728, ZN => n5440);
   U1866 : OAI22_X1 port map( A1 => n12707, A2 => n13181, B1 => n1941, B2 => 
                           n13727, ZN => n5441);
   U1867 : OAI22_X1 port map( A1 => n12706, A2 => n13184, B1 => n1941, B2 => 
                           n13726, ZN => n5442);
   U1868 : OAI22_X1 port map( A1 => n12706, A2 => n13187, B1 => n1941, B2 => 
                           n13725, ZN => n5443);
   U1869 : OAI22_X1 port map( A1 => n12706, A2 => n13190, B1 => n1941, B2 => 
                           n13724, ZN => n5444);
   U1870 : OAI22_X1 port map( A1 => n12706, A2 => n13193, B1 => n1941, B2 => 
                           n13723, ZN => n5445);
   U1871 : OAI22_X1 port map( A1 => n12706, A2 => n13196, B1 => n12691, B2 => 
                           n13722, ZN => n5446);
   U1872 : OAI22_X1 port map( A1 => n12705, A2 => n13199, B1 => n12691, B2 => 
                           n13721, ZN => n5447);
   U1873 : OAI22_X1 port map( A1 => n12705, A2 => n13202, B1 => n12691, B2 => 
                           n13720, ZN => n5448);
   U1874 : OAI22_X1 port map( A1 => n12705, A2 => n13205, B1 => n12691, B2 => 
                           n13719, ZN => n5449);
   U1875 : OAI22_X1 port map( A1 => n12705, A2 => n13208, B1 => n12693, B2 => 
                           n13718, ZN => n5450);
   U1876 : OAI22_X1 port map( A1 => n12705, A2 => n13211, B1 => n12694, B2 => 
                           n13717, ZN => n5451);
   U1877 : OAI22_X1 port map( A1 => n12704, A2 => n13214, B1 => n12692, B2 => 
                           n13716, ZN => n5452);
   U1878 : OAI22_X1 port map( A1 => n12704, A2 => n13217, B1 => n12693, B2 => 
                           n13715, ZN => n5453);
   U1879 : OAI22_X1 port map( A1 => n12704, A2 => n13220, B1 => n12694, B2 => 
                           n13714, ZN => n5454);
   U1880 : OAI22_X1 port map( A1 => n12704, A2 => n13223, B1 => n12691, B2 => 
                           n13713, ZN => n5455);
   U1881 : OAI22_X1 port map( A1 => n12704, A2 => n13226, B1 => n1941, B2 => 
                           n13712, ZN => n5456);
   U1882 : OAI22_X1 port map( A1 => n12703, A2 => n13229, B1 => n1941, B2 => 
                           n13711, ZN => n5457);
   U1883 : OAI22_X1 port map( A1 => n12703, A2 => n13232, B1 => n1941, B2 => 
                           n13710, ZN => n5458);
   U1884 : OAI22_X1 port map( A1 => n12703, A2 => n13235, B1 => n1941, B2 => 
                           n13709, ZN => n5459);
   U1885 : OAI22_X1 port map( A1 => n12703, A2 => n13238, B1 => n1941, B2 => 
                           n13708, ZN => n5460);
   U1886 : OAI22_X1 port map( A1 => n12703, A2 => n13241, B1 => n1941, B2 => 
                           n13707, ZN => n5461);
   U1887 : OAI22_X1 port map( A1 => n12887, A2 => n13171, B1 => n12871, B2 => 
                           n13650, ZN => n6014);
   U1888 : OAI22_X1 port map( A1 => n12887, A2 => n13174, B1 => n12871, B2 => 
                           n13649, ZN => n6015);
   U1889 : OAI22_X1 port map( A1 => n12887, A2 => n13177, B1 => n12871, B2 => 
                           n13648, ZN => n6016);
   U1890 : OAI22_X1 port map( A1 => n12887, A2 => n13180, B1 => n12871, B2 => 
                           n13647, ZN => n6017);
   U1891 : OAI22_X1 port map( A1 => n12884, A2 => n13219, B1 => n1931, B2 => 
                           n13646, ZN => n6030);
   U1892 : OAI22_X1 port map( A1 => n12883, A2 => n13237, B1 => n1931, B2 => 
                           n13645, ZN => n6036);
   U1893 : OAI22_X1 port map( A1 => n12883, A2 => n13240, B1 => n1931, B2 => 
                           n13644, ZN => n6037);
   U1894 : OAI22_X1 port map( A1 => n12907, A2 => n13171, B1 => n12891, B2 => 
                           n13603, ZN => n6078);
   U1895 : OAI22_X1 port map( A1 => n12907, A2 => n13174, B1 => n12891, B2 => 
                           n13602, ZN => n6079);
   U1896 : OAI22_X1 port map( A1 => n12907, A2 => n13177, B1 => n12891, B2 => 
                           n13601, ZN => n6080);
   U1897 : OAI22_X1 port map( A1 => n12907, A2 => n13180, B1 => n12891, B2 => 
                           n13600, ZN => n6081);
   U1898 : OAI22_X1 port map( A1 => n12906, A2 => n13183, B1 => n12891, B2 => 
                           n13599, ZN => n6082);
   U1899 : OAI22_X1 port map( A1 => n12906, A2 => n13186, B1 => n12891, B2 => 
                           n13598, ZN => n6083);
   U1900 : OAI22_X1 port map( A1 => n12906, A2 => n13189, B1 => n12891, B2 => 
                           n13597, ZN => n6084);
   U1901 : OAI22_X1 port map( A1 => n12906, A2 => n13192, B1 => n12891, B2 => 
                           n13596, ZN => n6085);
   U1902 : OAI22_X1 port map( A1 => n12906, A2 => n13195, B1 => n12891, B2 => 
                           n13595, ZN => n6086);
   U1903 : OAI22_X1 port map( A1 => n12905, A2 => n13198, B1 => n12891, B2 => 
                           n13594, ZN => n6087);
   U1904 : OAI22_X1 port map( A1 => n12905, A2 => n13201, B1 => n12891, B2 => 
                           n13593, ZN => n6088);
   U1905 : OAI22_X1 port map( A1 => n12905, A2 => n13204, B1 => n12891, B2 => 
                           n13592, ZN => n6089);
   U1906 : OAI22_X1 port map( A1 => n12905, A2 => n13207, B1 => n12893, B2 => 
                           n13591, ZN => n6090);
   U1907 : OAI22_X1 port map( A1 => n12905, A2 => n13210, B1 => n12894, B2 => 
                           n13590, ZN => n6091);
   U1908 : OAI22_X1 port map( A1 => n12904, A2 => n13213, B1 => n12891, B2 => 
                           n13589, ZN => n6092);
   U1909 : OAI22_X1 port map( A1 => n12904, A2 => n13216, B1 => n12893, B2 => 
                           n13588, ZN => n6093);
   U1910 : OAI22_X1 port map( A1 => n12904, A2 => n13219, B1 => n12894, B2 => 
                           n13587, ZN => n6094);
   U1911 : OAI22_X1 port map( A1 => n12904, A2 => n13222, B1 => n12890, B2 => 
                           n13586, ZN => n6095);
   U1912 : OAI22_X1 port map( A1 => n12904, A2 => n13225, B1 => n1930, B2 => 
                           n13585, ZN => n6096);
   U1913 : OAI22_X1 port map( A1 => n12903, A2 => n13228, B1 => n1930, B2 => 
                           n13584, ZN => n6097);
   U1914 : OAI22_X1 port map( A1 => n12903, A2 => n13231, B1 => n1930, B2 => 
                           n13583, ZN => n6098);
   U1915 : OAI22_X1 port map( A1 => n12903, A2 => n13234, B1 => n1930, B2 => 
                           n13582, ZN => n6099);
   U1916 : OAI22_X1 port map( A1 => n12903, A2 => n13237, B1 => n1930, B2 => 
                           n13581, ZN => n6100);
   U1917 : OAI22_X1 port map( A1 => n12903, A2 => n13240, B1 => n1930, B2 => 
                           n13580, ZN => n6101);
   U1918 : OAI22_X1 port map( A1 => n12967, A2 => n13170, B1 => n12951, B2 => 
                           n13539, ZN => n6270);
   U1919 : OAI22_X1 port map( A1 => n12967, A2 => n13173, B1 => n12951, B2 => 
                           n13538, ZN => n6271);
   U1920 : OAI22_X1 port map( A1 => n12967, A2 => n13176, B1 => n12951, B2 => 
                           n13537, ZN => n6272);
   U1921 : OAI22_X1 port map( A1 => n12967, A2 => n13179, B1 => n12951, B2 => 
                           n13536, ZN => n6273);
   U1922 : OAI22_X1 port map( A1 => n12964, A2 => n13218, B1 => n1927, B2 => 
                           n13535, ZN => n6286);
   U1923 : OAI22_X1 port map( A1 => n12963, A2 => n13230, B1 => n1927, B2 => 
                           n13534, ZN => n6290);
   U1924 : OAI22_X1 port map( A1 => n12963, A2 => n13233, B1 => n1927, B2 => 
                           n13533, ZN => n6291);
   U1925 : OAI22_X1 port map( A1 => n12963, A2 => n13236, B1 => n1927, B2 => 
                           n13532, ZN => n6292);
   U1926 : OAI22_X1 port map( A1 => n12963, A2 => n13239, B1 => n1927, B2 => 
                           n13531, ZN => n6293);
   U1927 : OAI22_X1 port map( A1 => n12987, A2 => n13170, B1 => n12971, B2 => 
                           n13494, ZN => n6334);
   U1928 : OAI22_X1 port map( A1 => n12987, A2 => n13173, B1 => n12971, B2 => 
                           n13493, ZN => n6335);
   U1929 : OAI22_X1 port map( A1 => n12987, A2 => n13176, B1 => n12971, B2 => 
                           n13492, ZN => n6336);
   U1930 : OAI22_X1 port map( A1 => n12987, A2 => n13179, B1 => n12971, B2 => 
                           n13491, ZN => n6337);
   U1931 : OAI22_X1 port map( A1 => n12986, A2 => n13182, B1 => n12971, B2 => 
                           n13490, ZN => n6338);
   U1932 : OAI22_X1 port map( A1 => n12986, A2 => n13185, B1 => n12971, B2 => 
                           n13489, ZN => n6339);
   U1933 : OAI22_X1 port map( A1 => n12986, A2 => n13188, B1 => n12971, B2 => 
                           n13488, ZN => n6340);
   U1934 : OAI22_X1 port map( A1 => n12986, A2 => n13191, B1 => n12971, B2 => 
                           n13487, ZN => n6341);
   U1935 : OAI22_X1 port map( A1 => n12986, A2 => n13194, B1 => n12971, B2 => 
                           n13486, ZN => n6342);
   U1936 : OAI22_X1 port map( A1 => n12985, A2 => n13197, B1 => n12971, B2 => 
                           n13485, ZN => n6343);
   U1937 : OAI22_X1 port map( A1 => n12985, A2 => n13200, B1 => n12971, B2 => 
                           n13484, ZN => n6344);
   U1938 : OAI22_X1 port map( A1 => n12985, A2 => n13203, B1 => n12971, B2 => 
                           n13483, ZN => n6345);
   U1939 : OAI22_X1 port map( A1 => n12985, A2 => n13206, B1 => n12973, B2 => 
                           n13482, ZN => n6346);
   U1940 : OAI22_X1 port map( A1 => n12985, A2 => n13209, B1 => n12974, B2 => 
                           n13481, ZN => n6347);
   U1941 : OAI22_X1 port map( A1 => n12984, A2 => n13212, B1 => n12971, B2 => 
                           n13480, ZN => n6348);
   U1942 : OAI22_X1 port map( A1 => n12984, A2 => n13215, B1 => n12973, B2 => 
                           n13479, ZN => n6349);
   U1943 : OAI22_X1 port map( A1 => n12984, A2 => n13218, B1 => n12974, B2 => 
                           n13478, ZN => n6350);
   U1944 : OAI22_X1 port map( A1 => n12984, A2 => n13221, B1 => n12970, B2 => 
                           n13477, ZN => n6351);
   U1945 : OAI22_X1 port map( A1 => n12984, A2 => n13224, B1 => n1926, B2 => 
                           n13476, ZN => n6352);
   U1946 : OAI22_X1 port map( A1 => n12983, A2 => n13227, B1 => n1926, B2 => 
                           n13475, ZN => n6353);
   U1947 : OAI22_X1 port map( A1 => n12983, A2 => n13230, B1 => n1926, B2 => 
                           n13474, ZN => n6354);
   U1948 : OAI22_X1 port map( A1 => n12983, A2 => n13233, B1 => n1926, B2 => 
                           n13473, ZN => n6355);
   U1949 : OAI22_X1 port map( A1 => n12983, A2 => n13236, B1 => n1926, B2 => 
                           n13472, ZN => n6356);
   U1950 : OAI22_X1 port map( A1 => n12983, A2 => n13239, B1 => n1926, B2 => 
                           n13471, ZN => n6357);
   U1951 : OAI22_X1 port map( A1 => n13167, A2 => n13170, B1 => n13151, B2 => 
                           n13430, ZN => n6910);
   U1952 : OAI22_X1 port map( A1 => n13167, A2 => n13173, B1 => n13151, B2 => 
                           n13429, ZN => n6911);
   U1953 : OAI22_X1 port map( A1 => n13167, A2 => n13176, B1 => n13151, B2 => 
                           n13428, ZN => n6912);
   U1954 : OAI22_X1 port map( A1 => n13167, A2 => n13179, B1 => n13151, B2 => 
                           n13427, ZN => n6913);
   U1955 : OAI22_X1 port map( A1 => n13166, A2 => n13182, B1 => n13151, B2 => 
                           n13426, ZN => n6914);
   U1956 : OAI22_X1 port map( A1 => n13166, A2 => n13185, B1 => n13151, B2 => 
                           n13425, ZN => n6915);
   U1957 : OAI22_X1 port map( A1 => n13166, A2 => n13188, B1 => n13151, B2 => 
                           n13424, ZN => n6916);
   U1958 : OAI22_X1 port map( A1 => n13166, A2 => n13191, B1 => n13151, B2 => 
                           n13423, ZN => n6917);
   U1959 : OAI22_X1 port map( A1 => n13166, A2 => n13194, B1 => n13151, B2 => 
                           n13422, ZN => n6918);
   U1960 : OAI22_X1 port map( A1 => n13165, A2 => n13197, B1 => n13151, B2 => 
                           n13421, ZN => n6919);
   U1961 : OAI22_X1 port map( A1 => n13165, A2 => n13200, B1 => n13151, B2 => 
                           n13420, ZN => n6920);
   U1962 : OAI22_X1 port map( A1 => n13165, A2 => n13203, B1 => n13151, B2 => 
                           n13419, ZN => n6921);
   U1963 : OAI22_X1 port map( A1 => n13165, A2 => n13206, B1 => n13153, B2 => 
                           n13418, ZN => n6922);
   U1964 : OAI22_X1 port map( A1 => n13165, A2 => n13209, B1 => n13152, B2 => 
                           n13417, ZN => n6923);
   U1965 : OAI22_X1 port map( A1 => n13164, A2 => n13212, B1 => n13151, B2 => 
                           n13416, ZN => n6924);
   U1966 : OAI22_X1 port map( A1 => n13164, A2 => n13215, B1 => n13153, B2 => 
                           n13415, ZN => n6925);
   U1967 : OAI22_X1 port map( A1 => n13164, A2 => n13218, B1 => n13152, B2 => 
                           n13414, ZN => n6926);
   U1968 : OAI22_X1 port map( A1 => n13164, A2 => n13221, B1 => n13150, B2 => 
                           n13413, ZN => n6927);
   U1969 : OAI22_X1 port map( A1 => n13164, A2 => n13224, B1 => n1908, B2 => 
                           n13412, ZN => n6928);
   U1970 : OAI22_X1 port map( A1 => n13163, A2 => n13227, B1 => n1908, B2 => 
                           n13411, ZN => n6929);
   U1971 : OAI22_X1 port map( A1 => n13163, A2 => n13230, B1 => n1908, B2 => 
                           n13410, ZN => n6930);
   U1972 : OAI22_X1 port map( A1 => n13163, A2 => n13233, B1 => n1908, B2 => 
                           n13409, ZN => n6931);
   U1973 : OAI22_X1 port map( A1 => n13163, A2 => n13236, B1 => n1908, B2 => 
                           n13408, ZN => n6932);
   U1974 : OAI22_X1 port map( A1 => n13163, A2 => n13239, B1 => n1908, B2 => 
                           n13407, ZN => n6933);
   U1975 : OAI22_X1 port map( A1 => n12959, A2 => n13287, B1 => n12953, B2 => 
                           n14460, ZN => n6309);
   U1976 : OAI22_X1 port map( A1 => n12959, A2 => n13290, B1 => n12953, B2 => 
                           n14459, ZN => n6310);
   U1977 : OAI22_X1 port map( A1 => n12959, A2 => n13293, B1 => n12953, B2 => 
                           n14458, ZN => n6311);
   U1978 : OAI22_X1 port map( A1 => n12959, A2 => n13296, B1 => n12953, B2 => 
                           n14457, ZN => n6312);
   U1979 : OAI22_X1 port map( A1 => n13370, A2 => n13260, B1 => n13361, B2 => 
                           n14456, ZN => n7004);
   U1980 : OAI22_X1 port map( A1 => n13370, A2 => n13263, B1 => n13361, B2 => 
                           n14455, ZN => n7005);
   U1981 : OAI22_X1 port map( A1 => n13370, A2 => n13266, B1 => n13361, B2 => 
                           n14454, ZN => n7006);
   U1982 : OAI22_X1 port map( A1 => n13370, A2 => n13269, B1 => n13361, B2 => 
                           n14453, ZN => n7007);
   U1983 : OAI22_X1 port map( A1 => n13369, A2 => n13272, B1 => n13361, B2 => 
                           n14452, ZN => n7008);
   U1984 : OAI22_X1 port map( A1 => n13369, A2 => n13275, B1 => n13361, B2 => 
                           n14451, ZN => n7009);
   U1985 : OAI22_X1 port map( A1 => n13369, A2 => n13278, B1 => n13362, B2 => 
                           n14450, ZN => n7010);
   U1986 : OAI22_X1 port map( A1 => n13369, A2 => n13281, B1 => n13362, B2 => 
                           n14449, ZN => n7011);
   U1987 : OAI22_X1 port map( A1 => n13369, A2 => n13284, B1 => n13362, B2 => 
                           n14448, ZN => n7012);
   U1988 : OAI22_X1 port map( A1 => n13368, A2 => n13287, B1 => n13362, B2 => 
                           n14447, ZN => n7013);
   U1989 : OAI22_X1 port map( A1 => n13368, A2 => n13290, B1 => n13362, B2 => 
                           n14446, ZN => n7014);
   U1990 : OAI22_X1 port map( A1 => n13368, A2 => n13293, B1 => n13362, B2 => 
                           n14445, ZN => n7015);
   U1991 : OAI22_X1 port map( A1 => n13368, A2 => n13296, B1 => n13362, B2 => 
                           n14444, ZN => n7016);
   U1992 : OAI22_X1 port map( A1 => n13368, A2 => n13299, B1 => n13362, B2 => 
                           n14443, ZN => n7017);
   U1993 : OAI22_X1 port map( A1 => n13367, A2 => n13302, B1 => n13362, B2 => 
                           n14442, ZN => n7018);
   U1994 : OAI22_X1 port map( A1 => n13367, A2 => n13305, B1 => n13362, B2 => 
                           n14441, ZN => n7019);
   U1995 : OAI22_X1 port map( A1 => n13365, A2 => n13335, B1 => n13363, B2 => 
                           n14440, ZN => n7029);
   U1996 : OAI22_X1 port map( A1 => n13365, A2 => n13338, B1 => n13363, B2 => 
                           n14439, ZN => n7030);
   U1997 : OAI22_X1 port map( A1 => n13365, A2 => n13341, B1 => n13363, B2 => 
                           n14438, ZN => n7031);
   U1998 : OAI22_X1 port map( A1 => n13365, A2 => n13344, B1 => n13363, B2 => 
                           n14437, ZN => n7032);
   U1999 : OAI22_X1 port map( A1 => n13364, A2 => n13347, B1 => n13363, B2 => 
                           n14436, ZN => n7033);
   U2000 : OAI22_X1 port map( A1 => n13159, A2 => n13290, B1 => n13153, B2 => 
                           n14432, ZN => n6950);
   U2001 : OAI22_X1 port map( A1 => n13159, A2 => n13293, B1 => n13153, B2 => 
                           n14431, ZN => n6951);
   U2002 : OAI22_X1 port map( A1 => n13159, A2 => n13296, B1 => n13153, B2 => 
                           n14430, ZN => n6952);
   U2003 : OAI22_X1 port map( A1 => n13159, A2 => n13299, B1 => n13153, B2 => 
                           n14429, ZN => n6953);
   U2004 : OAI22_X1 port map( A1 => n13158, A2 => n13302, B1 => n13153, B2 => 
                           n14428, ZN => n6954);
   U2005 : OAI22_X1 port map( A1 => n13158, A2 => n13305, B1 => n13153, B2 => 
                           n14427, ZN => n6955);
   U2006 : OAI22_X1 port map( A1 => n13158, A2 => n13308, B1 => n13153, B2 => 
                           n14426, ZN => n6956);
   U2007 : OAI22_X1 port map( A1 => n13158, A2 => n13311, B1 => n13153, B2 => 
                           n14425, ZN => n6957);
   U2008 : OAI22_X1 port map( A1 => n13158, A2 => n13314, B1 => n13154, B2 => 
                           n14424, ZN => n6958);
   U2009 : OAI22_X1 port map( A1 => n13157, A2 => n13317, B1 => n13154, B2 => 
                           n14423, ZN => n6959);
   U2010 : OAI22_X1 port map( A1 => n13157, A2 => n13320, B1 => n13154, B2 => 
                           n14422, ZN => n6960);
   U2011 : OAI22_X1 port map( A1 => n13157, A2 => n13323, B1 => n13154, B2 => 
                           n14421, ZN => n6961);
   U2012 : OAI22_X1 port map( A1 => n13157, A2 => n13326, B1 => n13154, B2 => 
                           n14420, ZN => n6962);
   U2013 : OAI22_X1 port map( A1 => n13157, A2 => n13329, B1 => n13154, B2 => 
                           n14419, ZN => n6963);
   U2014 : OAI22_X1 port map( A1 => n13156, A2 => n13332, B1 => n13154, B2 => 
                           n14418, ZN => n6964);
   U2015 : OAI22_X1 port map( A1 => n13156, A2 => n13335, B1 => n13154, B2 => 
                           n14417, ZN => n6965);
   U2016 : OAI22_X1 port map( A1 => n13156, A2 => n13338, B1 => n13154, B2 => 
                           n14416, ZN => n6966);
   U2017 : OAI22_X1 port map( A1 => n13156, A2 => n13341, B1 => n13154, B2 => 
                           n14415, ZN => n6967);
   U2018 : OAI22_X1 port map( A1 => n13156, A2 => n13344, B1 => n13154, B2 => 
                           n14414, ZN => n6968);
   U2019 : OAI22_X1 port map( A1 => n13155, A2 => n13347, B1 => n13154, B2 => 
                           n14413, ZN => n6969);
   U2020 : OAI22_X1 port map( A1 => n13161, A2 => n13257, B1 => n13152, B2 => 
                           n14322, ZN => n6939);
   U2021 : OAI22_X1 port map( A1 => n13161, A2 => n13260, B1 => n13152, B2 => 
                           n14321, ZN => n6940);
   U2022 : OAI22_X1 port map( A1 => n13161, A2 => n13263, B1 => n13152, B2 => 
                           n14320, ZN => n6941);
   U2023 : OAI22_X1 port map( A1 => n13161, A2 => n13266, B1 => n13152, B2 => 
                           n14319, ZN => n6942);
   U2024 : OAI22_X1 port map( A1 => n13161, A2 => n13269, B1 => n13152, B2 => 
                           n14318, ZN => n6943);
   U2025 : OAI22_X1 port map( A1 => n13160, A2 => n13272, B1 => n13152, B2 => 
                           n14317, ZN => n6944);
   U2026 : OAI22_X1 port map( A1 => n13160, A2 => n13275, B1 => n13152, B2 => 
                           n14316, ZN => n6945);
   U2027 : OAI22_X1 port map( A1 => n13160, A2 => n13278, B1 => n13153, B2 => 
                           n14315, ZN => n6946);
   U2028 : OAI22_X1 port map( A1 => n13160, A2 => n13281, B1 => n13153, B2 => 
                           n14314, ZN => n6947);
   U2029 : OAI22_X1 port map( A1 => n13160, A2 => n13284, B1 => n13153, B2 => 
                           n14313, ZN => n6948);
   U2030 : OAI22_X1 port map( A1 => n13159, A2 => n13287, B1 => n13153, B2 => 
                           n14312, ZN => n6949);
   U2031 : OAI22_X1 port map( A1 => n13371, A2 => n13242, B1 => n13361, B2 => 
                           n14294, ZN => n6998);
   U2032 : OAI22_X1 port map( A1 => n13371, A2 => n13245, B1 => n13361, B2 => 
                           n14293, ZN => n6999);
   U2033 : OAI22_X1 port map( A1 => n13371, A2 => n13248, B1 => n13361, B2 => 
                           n14292, ZN => n7000);
   U2034 : OAI22_X1 port map( A1 => n13371, A2 => n13251, B1 => n13361, B2 => 
                           n14291, ZN => n7001);
   U2035 : OAI22_X1 port map( A1 => n13371, A2 => n13254, B1 => n13361, B2 => 
                           n14290, ZN => n7002);
   U2036 : OAI22_X1 port map( A1 => n13370, A2 => n13257, B1 => n13361, B2 => 
                           n14289, ZN => n7003);
   U2037 : OAI22_X1 port map( A1 => n13102, A2 => n13242, B1 => n13092, B2 => 
                           n14288, ZN => n6742);
   U2038 : OAI22_X1 port map( A1 => n13102, A2 => n13245, B1 => n13092, B2 => 
                           n14287, ZN => n6743);
   U2039 : OAI22_X1 port map( A1 => n13102, A2 => n13248, B1 => n13092, B2 => 
                           n14286, ZN => n6744);
   U2040 : OAI22_X1 port map( A1 => n13102, A2 => n13251, B1 => n13092, B2 => 
                           n14285, ZN => n6745);
   U2041 : OAI22_X1 port map( A1 => n13102, A2 => n13254, B1 => n13092, B2 => 
                           n14284, ZN => n6746);
   U2042 : OAI22_X1 port map( A1 => n13101, A2 => n13257, B1 => n13092, B2 => 
                           n14283, ZN => n6747);
   U2043 : OAI22_X1 port map( A1 => n13101, A2 => n13260, B1 => n13092, B2 => 
                           n14282, ZN => n6748);
   U2044 : OAI22_X1 port map( A1 => n13101, A2 => n13263, B1 => n13092, B2 => 
                           n14281, ZN => n6749);
   U2045 : OAI22_X1 port map( A1 => n13101, A2 => n13266, B1 => n13092, B2 => 
                           n14280, ZN => n6750);
   U2046 : OAI22_X1 port map( A1 => n13101, A2 => n13269, B1 => n13092, B2 => 
                           n14279, ZN => n6751);
   U2047 : OAI22_X1 port map( A1 => n13100, A2 => n13272, B1 => n13092, B2 => 
                           n14278, ZN => n6752);
   U2048 : OAI22_X1 port map( A1 => n13100, A2 => n13275, B1 => n13092, B2 => 
                           n14277, ZN => n6753);
   U2049 : OAI22_X1 port map( A1 => n13100, A2 => n13278, B1 => n13093, B2 => 
                           n14276, ZN => n6754);
   U2050 : OAI22_X1 port map( A1 => n13100, A2 => n13281, B1 => n13093, B2 => 
                           n14275, ZN => n6755);
   U2051 : OAI22_X1 port map( A1 => n13100, A2 => n13284, B1 => n13093, B2 => 
                           n14274, ZN => n6756);
   U2052 : OAI22_X1 port map( A1 => n13099, A2 => n13287, B1 => n13093, B2 => 
                           n14273, ZN => n6757);
   U2053 : OAI22_X1 port map( A1 => n13099, A2 => n13290, B1 => n13093, B2 => 
                           n14272, ZN => n6758);
   U2054 : OAI22_X1 port map( A1 => n13099, A2 => n13293, B1 => n13093, B2 => 
                           n14271, ZN => n6759);
   U2055 : OAI22_X1 port map( A1 => n13099, A2 => n13296, B1 => n13093, B2 => 
                           n14270, ZN => n6760);
   U2056 : OAI22_X1 port map( A1 => n13099, A2 => n13299, B1 => n13093, B2 => 
                           n14269, ZN => n6761);
   U2057 : OAI22_X1 port map( A1 => n13098, A2 => n13302, B1 => n13093, B2 => 
                           n14268, ZN => n6762);
   U2058 : OAI22_X1 port map( A1 => n13098, A2 => n13305, B1 => n13093, B2 => 
                           n14267, ZN => n6763);
   U2059 : OAI22_X1 port map( A1 => n13098, A2 => n13308, B1 => n13093, B2 => 
                           n14266, ZN => n6764);
   U2060 : OAI22_X1 port map( A1 => n13098, A2 => n13311, B1 => n13093, B2 => 
                           n14265, ZN => n6765);
   U2061 : OAI22_X1 port map( A1 => n13098, A2 => n13314, B1 => n13094, B2 => 
                           n14264, ZN => n6766);
   U2062 : OAI22_X1 port map( A1 => n13097, A2 => n13317, B1 => n13094, B2 => 
                           n14263, ZN => n6767);
   U2063 : OAI22_X1 port map( A1 => n13097, A2 => n13320, B1 => n13094, B2 => 
                           n14262, ZN => n6768);
   U2064 : OAI22_X1 port map( A1 => n13097, A2 => n13323, B1 => n13094, B2 => 
                           n14261, ZN => n6769);
   U2065 : OAI22_X1 port map( A1 => n13097, A2 => n13326, B1 => n13094, B2 => 
                           n14260, ZN => n6770);
   U2066 : OAI22_X1 port map( A1 => n13097, A2 => n13329, B1 => n13094, B2 => 
                           n14259, ZN => n6771);
   U2067 : OAI22_X1 port map( A1 => n13096, A2 => n13332, B1 => n13094, B2 => 
                           n14258, ZN => n6772);
   U2068 : OAI22_X1 port map( A1 => n13096, A2 => n13335, B1 => n13094, B2 => 
                           n14257, ZN => n6773);
   U2069 : OAI22_X1 port map( A1 => n13096, A2 => n13338, B1 => n13094, B2 => 
                           n14256, ZN => n6774);
   U2070 : OAI22_X1 port map( A1 => n13096, A2 => n13341, B1 => n13094, B2 => 
                           n14255, ZN => n6775);
   U2071 : OAI22_X1 port map( A1 => n13096, A2 => n13344, B1 => n13094, B2 => 
                           n14254, ZN => n6776);
   U2072 : OAI22_X1 port map( A1 => n13095, A2 => n13347, B1 => n13094, B2 => 
                           n14253, ZN => n6777);
   U2073 : OAI22_X1 port map( A1 => n13082, A2 => n13242, B1 => n13072, B2 => 
                           n14252, ZN => n6678);
   U2074 : OAI22_X1 port map( A1 => n13082, A2 => n13245, B1 => n13072, B2 => 
                           n14251, ZN => n6679);
   U2075 : OAI22_X1 port map( A1 => n13082, A2 => n13248, B1 => n13072, B2 => 
                           n14250, ZN => n6680);
   U2076 : OAI22_X1 port map( A1 => n13082, A2 => n13251, B1 => n13072, B2 => 
                           n14249, ZN => n6681);
   U2077 : OAI22_X1 port map( A1 => n13082, A2 => n13254, B1 => n13072, B2 => 
                           n14248, ZN => n6682);
   U2078 : OAI22_X1 port map( A1 => n13081, A2 => n13257, B1 => n13072, B2 => 
                           n14247, ZN => n6683);
   U2079 : OAI22_X1 port map( A1 => n13081, A2 => n13260, B1 => n13072, B2 => 
                           n14246, ZN => n6684);
   U2080 : OAI22_X1 port map( A1 => n13081, A2 => n13263, B1 => n13072, B2 => 
                           n14245, ZN => n6685);
   U2081 : OAI22_X1 port map( A1 => n13081, A2 => n13266, B1 => n13072, B2 => 
                           n14244, ZN => n6686);
   U2082 : OAI22_X1 port map( A1 => n13081, A2 => n13269, B1 => n13072, B2 => 
                           n14243, ZN => n6687);
   U2083 : OAI22_X1 port map( A1 => n13080, A2 => n13272, B1 => n13072, B2 => 
                           n14242, ZN => n6688);
   U2084 : OAI22_X1 port map( A1 => n13080, A2 => n13275, B1 => n13072, B2 => 
                           n14241, ZN => n6689);
   U2085 : OAI22_X1 port map( A1 => n13080, A2 => n13278, B1 => n13073, B2 => 
                           n14240, ZN => n6690);
   U2086 : OAI22_X1 port map( A1 => n13080, A2 => n13281, B1 => n13073, B2 => 
                           n14239, ZN => n6691);
   U2087 : OAI22_X1 port map( A1 => n13080, A2 => n13284, B1 => n13073, B2 => 
                           n14238, ZN => n6692);
   U2088 : OAI22_X1 port map( A1 => n13079, A2 => n13287, B1 => n13073, B2 => 
                           n14237, ZN => n6693);
   U2089 : OAI22_X1 port map( A1 => n13079, A2 => n13290, B1 => n13073, B2 => 
                           n14236, ZN => n6694);
   U2090 : OAI22_X1 port map( A1 => n13079, A2 => n13293, B1 => n13073, B2 => 
                           n14235, ZN => n6695);
   U2091 : OAI22_X1 port map( A1 => n13079, A2 => n13296, B1 => n13073, B2 => 
                           n14234, ZN => n6696);
   U2092 : OAI22_X1 port map( A1 => n13079, A2 => n13299, B1 => n13073, B2 => 
                           n14233, ZN => n6697);
   U2093 : OAI22_X1 port map( A1 => n13078, A2 => n13302, B1 => n13073, B2 => 
                           n14232, ZN => n6698);
   U2094 : OAI22_X1 port map( A1 => n13078, A2 => n13305, B1 => n13073, B2 => 
                           n14231, ZN => n6699);
   U2095 : OAI22_X1 port map( A1 => n13078, A2 => n13308, B1 => n13073, B2 => 
                           n14230, ZN => n6700);
   U2096 : OAI22_X1 port map( A1 => n13078, A2 => n13311, B1 => n13073, B2 => 
                           n14229, ZN => n6701);
   U2097 : OAI22_X1 port map( A1 => n13078, A2 => n13314, B1 => n13074, B2 => 
                           n14228, ZN => n6702);
   U2098 : OAI22_X1 port map( A1 => n13077, A2 => n13317, B1 => n13074, B2 => 
                           n14227, ZN => n6703);
   U2099 : OAI22_X1 port map( A1 => n13077, A2 => n13320, B1 => n13074, B2 => 
                           n14226, ZN => n6704);
   U2100 : OAI22_X1 port map( A1 => n13077, A2 => n13323, B1 => n13074, B2 => 
                           n14225, ZN => n6705);
   U2101 : OAI22_X1 port map( A1 => n13077, A2 => n13326, B1 => n13074, B2 => 
                           n14224, ZN => n6706);
   U2102 : OAI22_X1 port map( A1 => n13077, A2 => n13329, B1 => n13074, B2 => 
                           n14223, ZN => n6707);
   U2103 : OAI22_X1 port map( A1 => n13076, A2 => n13332, B1 => n13074, B2 => 
                           n14222, ZN => n6708);
   U2104 : OAI22_X1 port map( A1 => n13076, A2 => n13335, B1 => n13074, B2 => 
                           n14221, ZN => n6709);
   U2105 : OAI22_X1 port map( A1 => n13076, A2 => n13338, B1 => n13074, B2 => 
                           n14220, ZN => n6710);
   U2106 : OAI22_X1 port map( A1 => n13076, A2 => n13341, B1 => n13074, B2 => 
                           n14219, ZN => n6711);
   U2107 : OAI22_X1 port map( A1 => n13076, A2 => n13344, B1 => n13074, B2 => 
                           n14218, ZN => n6712);
   U2108 : OAI22_X1 port map( A1 => n13075, A2 => n13347, B1 => n13074, B2 => 
                           n14217, ZN => n6713);
   U2109 : OAI22_X1 port map( A1 => n12604, A2 => n13292, B1 => n12598, B2 => 
                           n14106, ZN => n5158);
   U2110 : OAI22_X1 port map( A1 => n12604, A2 => n13295, B1 => n12598, B2 => 
                           n14105, ZN => n5159);
   U2111 : OAI22_X1 port map( A1 => n12604, A2 => n13298, B1 => n12598, B2 => 
                           n14104, ZN => n5160);
   U2112 : OAI22_X1 port map( A1 => n12604, A2 => n13301, B1 => n12598, B2 => 
                           n14103, ZN => n5161);
   U2113 : OAI22_X1 port map( A1 => n12603, A2 => n13304, B1 => n12598, B2 => 
                           n14102, ZN => n5162);
   U2114 : OAI22_X1 port map( A1 => n12603, A2 => n13307, B1 => n12598, B2 => 
                           n14101, ZN => n5163);
   U2115 : OAI22_X1 port map( A1 => n12603, A2 => n13310, B1 => n12598, B2 => 
                           n14100, ZN => n5164);
   U2116 : OAI22_X1 port map( A1 => n12603, A2 => n13313, B1 => n12598, B2 => 
                           n14099, ZN => n5165);
   U2117 : OAI22_X1 port map( A1 => n12603, A2 => n13316, B1 => n12599, B2 => 
                           n14098, ZN => n5166);
   U2118 : OAI22_X1 port map( A1 => n12602, A2 => n13319, B1 => n12599, B2 => 
                           n14097, ZN => n5167);
   U2119 : OAI22_X1 port map( A1 => n12602, A2 => n13322, B1 => n12599, B2 => 
                           n14096, ZN => n5168);
   U2120 : OAI22_X1 port map( A1 => n12602, A2 => n13325, B1 => n12599, B2 => 
                           n14095, ZN => n5169);
   U2121 : OAI22_X1 port map( A1 => n12602, A2 => n13328, B1 => n12599, B2 => 
                           n14094, ZN => n5170);
   U2122 : OAI22_X1 port map( A1 => n12602, A2 => n13331, B1 => n12599, B2 => 
                           n14093, ZN => n5171);
   U2123 : OAI22_X1 port map( A1 => n12601, A2 => n13334, B1 => n12599, B2 => 
                           n14092, ZN => n5172);
   U2124 : OAI22_X1 port map( A1 => n12601, A2 => n13337, B1 => n12599, B2 => 
                           n14091, ZN => n5173);
   U2125 : OAI22_X1 port map( A1 => n12601, A2 => n13340, B1 => n12599, B2 => 
                           n14090, ZN => n5174);
   U2126 : OAI22_X1 port map( A1 => n12601, A2 => n13343, B1 => n12599, B2 => 
                           n14089, ZN => n5175);
   U2127 : OAI22_X1 port map( A1 => n12601, A2 => n13346, B1 => n12599, B2 => 
                           n14088, ZN => n5176);
   U2128 : OAI22_X1 port map( A1 => n12600, A2 => n13349, B1 => n12599, B2 => 
                           n14087, ZN => n5177);
   U2129 : OAI22_X1 port map( A1 => n12683, A2 => n13256, B1 => n12673, B2 => 
                           n14059, ZN => n5402);
   U2130 : OAI22_X1 port map( A1 => n12682, A2 => n13259, B1 => n12673, B2 => 
                           n14058, ZN => n5403);
   U2131 : OAI22_X1 port map( A1 => n12682, A2 => n13262, B1 => n12673, B2 => 
                           n14057, ZN => n5404);
   U2132 : OAI22_X1 port map( A1 => n12682, A2 => n13265, B1 => n12673, B2 => 
                           n14056, ZN => n5405);
   U2133 : OAI22_X1 port map( A1 => n12682, A2 => n13268, B1 => n12673, B2 => 
                           n14055, ZN => n5406);
   U2134 : OAI22_X1 port map( A1 => n12682, A2 => n13271, B1 => n12673, B2 => 
                           n14054, ZN => n5407);
   U2135 : OAI22_X1 port map( A1 => n12681, A2 => n13274, B1 => n12673, B2 => 
                           n14053, ZN => n5408);
   U2136 : OAI22_X1 port map( A1 => n12681, A2 => n13277, B1 => n12673, B2 => 
                           n14052, ZN => n5409);
   U2137 : OAI22_X1 port map( A1 => n12681, A2 => n13280, B1 => n12674, B2 => 
                           n14051, ZN => n5410);
   U2138 : OAI22_X1 port map( A1 => n12681, A2 => n13283, B1 => n12674, B2 => 
                           n14050, ZN => n5411);
   U2139 : OAI22_X1 port map( A1 => n12681, A2 => n13286, B1 => n12674, B2 => 
                           n14049, ZN => n5412);
   U2140 : OAI22_X1 port map( A1 => n12680, A2 => n13289, B1 => n12674, B2 => 
                           n14048, ZN => n5413);
   U2141 : OAI22_X1 port map( A1 => n12680, A2 => n13292, B1 => n12674, B2 => 
                           n14047, ZN => n5414);
   U2142 : OAI22_X1 port map( A1 => n12680, A2 => n13295, B1 => n12674, B2 => 
                           n14046, ZN => n5415);
   U2143 : OAI22_X1 port map( A1 => n12680, A2 => n13298, B1 => n12674, B2 => 
                           n14045, ZN => n5416);
   U2144 : OAI22_X1 port map( A1 => n12680, A2 => n13301, B1 => n12674, B2 => 
                           n14044, ZN => n5417);
   U2145 : OAI22_X1 port map( A1 => n12679, A2 => n13304, B1 => n12674, B2 => 
                           n14043, ZN => n5418);
   U2146 : OAI22_X1 port map( A1 => n12679, A2 => n13307, B1 => n12674, B2 => 
                           n14042, ZN => n5419);
   U2147 : OAI22_X1 port map( A1 => n12679, A2 => n13310, B1 => n12674, B2 => 
                           n14041, ZN => n5420);
   U2148 : OAI22_X1 port map( A1 => n12679, A2 => n13313, B1 => n12674, B2 => 
                           n14040, ZN => n5421);
   U2149 : OAI22_X1 port map( A1 => n12679, A2 => n13316, B1 => n12675, B2 => 
                           n14039, ZN => n5422);
   U2150 : OAI22_X1 port map( A1 => n12678, A2 => n13319, B1 => n12675, B2 => 
                           n14038, ZN => n5423);
   U2151 : OAI22_X1 port map( A1 => n12678, A2 => n13322, B1 => n12675, B2 => 
                           n14037, ZN => n5424);
   U2152 : OAI22_X1 port map( A1 => n12678, A2 => n13325, B1 => n12675, B2 => 
                           n14036, ZN => n5425);
   U2153 : OAI22_X1 port map( A1 => n12607, A2 => n13244, B1 => n12597, B2 => 
                           n13944, ZN => n5142);
   U2154 : OAI22_X1 port map( A1 => n12607, A2 => n13247, B1 => n12597, B2 => 
                           n13943, ZN => n5143);
   U2155 : OAI22_X1 port map( A1 => n12607, A2 => n13250, B1 => n12597, B2 => 
                           n13942, ZN => n5144);
   U2156 : OAI22_X1 port map( A1 => n12607, A2 => n13253, B1 => n12597, B2 => 
                           n13941, ZN => n5145);
   U2157 : OAI22_X1 port map( A1 => n12607, A2 => n13256, B1 => n12597, B2 => 
                           n13940, ZN => n5146);
   U2158 : OAI22_X1 port map( A1 => n12606, A2 => n13259, B1 => n12597, B2 => 
                           n13939, ZN => n5147);
   U2159 : OAI22_X1 port map( A1 => n12606, A2 => n13262, B1 => n12597, B2 => 
                           n13938, ZN => n5148);
   U2160 : OAI22_X1 port map( A1 => n12606, A2 => n13265, B1 => n12597, B2 => 
                           n13937, ZN => n5149);
   U2161 : OAI22_X1 port map( A1 => n12606, A2 => n13268, B1 => n12597, B2 => 
                           n13936, ZN => n5150);
   U2162 : OAI22_X1 port map( A1 => n12606, A2 => n13271, B1 => n12597, B2 => 
                           n13935, ZN => n5151);
   U2163 : OAI22_X1 port map( A1 => n12605, A2 => n13274, B1 => n12597, B2 => 
                           n13934, ZN => n5152);
   U2164 : OAI22_X1 port map( A1 => n12605, A2 => n13277, B1 => n12597, B2 => 
                           n13933, ZN => n5153);
   U2165 : OAI22_X1 port map( A1 => n12605, A2 => n13280, B1 => n12598, B2 => 
                           n13932, ZN => n5154);
   U2166 : OAI22_X1 port map( A1 => n12605, A2 => n13283, B1 => n12598, B2 => 
                           n13931, ZN => n5155);
   U2167 : OAI22_X1 port map( A1 => n12605, A2 => n13286, B1 => n12598, B2 => 
                           n13930, ZN => n5156);
   U2168 : OAI22_X1 port map( A1 => n12604, A2 => n13289, B1 => n12598, B2 => 
                           n13929, ZN => n5157);
   U2169 : OAI22_X1 port map( A1 => n12683, A2 => n13244, B1 => n12673, B2 => 
                           n13872, ZN => n5398);
   U2170 : OAI22_X1 port map( A1 => n12683, A2 => n13247, B1 => n12673, B2 => 
                           n13871, ZN => n5399);
   U2171 : OAI22_X1 port map( A1 => n12683, A2 => n13250, B1 => n12673, B2 => 
                           n13870, ZN => n5400);
   U2172 : OAI22_X1 port map( A1 => n12683, A2 => n13253, B1 => n12673, B2 => 
                           n13869, ZN => n5401);
   U2173 : OAI22_X1 port map( A1 => n12626, A2 => n13244, B1 => n12616, B2 => 
                           n13786, ZN => n5206);
   U2174 : OAI22_X1 port map( A1 => n12626, A2 => n13247, B1 => n12616, B2 => 
                           n13785, ZN => n5207);
   U2175 : OAI22_X1 port map( A1 => n12626, A2 => n13250, B1 => n12616, B2 => 
                           n13784, ZN => n5208);
   U2176 : OAI22_X1 port map( A1 => n12626, A2 => n13253, B1 => n12616, B2 => 
                           n13783, ZN => n5209);
   U2177 : OAI22_X1 port map( A1 => n12626, A2 => n13256, B1 => n12616, B2 => 
                           n13782, ZN => n5210);
   U2178 : OAI22_X1 port map( A1 => n12625, A2 => n13259, B1 => n12616, B2 => 
                           n13781, ZN => n5211);
   U2179 : OAI22_X1 port map( A1 => n12625, A2 => n13262, B1 => n12616, B2 => 
                           n13780, ZN => n5212);
   U2180 : OAI22_X1 port map( A1 => n12625, A2 => n13265, B1 => n12616, B2 => 
                           n13779, ZN => n5213);
   U2181 : OAI22_X1 port map( A1 => n12625, A2 => n13268, B1 => n12616, B2 => 
                           n13778, ZN => n5214);
   U2182 : OAI22_X1 port map( A1 => n12625, A2 => n13271, B1 => n12616, B2 => 
                           n13777, ZN => n5215);
   U2183 : OAI22_X1 port map( A1 => n12624, A2 => n13274, B1 => n12616, B2 => 
                           n13776, ZN => n5216);
   U2184 : OAI22_X1 port map( A1 => n12624, A2 => n13277, B1 => n12616, B2 => 
                           n13775, ZN => n5217);
   U2185 : OAI22_X1 port map( A1 => n12624, A2 => n13280, B1 => n12617, B2 => 
                           n13774, ZN => n5218);
   U2186 : OAI22_X1 port map( A1 => n12624, A2 => n13283, B1 => n12617, B2 => 
                           n13773, ZN => n5219);
   U2187 : OAI22_X1 port map( A1 => n12624, A2 => n13286, B1 => n12617, B2 => 
                           n13772, ZN => n5220);
   U2188 : OAI22_X1 port map( A1 => n12623, A2 => n13289, B1 => n12617, B2 => 
                           n13771, ZN => n5221);
   U2189 : OAI22_X1 port map( A1 => n12623, A2 => n13292, B1 => n12617, B2 => 
                           n13770, ZN => n5222);
   U2190 : OAI22_X1 port map( A1 => n12623, A2 => n13295, B1 => n12617, B2 => 
                           n13769, ZN => n5223);
   U2191 : OAI22_X1 port map( A1 => n12623, A2 => n13298, B1 => n12617, B2 => 
                           n13768, ZN => n5224);
   U2192 : OAI22_X1 port map( A1 => n12623, A2 => n13301, B1 => n12617, B2 => 
                           n13767, ZN => n5225);
   U2193 : OAI22_X1 port map( A1 => n12622, A2 => n13304, B1 => n12617, B2 => 
                           n13766, ZN => n5226);
   U2194 : OAI22_X1 port map( A1 => n12622, A2 => n13307, B1 => n12617, B2 => 
                           n13765, ZN => n5227);
   U2195 : OAI22_X1 port map( A1 => n12622, A2 => n13310, B1 => n12617, B2 => 
                           n13764, ZN => n5228);
   U2196 : OAI22_X1 port map( A1 => n12622, A2 => n13313, B1 => n12617, B2 => 
                           n13763, ZN => n5229);
   U2197 : OAI22_X1 port map( A1 => n12622, A2 => n13316, B1 => n12618, B2 => 
                           n13762, ZN => n5230);
   U2198 : OAI22_X1 port map( A1 => n12621, A2 => n13319, B1 => n12618, B2 => 
                           n13761, ZN => n5231);
   U2199 : OAI22_X1 port map( A1 => n12621, A2 => n13322, B1 => n12618, B2 => 
                           n13760, ZN => n5232);
   U2200 : OAI22_X1 port map( A1 => n12621, A2 => n13325, B1 => n12618, B2 => 
                           n13759, ZN => n5233);
   U2201 : OAI22_X1 port map( A1 => n12621, A2 => n13328, B1 => n12618, B2 => 
                           n13758, ZN => n5234);
   U2202 : OAI22_X1 port map( A1 => n12621, A2 => n13331, B1 => n12618, B2 => 
                           n13757, ZN => n5235);
   U2203 : OAI22_X1 port map( A1 => n12620, A2 => n13334, B1 => n12618, B2 => 
                           n13756, ZN => n5236);
   U2204 : OAI22_X1 port map( A1 => n12620, A2 => n13337, B1 => n12618, B2 => 
                           n13755, ZN => n5237);
   U2205 : OAI22_X1 port map( A1 => n12620, A2 => n13340, B1 => n12618, B2 => 
                           n13754, ZN => n5238);
   U2206 : OAI22_X1 port map( A1 => n12620, A2 => n13343, B1 => n12618, B2 => 
                           n13753, ZN => n5239);
   U2207 : OAI22_X1 port map( A1 => n12620, A2 => n13346, B1 => n12618, B2 => 
                           n13752, ZN => n5240);
   U2208 : OAI22_X1 port map( A1 => n12619, A2 => n13349, B1 => n12618, B2 => 
                           n13751, ZN => n5241);
   U2209 : OAI22_X1 port map( A1 => n12678, A2 => n13328, B1 => n12675, B2 => 
                           n13742, ZN => n5426);
   U2210 : OAI22_X1 port map( A1 => n12678, A2 => n13331, B1 => n12675, B2 => 
                           n13741, ZN => n5427);
   U2211 : OAI22_X1 port map( A1 => n12677, A2 => n13334, B1 => n12675, B2 => 
                           n13740, ZN => n5428);
   U2212 : OAI22_X1 port map( A1 => n12677, A2 => n13337, B1 => n12675, B2 => 
                           n13739, ZN => n5429);
   U2213 : OAI22_X1 port map( A1 => n12677, A2 => n13340, B1 => n12675, B2 => 
                           n13738, ZN => n5430);
   U2214 : OAI22_X1 port map( A1 => n12677, A2 => n13343, B1 => n12675, B2 => 
                           n13737, ZN => n5431);
   U2215 : OAI22_X1 port map( A1 => n12677, A2 => n13346, B1 => n12675, B2 => 
                           n13736, ZN => n5432);
   U2216 : OAI22_X1 port map( A1 => n12676, A2 => n13349, B1 => n12675, B2 => 
                           n13735, ZN => n5433);
   U2217 : OAI22_X1 port map( A1 => n12702, A2 => n13244, B1 => n12692, B2 => 
                           n13706, ZN => n5462);
   U2218 : OAI22_X1 port map( A1 => n12702, A2 => n13247, B1 => n12692, B2 => 
                           n13705, ZN => n5463);
   U2219 : OAI22_X1 port map( A1 => n12702, A2 => n13250, B1 => n12692, B2 => 
                           n13704, ZN => n5464);
   U2220 : OAI22_X1 port map( A1 => n12702, A2 => n13253, B1 => n12692, B2 => 
                           n13703, ZN => n5465);
   U2221 : OAI22_X1 port map( A1 => n12702, A2 => n13256, B1 => n12692, B2 => 
                           n13702, ZN => n5466);
   U2222 : OAI22_X1 port map( A1 => n12701, A2 => n13259, B1 => n12692, B2 => 
                           n13701, ZN => n5467);
   U2223 : OAI22_X1 port map( A1 => n12701, A2 => n13262, B1 => n12692, B2 => 
                           n13700, ZN => n5468);
   U2224 : OAI22_X1 port map( A1 => n12701, A2 => n13265, B1 => n12692, B2 => 
                           n13699, ZN => n5469);
   U2225 : OAI22_X1 port map( A1 => n12701, A2 => n13268, B1 => n12692, B2 => 
                           n13698, ZN => n5470);
   U2226 : OAI22_X1 port map( A1 => n12701, A2 => n13271, B1 => n12692, B2 => 
                           n13697, ZN => n5471);
   U2227 : OAI22_X1 port map( A1 => n12700, A2 => n13274, B1 => n12692, B2 => 
                           n13696, ZN => n5472);
   U2228 : OAI22_X1 port map( A1 => n12700, A2 => n13277, B1 => n12692, B2 => 
                           n13695, ZN => n5473);
   U2229 : OAI22_X1 port map( A1 => n12700, A2 => n13280, B1 => n12693, B2 => 
                           n13694, ZN => n5474);
   U2230 : OAI22_X1 port map( A1 => n12700, A2 => n13283, B1 => n12693, B2 => 
                           n13693, ZN => n5475);
   U2231 : OAI22_X1 port map( A1 => n12700, A2 => n13286, B1 => n12693, B2 => 
                           n13692, ZN => n5476);
   U2232 : OAI22_X1 port map( A1 => n12699, A2 => n13289, B1 => n12693, B2 => 
                           n13691, ZN => n5477);
   U2233 : OAI22_X1 port map( A1 => n12699, A2 => n13292, B1 => n12693, B2 => 
                           n13690, ZN => n5478);
   U2234 : OAI22_X1 port map( A1 => n12699, A2 => n13295, B1 => n12693, B2 => 
                           n13689, ZN => n5479);
   U2235 : OAI22_X1 port map( A1 => n12699, A2 => n13298, B1 => n12693, B2 => 
                           n13688, ZN => n5480);
   U2236 : OAI22_X1 port map( A1 => n12699, A2 => n13301, B1 => n12693, B2 => 
                           n13687, ZN => n5481);
   U2237 : OAI22_X1 port map( A1 => n12698, A2 => n13304, B1 => n12693, B2 => 
                           n13686, ZN => n5482);
   U2238 : OAI22_X1 port map( A1 => n12698, A2 => n13307, B1 => n12693, B2 => 
                           n13685, ZN => n5483);
   U2239 : OAI22_X1 port map( A1 => n12698, A2 => n13310, B1 => n12693, B2 => 
                           n13684, ZN => n5484);
   U2240 : OAI22_X1 port map( A1 => n12698, A2 => n13313, B1 => n12693, B2 => 
                           n13683, ZN => n5485);
   U2241 : OAI22_X1 port map( A1 => n12698, A2 => n13316, B1 => n12694, B2 => 
                           n13682, ZN => n5486);
   U2242 : OAI22_X1 port map( A1 => n12697, A2 => n13319, B1 => n12694, B2 => 
                           n13681, ZN => n5487);
   U2243 : OAI22_X1 port map( A1 => n12697, A2 => n13322, B1 => n12694, B2 => 
                           n13680, ZN => n5488);
   U2244 : OAI22_X1 port map( A1 => n12697, A2 => n13325, B1 => n12694, B2 => 
                           n13679, ZN => n5489);
   U2245 : OAI22_X1 port map( A1 => n12697, A2 => n13328, B1 => n12694, B2 => 
                           n13678, ZN => n5490);
   U2246 : OAI22_X1 port map( A1 => n12697, A2 => n13331, B1 => n12694, B2 => 
                           n13677, ZN => n5491);
   U2247 : OAI22_X1 port map( A1 => n12696, A2 => n13334, B1 => n12694, B2 => 
                           n13676, ZN => n5492);
   U2248 : OAI22_X1 port map( A1 => n12696, A2 => n13337, B1 => n12694, B2 => 
                           n13675, ZN => n5493);
   U2249 : OAI22_X1 port map( A1 => n12696, A2 => n13340, B1 => n12694, B2 => 
                           n13674, ZN => n5494);
   U2250 : OAI22_X1 port map( A1 => n12696, A2 => n13343, B1 => n12694, B2 => 
                           n13673, ZN => n5495);
   U2251 : OAI22_X1 port map( A1 => n12696, A2 => n13346, B1 => n12694, B2 => 
                           n13672, ZN => n5496);
   U2252 : OAI22_X1 port map( A1 => n12695, A2 => n13349, B1 => n12694, B2 => 
                           n13671, ZN => n5497);
   U2253 : OAI22_X1 port map( A1 => n12882, A2 => n13243, B1 => n12872, B2 => 
                           n13643, ZN => n6038);
   U2254 : OAI22_X1 port map( A1 => n12882, A2 => n13246, B1 => n12872, B2 => 
                           n13642, ZN => n6039);
   U2255 : OAI22_X1 port map( A1 => n12882, A2 => n13249, B1 => n12872, B2 => 
                           n13641, ZN => n6040);
   U2256 : OAI22_X1 port map( A1 => n12882, A2 => n13252, B1 => n12872, B2 => 
                           n13640, ZN => n6041);
   U2257 : OAI22_X1 port map( A1 => n12882, A2 => n13255, B1 => n12872, B2 => 
                           n13639, ZN => n6042);
   U2258 : OAI22_X1 port map( A1 => n12881, A2 => n13258, B1 => n12872, B2 => 
                           n13638, ZN => n6043);
   U2259 : OAI22_X1 port map( A1 => n12881, A2 => n13261, B1 => n12872, B2 => 
                           n13637, ZN => n6044);
   U2260 : OAI22_X1 port map( A1 => n12881, A2 => n13264, B1 => n12872, B2 => 
                           n13636, ZN => n6045);
   U2261 : OAI22_X1 port map( A1 => n12881, A2 => n13267, B1 => n12872, B2 => 
                           n13635, ZN => n6046);
   U2262 : OAI22_X1 port map( A1 => n12881, A2 => n13270, B1 => n12872, B2 => 
                           n13634, ZN => n6047);
   U2263 : OAI22_X1 port map( A1 => n12880, A2 => n13273, B1 => n12872, B2 => 
                           n13633, ZN => n6048);
   U2264 : OAI22_X1 port map( A1 => n12880, A2 => n13276, B1 => n12872, B2 => 
                           n13632, ZN => n6049);
   U2265 : OAI22_X1 port map( A1 => n12880, A2 => n13279, B1 => n12873, B2 => 
                           n13631, ZN => n6050);
   U2266 : OAI22_X1 port map( A1 => n12880, A2 => n13282, B1 => n12873, B2 => 
                           n13630, ZN => n6051);
   U2267 : OAI22_X1 port map( A1 => n12880, A2 => n13285, B1 => n12873, B2 => 
                           n13629, ZN => n6052);
   U2268 : OAI22_X1 port map( A1 => n12879, A2 => n13288, B1 => n12873, B2 => 
                           n13628, ZN => n6053);
   U2269 : OAI22_X1 port map( A1 => n12879, A2 => n13291, B1 => n12873, B2 => 
                           n13627, ZN => n6054);
   U2270 : OAI22_X1 port map( A1 => n12879, A2 => n13294, B1 => n12873, B2 => 
                           n13626, ZN => n6055);
   U2271 : OAI22_X1 port map( A1 => n12879, A2 => n13297, B1 => n12873, B2 => 
                           n13625, ZN => n6056);
   U2272 : OAI22_X1 port map( A1 => n12879, A2 => n13300, B1 => n12873, B2 => 
                           n13624, ZN => n6057);
   U2273 : OAI22_X1 port map( A1 => n12878, A2 => n13303, B1 => n12873, B2 => 
                           n13623, ZN => n6058);
   U2274 : OAI22_X1 port map( A1 => n12878, A2 => n13306, B1 => n12873, B2 => 
                           n13622, ZN => n6059);
   U2275 : OAI22_X1 port map( A1 => n12878, A2 => n13309, B1 => n12873, B2 => 
                           n13621, ZN => n6060);
   U2276 : OAI22_X1 port map( A1 => n12878, A2 => n13312, B1 => n12873, B2 => 
                           n13620, ZN => n6061);
   U2277 : OAI22_X1 port map( A1 => n12878, A2 => n13315, B1 => n12874, B2 => 
                           n13619, ZN => n6062);
   U2278 : OAI22_X1 port map( A1 => n12877, A2 => n13318, B1 => n12874, B2 => 
                           n13618, ZN => n6063);
   U2279 : OAI22_X1 port map( A1 => n12877, A2 => n13321, B1 => n12874, B2 => 
                           n13617, ZN => n6064);
   U2280 : OAI22_X1 port map( A1 => n12877, A2 => n13324, B1 => n12874, B2 => 
                           n13616, ZN => n6065);
   U2281 : OAI22_X1 port map( A1 => n12877, A2 => n13327, B1 => n12874, B2 => 
                           n13615, ZN => n6066);
   U2282 : OAI22_X1 port map( A1 => n12877, A2 => n13330, B1 => n12874, B2 => 
                           n13614, ZN => n6067);
   U2283 : OAI22_X1 port map( A1 => n12876, A2 => n13333, B1 => n12874, B2 => 
                           n13613, ZN => n6068);
   U2284 : OAI22_X1 port map( A1 => n12876, A2 => n13336, B1 => n12874, B2 => 
                           n13612, ZN => n6069);
   U2285 : OAI22_X1 port map( A1 => n12876, A2 => n13339, B1 => n12874, B2 => 
                           n13611, ZN => n6070);
   U2286 : OAI22_X1 port map( A1 => n12876, A2 => n13342, B1 => n12874, B2 => 
                           n13610, ZN => n6071);
   U2287 : OAI22_X1 port map( A1 => n12876, A2 => n13345, B1 => n12874, B2 => 
                           n13609, ZN => n6072);
   U2288 : OAI22_X1 port map( A1 => n12875, A2 => n13348, B1 => n12874, B2 => 
                           n13608, ZN => n6073);
   U2289 : OAI22_X1 port map( A1 => n12902, A2 => n13243, B1 => n12892, B2 => 
                           n13579, ZN => n6102);
   U2290 : OAI22_X1 port map( A1 => n12902, A2 => n13246, B1 => n12892, B2 => 
                           n13578, ZN => n6103);
   U2291 : OAI22_X1 port map( A1 => n12902, A2 => n13249, B1 => n12892, B2 => 
                           n13577, ZN => n6104);
   U2292 : OAI22_X1 port map( A1 => n12902, A2 => n13252, B1 => n12892, B2 => 
                           n13576, ZN => n6105);
   U2293 : OAI22_X1 port map( A1 => n12902, A2 => n13255, B1 => n12892, B2 => 
                           n13575, ZN => n6106);
   U2294 : OAI22_X1 port map( A1 => n12901, A2 => n13258, B1 => n12892, B2 => 
                           n13574, ZN => n6107);
   U2295 : OAI22_X1 port map( A1 => n12901, A2 => n13261, B1 => n12892, B2 => 
                           n13573, ZN => n6108);
   U2296 : OAI22_X1 port map( A1 => n12901, A2 => n13264, B1 => n12892, B2 => 
                           n13572, ZN => n6109);
   U2297 : OAI22_X1 port map( A1 => n12901, A2 => n13267, B1 => n12892, B2 => 
                           n13571, ZN => n6110);
   U2298 : OAI22_X1 port map( A1 => n12901, A2 => n13270, B1 => n12892, B2 => 
                           n13570, ZN => n6111);
   U2299 : OAI22_X1 port map( A1 => n12900, A2 => n13273, B1 => n12892, B2 => 
                           n13569, ZN => n6112);
   U2300 : OAI22_X1 port map( A1 => n12900, A2 => n13276, B1 => n12892, B2 => 
                           n13568, ZN => n6113);
   U2301 : OAI22_X1 port map( A1 => n12900, A2 => n13279, B1 => n12893, B2 => 
                           n13567, ZN => n6114);
   U2302 : OAI22_X1 port map( A1 => n12900, A2 => n13282, B1 => n12893, B2 => 
                           n13566, ZN => n6115);
   U2303 : OAI22_X1 port map( A1 => n12900, A2 => n13285, B1 => n12893, B2 => 
                           n13565, ZN => n6116);
   U2304 : OAI22_X1 port map( A1 => n12899, A2 => n13288, B1 => n12893, B2 => 
                           n13564, ZN => n6117);
   U2305 : OAI22_X1 port map( A1 => n12899, A2 => n13291, B1 => n12893, B2 => 
                           n13563, ZN => n6118);
   U2306 : OAI22_X1 port map( A1 => n12899, A2 => n13294, B1 => n12893, B2 => 
                           n13562, ZN => n6119);
   U2307 : OAI22_X1 port map( A1 => n12899, A2 => n13297, B1 => n12893, B2 => 
                           n13561, ZN => n6120);
   U2308 : OAI22_X1 port map( A1 => n12899, A2 => n13300, B1 => n12893, B2 => 
                           n13560, ZN => n6121);
   U2309 : OAI22_X1 port map( A1 => n12898, A2 => n13303, B1 => n12893, B2 => 
                           n13559, ZN => n6122);
   U2310 : OAI22_X1 port map( A1 => n12898, A2 => n13306, B1 => n12893, B2 => 
                           n13558, ZN => n6123);
   U2311 : OAI22_X1 port map( A1 => n12898, A2 => n13309, B1 => n12893, B2 => 
                           n13557, ZN => n6124);
   U2312 : OAI22_X1 port map( A1 => n12898, A2 => n13312, B1 => n12893, B2 => 
                           n13556, ZN => n6125);
   U2313 : OAI22_X1 port map( A1 => n12898, A2 => n13315, B1 => n12894, B2 => 
                           n13555, ZN => n6126);
   U2314 : OAI22_X1 port map( A1 => n12897, A2 => n13318, B1 => n12894, B2 => 
                           n13554, ZN => n6127);
   U2315 : OAI22_X1 port map( A1 => n12897, A2 => n13321, B1 => n12894, B2 => 
                           n13553, ZN => n6128);
   U2316 : OAI22_X1 port map( A1 => n12897, A2 => n13324, B1 => n12894, B2 => 
                           n13552, ZN => n6129);
   U2317 : OAI22_X1 port map( A1 => n12897, A2 => n13327, B1 => n12894, B2 => 
                           n13551, ZN => n6130);
   U2318 : OAI22_X1 port map( A1 => n12897, A2 => n13330, B1 => n12894, B2 => 
                           n13550, ZN => n6131);
   U2319 : OAI22_X1 port map( A1 => n12896, A2 => n13333, B1 => n12894, B2 => 
                           n13549, ZN => n6132);
   U2320 : OAI22_X1 port map( A1 => n12896, A2 => n13336, B1 => n12894, B2 => 
                           n13548, ZN => n6133);
   U2321 : OAI22_X1 port map( A1 => n12896, A2 => n13339, B1 => n12894, B2 => 
                           n13547, ZN => n6134);
   U2322 : OAI22_X1 port map( A1 => n12896, A2 => n13342, B1 => n12894, B2 => 
                           n13546, ZN => n6135);
   U2323 : OAI22_X1 port map( A1 => n12896, A2 => n13345, B1 => n12894, B2 => 
                           n13545, ZN => n6136);
   U2324 : OAI22_X1 port map( A1 => n12895, A2 => n13348, B1 => n12894, B2 => 
                           n13544, ZN => n6137);
   U2325 : OAI22_X1 port map( A1 => n12962, A2 => n13242, B1 => n12952, B2 => 
                           n13530, ZN => n6294);
   U2326 : OAI22_X1 port map( A1 => n12962, A2 => n13245, B1 => n12952, B2 => 
                           n13529, ZN => n6295);
   U2327 : OAI22_X1 port map( A1 => n12962, A2 => n13248, B1 => n12952, B2 => 
                           n13528, ZN => n6296);
   U2328 : OAI22_X1 port map( A1 => n12962, A2 => n13251, B1 => n12952, B2 => 
                           n13527, ZN => n6297);
   U2329 : OAI22_X1 port map( A1 => n12962, A2 => n13254, B1 => n12952, B2 => 
                           n13526, ZN => n6298);
   U2330 : OAI22_X1 port map( A1 => n12961, A2 => n13257, B1 => n12952, B2 => 
                           n13525, ZN => n6299);
   U2331 : OAI22_X1 port map( A1 => n12961, A2 => n13260, B1 => n12952, B2 => 
                           n13524, ZN => n6300);
   U2332 : OAI22_X1 port map( A1 => n12961, A2 => n13263, B1 => n12952, B2 => 
                           n13523, ZN => n6301);
   U2333 : OAI22_X1 port map( A1 => n12961, A2 => n13266, B1 => n12952, B2 => 
                           n13522, ZN => n6302);
   U2334 : OAI22_X1 port map( A1 => n12961, A2 => n13269, B1 => n12952, B2 => 
                           n13521, ZN => n6303);
   U2335 : OAI22_X1 port map( A1 => n12960, A2 => n13272, B1 => n12952, B2 => 
                           n13520, ZN => n6304);
   U2336 : OAI22_X1 port map( A1 => n12960, A2 => n13275, B1 => n12952, B2 => 
                           n13519, ZN => n6305);
   U2337 : OAI22_X1 port map( A1 => n12960, A2 => n13278, B1 => n12953, B2 => 
                           n13518, ZN => n6306);
   U2338 : OAI22_X1 port map( A1 => n12960, A2 => n13281, B1 => n12953, B2 => 
                           n13517, ZN => n6307);
   U2339 : OAI22_X1 port map( A1 => n12960, A2 => n13284, B1 => n12953, B2 => 
                           n13516, ZN => n6308);
   U2340 : OAI22_X1 port map( A1 => n12959, A2 => n13299, B1 => n12953, B2 => 
                           n13515, ZN => n6313);
   U2341 : OAI22_X1 port map( A1 => n12958, A2 => n13302, B1 => n12953, B2 => 
                           n13514, ZN => n6314);
   U2342 : OAI22_X1 port map( A1 => n12958, A2 => n13305, B1 => n12953, B2 => 
                           n13513, ZN => n6315);
   U2343 : OAI22_X1 port map( A1 => n12958, A2 => n13308, B1 => n12953, B2 => 
                           n13512, ZN => n6316);
   U2344 : OAI22_X1 port map( A1 => n12958, A2 => n13311, B1 => n12953, B2 => 
                           n13511, ZN => n6317);
   U2345 : OAI22_X1 port map( A1 => n12958, A2 => n13314, B1 => n12954, B2 => 
                           n13510, ZN => n6318);
   U2346 : OAI22_X1 port map( A1 => n12957, A2 => n13317, B1 => n12954, B2 => 
                           n13509, ZN => n6319);
   U2347 : OAI22_X1 port map( A1 => n12957, A2 => n13320, B1 => n12954, B2 => 
                           n13508, ZN => n6320);
   U2348 : OAI22_X1 port map( A1 => n12957, A2 => n13323, B1 => n12954, B2 => 
                           n13507, ZN => n6321);
   U2349 : OAI22_X1 port map( A1 => n12957, A2 => n13326, B1 => n12954, B2 => 
                           n13506, ZN => n6322);
   U2350 : OAI22_X1 port map( A1 => n12957, A2 => n13329, B1 => n12954, B2 => 
                           n13505, ZN => n6323);
   U2351 : OAI22_X1 port map( A1 => n12956, A2 => n13332, B1 => n12954, B2 => 
                           n13504, ZN => n6324);
   U2352 : OAI22_X1 port map( A1 => n12956, A2 => n13335, B1 => n12954, B2 => 
                           n13503, ZN => n6325);
   U2353 : OAI22_X1 port map( A1 => n12956, A2 => n13338, B1 => n12954, B2 => 
                           n13502, ZN => n6326);
   U2354 : OAI22_X1 port map( A1 => n12956, A2 => n13341, B1 => n12954, B2 => 
                           n13501, ZN => n6327);
   U2355 : OAI22_X1 port map( A1 => n12956, A2 => n13344, B1 => n12954, B2 => 
                           n13500, ZN => n6328);
   U2356 : OAI22_X1 port map( A1 => n12955, A2 => n13347, B1 => n12954, B2 => 
                           n13499, ZN => n6329);
   U2357 : OAI22_X1 port map( A1 => n12982, A2 => n13242, B1 => n12972, B2 => 
                           n13470, ZN => n6358);
   U2358 : OAI22_X1 port map( A1 => n12982, A2 => n13245, B1 => n12972, B2 => 
                           n13469, ZN => n6359);
   U2359 : OAI22_X1 port map( A1 => n12982, A2 => n13248, B1 => n12972, B2 => 
                           n13468, ZN => n6360);
   U2360 : OAI22_X1 port map( A1 => n12982, A2 => n13251, B1 => n12972, B2 => 
                           n13467, ZN => n6361);
   U2361 : OAI22_X1 port map( A1 => n12982, A2 => n13254, B1 => n12972, B2 => 
                           n13466, ZN => n6362);
   U2362 : OAI22_X1 port map( A1 => n12981, A2 => n13257, B1 => n12972, B2 => 
                           n13465, ZN => n6363);
   U2363 : OAI22_X1 port map( A1 => n12981, A2 => n13260, B1 => n12972, B2 => 
                           n13464, ZN => n6364);
   U2364 : OAI22_X1 port map( A1 => n12981, A2 => n13263, B1 => n12972, B2 => 
                           n13463, ZN => n6365);
   U2365 : OAI22_X1 port map( A1 => n12981, A2 => n13266, B1 => n12972, B2 => 
                           n13462, ZN => n6366);
   U2366 : OAI22_X1 port map( A1 => n12981, A2 => n13269, B1 => n12972, B2 => 
                           n13461, ZN => n6367);
   U2367 : OAI22_X1 port map( A1 => n12980, A2 => n13272, B1 => n12972, B2 => 
                           n13460, ZN => n6368);
   U2368 : OAI22_X1 port map( A1 => n12980, A2 => n13275, B1 => n12972, B2 => 
                           n13459, ZN => n6369);
   U2369 : OAI22_X1 port map( A1 => n12980, A2 => n13278, B1 => n12973, B2 => 
                           n13458, ZN => n6370);
   U2370 : OAI22_X1 port map( A1 => n12980, A2 => n13281, B1 => n12973, B2 => 
                           n13457, ZN => n6371);
   U2371 : OAI22_X1 port map( A1 => n12980, A2 => n13284, B1 => n12973, B2 => 
                           n13456, ZN => n6372);
   U2372 : OAI22_X1 port map( A1 => n12979, A2 => n13287, B1 => n12973, B2 => 
                           n13455, ZN => n6373);
   U2373 : OAI22_X1 port map( A1 => n12979, A2 => n13290, B1 => n12973, B2 => 
                           n13454, ZN => n6374);
   U2374 : OAI22_X1 port map( A1 => n12979, A2 => n13293, B1 => n12973, B2 => 
                           n13453, ZN => n6375);
   U2375 : OAI22_X1 port map( A1 => n12979, A2 => n13296, B1 => n12973, B2 => 
                           n13452, ZN => n6376);
   U2376 : OAI22_X1 port map( A1 => n12979, A2 => n13299, B1 => n12973, B2 => 
                           n13451, ZN => n6377);
   U2377 : OAI22_X1 port map( A1 => n12978, A2 => n13302, B1 => n12973, B2 => 
                           n13450, ZN => n6378);
   U2378 : OAI22_X1 port map( A1 => n12978, A2 => n13305, B1 => n12973, B2 => 
                           n13449, ZN => n6379);
   U2379 : OAI22_X1 port map( A1 => n12978, A2 => n13308, B1 => n12973, B2 => 
                           n13448, ZN => n6380);
   U2380 : OAI22_X1 port map( A1 => n12978, A2 => n13311, B1 => n12973, B2 => 
                           n13447, ZN => n6381);
   U2381 : OAI22_X1 port map( A1 => n12978, A2 => n13314, B1 => n12974, B2 => 
                           n13446, ZN => n6382);
   U2382 : OAI22_X1 port map( A1 => n12977, A2 => n13317, B1 => n12974, B2 => 
                           n13445, ZN => n6383);
   U2383 : OAI22_X1 port map( A1 => n12977, A2 => n13320, B1 => n12974, B2 => 
                           n13444, ZN => n6384);
   U2384 : OAI22_X1 port map( A1 => n12977, A2 => n13323, B1 => n12974, B2 => 
                           n13443, ZN => n6385);
   U2385 : OAI22_X1 port map( A1 => n12977, A2 => n13326, B1 => n12974, B2 => 
                           n13442, ZN => n6386);
   U2386 : OAI22_X1 port map( A1 => n12977, A2 => n13329, B1 => n12974, B2 => 
                           n13441, ZN => n6387);
   U2387 : OAI22_X1 port map( A1 => n12976, A2 => n13332, B1 => n12974, B2 => 
                           n13440, ZN => n6388);
   U2388 : OAI22_X1 port map( A1 => n12976, A2 => n13335, B1 => n12974, B2 => 
                           n13439, ZN => n6389);
   U2389 : OAI22_X1 port map( A1 => n12976, A2 => n13338, B1 => n12974, B2 => 
                           n13438, ZN => n6390);
   U2390 : OAI22_X1 port map( A1 => n12976, A2 => n13341, B1 => n12974, B2 => 
                           n13437, ZN => n6391);
   U2391 : OAI22_X1 port map( A1 => n12976, A2 => n13344, B1 => n12974, B2 => 
                           n13436, ZN => n6392);
   U2392 : OAI22_X1 port map( A1 => n12975, A2 => n13347, B1 => n12974, B2 => 
                           n13435, ZN => n6393);
   U2393 : OAI22_X1 port map( A1 => n13162, A2 => n13242, B1 => n13152, B2 => 
                           n13406, ZN => n6934);
   U2394 : OAI22_X1 port map( A1 => n13162, A2 => n13245, B1 => n13152, B2 => 
                           n13405, ZN => n6935);
   U2395 : OAI22_X1 port map( A1 => n13162, A2 => n13248, B1 => n13152, B2 => 
                           n13404, ZN => n6936);
   U2396 : OAI22_X1 port map( A1 => n13162, A2 => n13251, B1 => n13152, B2 => 
                           n13403, ZN => n6937);
   U2397 : OAI22_X1 port map( A1 => n13162, A2 => n13254, B1 => n13152, B2 => 
                           n13402, ZN => n6938);
   U2398 : OAI22_X1 port map( A1 => n13367, A2 => n13308, B1 => n13362, B2 => 
                           n13401, ZN => n7020);
   U2399 : OAI22_X1 port map( A1 => n13367, A2 => n13311, B1 => n13362, B2 => 
                           n13400, ZN => n7021);
   U2400 : OAI22_X1 port map( A1 => n13367, A2 => n13314, B1 => n13363, B2 => 
                           n13399, ZN => n7022);
   U2401 : OAI22_X1 port map( A1 => n13366, A2 => n13317, B1 => n13363, B2 => 
                           n13398, ZN => n7023);
   U2402 : OAI22_X1 port map( A1 => n13366, A2 => n13320, B1 => n13363, B2 => 
                           n13397, ZN => n7024);
   U2403 : OAI22_X1 port map( A1 => n13366, A2 => n13323, B1 => n13363, B2 => 
                           n13396, ZN => n7025);
   U2404 : OAI22_X1 port map( A1 => n13366, A2 => n13326, B1 => n13363, B2 => 
                           n13395, ZN => n7026);
   U2405 : OAI22_X1 port map( A1 => n13366, A2 => n13329, B1 => n13363, B2 => 
                           n13394, ZN => n7027);
   U2406 : OAI22_X1 port map( A1 => n13365, A2 => n13332, B1 => n13363, B2 => 
                           n13393, ZN => n7028);
   U2407 : OAI22_X1 port map( A1 => n13364, A2 => n13350, B1 => n13361, B2 => 
                           n14435, ZN => n7034);
   U2408 : OAI22_X1 port map( A1 => n13364, A2 => n13353, B1 => n13362, B2 => 
                           n14434, ZN => n7035);
   U2409 : OAI22_X1 port map( A1 => n13364, A2 => n13356, B1 => n13363, B2 => 
                           n14433, ZN => n7036);
   U2410 : OAI22_X1 port map( A1 => n13155, A2 => n13350, B1 => n13154, B2 => 
                           n14412, ZN => n6970);
   U2411 : OAI22_X1 port map( A1 => n13155, A2 => n13353, B1 => n13153, B2 => 
                           n14411, ZN => n6971);
   U2412 : OAI22_X1 port map( A1 => n13155, A2 => n13356, B1 => n13152, B2 => 
                           n14410, ZN => n6972);
   U2413 : OAI22_X1 port map( A1 => n13155, A2 => n13379, B1 => n13154, B2 => 
                           n14409, ZN => n6973);
   U2414 : OAI22_X1 port map( A1 => n12600, A2 => n13352, B1 => n12599, B2 => 
                           n14086, ZN => n5178);
   U2415 : OAI22_X1 port map( A1 => n12600, A2 => n13355, B1 => n12597, B2 => 
                           n14085, ZN => n5179);
   U2416 : OAI22_X1 port map( A1 => n12600, A2 => n13358, B1 => n12598, B2 => 
                           n14084, ZN => n5180);
   U2417 : OAI22_X1 port map( A1 => n12600, A2 => n13381, B1 => n12599, B2 => 
                           n14083, ZN => n5181);
   U2418 : OAI22_X1 port map( A1 => n13095, A2 => n13350, B1 => n13092, B2 => 
                           n13847, ZN => n6778);
   U2419 : OAI22_X1 port map( A1 => n13095, A2 => n13353, B1 => n13093, B2 => 
                           n13846, ZN => n6779);
   U2420 : OAI22_X1 port map( A1 => n13095, A2 => n13356, B1 => n13094, B2 => 
                           n13845, ZN => n6780);
   U2421 : OAI22_X1 port map( A1 => n13095, A2 => n13379, B1 => n13092, B2 => 
                           n13844, ZN => n6781);
   U2422 : OAI22_X1 port map( A1 => n13075, A2 => n13350, B1 => n13072, B2 => 
                           n13843, ZN => n6714);
   U2423 : OAI22_X1 port map( A1 => n13075, A2 => n13353, B1 => n13073, B2 => 
                           n13842, ZN => n6715);
   U2424 : OAI22_X1 port map( A1 => n13075, A2 => n13356, B1 => n13074, B2 => 
                           n13841, ZN => n6716);
   U2425 : OAI22_X1 port map( A1 => n13075, A2 => n13379, B1 => n13072, B2 => 
                           n13840, ZN => n6717);
   U2426 : OAI22_X1 port map( A1 => n12619, A2 => n13352, B1 => n12616, B2 => 
                           n13750, ZN => n5242);
   U2427 : OAI22_X1 port map( A1 => n12619, A2 => n13355, B1 => n12617, B2 => 
                           n13749, ZN => n5243);
   U2428 : OAI22_X1 port map( A1 => n12619, A2 => n13358, B1 => n12618, B2 => 
                           n13748, ZN => n5244);
   U2429 : OAI22_X1 port map( A1 => n12619, A2 => n13381, B1 => n12616, B2 => 
                           n13747, ZN => n5245);
   U2430 : OAI22_X1 port map( A1 => n12676, A2 => n13352, B1 => n12674, B2 => 
                           n13734, ZN => n5434);
   U2431 : OAI22_X1 port map( A1 => n12676, A2 => n13355, B1 => n12673, B2 => 
                           n13733, ZN => n5435);
   U2432 : OAI22_X1 port map( A1 => n12676, A2 => n13358, B1 => n12675, B2 => 
                           n13732, ZN => n5436);
   U2433 : OAI22_X1 port map( A1 => n12676, A2 => n13381, B1 => n12674, B2 => 
                           n13731, ZN => n5437);
   U2434 : OAI22_X1 port map( A1 => n12695, A2 => n13352, B1 => n12692, B2 => 
                           n13670, ZN => n5498);
   U2435 : OAI22_X1 port map( A1 => n12695, A2 => n13355, B1 => n12693, B2 => 
                           n13669, ZN => n5499);
   U2436 : OAI22_X1 port map( A1 => n12695, A2 => n13358, B1 => n12694, B2 => 
                           n13668, ZN => n5500);
   U2437 : OAI22_X1 port map( A1 => n12695, A2 => n13381, B1 => n12692, B2 => 
                           n13667, ZN => n5501);
   U2438 : OAI22_X1 port map( A1 => n12875, A2 => n13351, B1 => n12872, B2 => 
                           n13607, ZN => n6074);
   U2439 : OAI22_X1 port map( A1 => n12875, A2 => n13354, B1 => n12873, B2 => 
                           n13606, ZN => n6075);
   U2440 : OAI22_X1 port map( A1 => n12875, A2 => n13357, B1 => n12874, B2 => 
                           n13605, ZN => n6076);
   U2441 : OAI22_X1 port map( A1 => n12875, A2 => n13380, B1 => n12872, B2 => 
                           n13604, ZN => n6077);
   U2442 : OAI22_X1 port map( A1 => n12895, A2 => n13351, B1 => n12892, B2 => 
                           n13543, ZN => n6138);
   U2443 : OAI22_X1 port map( A1 => n12895, A2 => n13354, B1 => n12893, B2 => 
                           n13542, ZN => n6139);
   U2444 : OAI22_X1 port map( A1 => n12895, A2 => n13357, B1 => n12894, B2 => 
                           n13541, ZN => n6140);
   U2445 : OAI22_X1 port map( A1 => n12895, A2 => n13380, B1 => n12892, B2 => 
                           n13540, ZN => n6141);
   U2446 : OAI22_X1 port map( A1 => n12955, A2 => n13350, B1 => n12952, B2 => 
                           n13498, ZN => n6330);
   U2447 : OAI22_X1 port map( A1 => n12955, A2 => n13353, B1 => n12953, B2 => 
                           n13497, ZN => n6331);
   U2448 : OAI22_X1 port map( A1 => n12955, A2 => n13356, B1 => n12954, B2 => 
                           n13496, ZN => n6332);
   U2449 : OAI22_X1 port map( A1 => n12955, A2 => n13379, B1 => n12952, B2 => 
                           n13495, ZN => n6333);
   U2450 : OAI22_X1 port map( A1 => n12975, A2 => n13350, B1 => n12972, B2 => 
                           n13434, ZN => n6394);
   U2451 : OAI22_X1 port map( A1 => n12975, A2 => n13353, B1 => n12973, B2 => 
                           n13433, ZN => n6395);
   U2452 : OAI22_X1 port map( A1 => n12975, A2 => n13356, B1 => n12974, B2 => 
                           n13432, ZN => n6396);
   U2453 : OAI22_X1 port map( A1 => n12975, A2 => n13379, B1 => n12972, B2 => 
                           n13431, ZN => n6397);
   U2454 : OAI22_X1 port map( A1 => n13364, A2 => n13379, B1 => n13361, B2 => 
                           n13392, ZN => n7037);
   U2455 : INV_X1 port map( A => ADD_RD1(3), ZN => n14462);
   U2456 : INV_X1 port map( A => ADD_RD1(4), ZN => n14461);
   U2457 : INV_X1 port map( A => ADD_RD1(0), ZN => n14465);
   U2458 : INV_X1 port map( A => ADD_RD1(1), ZN => n14464);
   U2459 : INV_X1 port map( A => ADD_RD1(2), ZN => n14463);
   U2460 : INV_X1 port map( A => ADD_WR(2), ZN => n13384);
   U2461 : INV_X1 port map( A => ADD_WR(0), ZN => n13386);
   U2462 : INV_X1 port map( A => ADD_WR(1), ZN => n13385);
   U2463 : INV_X1 port map( A => ADD_WR(3), ZN => n13383);
   U2464 : NOR2_X1 port map( A1 => n13389, A2 => n13390, ZN => n4455);
   U2465 : NOR3_X1 port map( A1 => n13391, A2 => n13387, A3 => n13388, ZN => 
                           n4470);
   U2466 : AOI221_X1 port map( B1 => n12302, B2 => n11586, C1 => n12296, C2 => 
                           n11406, A => n4453, ZN => n4446);
   U2467 : OAI22_X1 port map( A1 => n14362, A2 => n12290, B1 => n14361, B2 => 
                           n12284, ZN => n4453);
   U2468 : AOI221_X1 port map( B1 => n12302, B2 => n11587, C1 => n12296, C2 => 
                           n11407, A => n4411, ZN => n4408);
   U2469 : OAI22_X1 port map( A1 => n14407, A2 => n12290, B1 => n14384, B2 => 
                           n12284, ZN => n4411);
   U2470 : AOI221_X1 port map( B1 => n12302, B2 => n11588, C1 => n12296, C2 => 
                           n11408, A => n4392, ZN => n4389);
   U2471 : OAI22_X1 port map( A1 => n14406, A2 => n12290, B1 => n14383, B2 => 
                           n12284, ZN => n4392);
   U2472 : AOI221_X1 port map( B1 => n12302, B2 => n11589, C1 => n12296, C2 => 
                           n11409, A => n4373, ZN => n4370);
   U2473 : OAI22_X1 port map( A1 => n14405, A2 => n12290, B1 => n14382, B2 => 
                           n12284, ZN => n4373);
   U2474 : AOI221_X1 port map( B1 => n12302, B2 => n11590, C1 => n12296, C2 => 
                           n11410, A => n4316, ZN => n4313);
   U2475 : OAI22_X1 port map( A1 => n14402, A2 => n12290, B1 => n14379, B2 => 
                           n12284, ZN => n4316);
   U2476 : AOI221_X1 port map( B1 => n12302, B2 => n11591, C1 => n12296, C2 => 
                           n11411, A => n4297, ZN => n4294);
   U2477 : OAI22_X1 port map( A1 => n14401, A2 => n12290, B1 => n14378, B2 => 
                           n12284, ZN => n4297);
   U2478 : AOI221_X1 port map( B1 => n12302, B2 => n11592, C1 => n12296, C2 => 
                           n11412, A => n4278, ZN => n4275);
   U2479 : OAI22_X1 port map( A1 => n14400, A2 => n12290, B1 => n14377, B2 => 
                           n12284, ZN => n4278);
   U2480 : AOI221_X1 port map( B1 => n12302, B2 => n11593, C1 => n12296, C2 => 
                           n11413, A => n4259, ZN => n4256);
   U2481 : OAI22_X1 port map( A1 => n14399, A2 => n12290, B1 => n14376, B2 => 
                           n12284, ZN => n4259);
   U2482 : AOI221_X1 port map( B1 => n12302, B2 => n11594, C1 => n12296, C2 => 
                           n11414, A => n4240, ZN => n4237);
   U2483 : OAI22_X1 port map( A1 => n14398, A2 => n12290, B1 => n14375, B2 => 
                           n12284, ZN => n4240);
   U2484 : AOI221_X1 port map( B1 => n12303, B2 => n11595, C1 => n12297, C2 => 
                           n11415, A => n4221, ZN => n4218);
   U2485 : OAI22_X1 port map( A1 => n14397, A2 => n12291, B1 => n14374, B2 => 
                           n12285, ZN => n4221);
   U2486 : AOI221_X1 port map( B1 => n12303, B2 => n11596, C1 => n12297, C2 => 
                           n11416, A => n4202, ZN => n4199);
   U2487 : OAI22_X1 port map( A1 => n14396, A2 => n12291, B1 => n14373, B2 => 
                           n12285, ZN => n4202);
   U2488 : AOI221_X1 port map( B1 => n12303, B2 => n11597, C1 => n12297, C2 => 
                           n11417, A => n4183, ZN => n4180);
   U2489 : OAI22_X1 port map( A1 => n14395, A2 => n12291, B1 => n14372, B2 => 
                           n12285, ZN => n4183);
   U2490 : AOI221_X1 port map( B1 => n12303, B2 => n11598, C1 => n12297, C2 => 
                           n11418, A => n4164, ZN => n4161);
   U2491 : OAI22_X1 port map( A1 => n14394, A2 => n12291, B1 => n14371, B2 => 
                           n12285, ZN => n4164);
   U2492 : AOI221_X1 port map( B1 => n12303, B2 => n11599, C1 => n12297, C2 => 
                           n11419, A => n4145, ZN => n4142);
   U2493 : OAI22_X1 port map( A1 => n14393, A2 => n12291, B1 => n14370, B2 => 
                           n12285, ZN => n4145);
   U2494 : AOI221_X1 port map( B1 => n12303, B2 => n11600, C1 => n12297, C2 => 
                           n11420, A => n4126, ZN => n4123);
   U2495 : OAI22_X1 port map( A1 => n14392, A2 => n12291, B1 => n14369, B2 => 
                           n12285, ZN => n4126);
   U2496 : AOI221_X1 port map( B1 => n12303, B2 => n11601, C1 => n12297, C2 => 
                           n11421, A => n4107, ZN => n4104);
   U2497 : OAI22_X1 port map( A1 => n14391, A2 => n12291, B1 => n14368, B2 => 
                           n12285, ZN => n4107);
   U2498 : AOI221_X1 port map( B1 => n12303, B2 => n11602, C1 => n12297, C2 => 
                           n11422, A => n4088, ZN => n4085);
   U2499 : OAI22_X1 port map( A1 => n14390, A2 => n12291, B1 => n14367, B2 => 
                           n12285, ZN => n4088);
   U2500 : AOI221_X1 port map( B1 => n12303, B2 => n11603, C1 => n12297, C2 => 
                           n11423, A => n4069, ZN => n4066);
   U2501 : OAI22_X1 port map( A1 => n14389, A2 => n12291, B1 => n14366, B2 => 
                           n12285, ZN => n4069);
   U2502 : AOI221_X1 port map( B1 => n12303, B2 => n11604, C1 => n12297, C2 => 
                           n11424, A => n4050, ZN => n4047);
   U2503 : OAI22_X1 port map( A1 => n14388, A2 => n12291, B1 => n14365, B2 => 
                           n12285, ZN => n4050);
   U2504 : AOI221_X1 port map( B1 => n12303, B2 => n11605, C1 => n12297, C2 => 
                           n11425, A => n4031, ZN => n4028);
   U2505 : OAI22_X1 port map( A1 => n14387, A2 => n12291, B1 => n14364, B2 => 
                           n12285, ZN => n4031);
   U2506 : AOI221_X1 port map( B1 => n12303, B2 => n11606, C1 => n12297, C2 => 
                           n11426, A => n4012, ZN => n4009);
   U2507 : OAI22_X1 port map( A1 => n14386, A2 => n12291, B1 => n14363, B2 => 
                           n12285, ZN => n4012);
   U2508 : AOI221_X1 port map( B1 => n12304, B2 => n11607, C1 => n12298, C2 => 
                           n11427, A => n3993, ZN => n3990);
   U2509 : OAI22_X1 port map( A1 => n14288, A2 => n12292, B1 => n14252, B2 => 
                           n12286, ZN => n3993);
   U2510 : AOI221_X1 port map( B1 => n12304, B2 => n11608, C1 => n12298, C2 => 
                           n11428, A => n3974, ZN => n3971);
   U2511 : OAI22_X1 port map( A1 => n14287, A2 => n12292, B1 => n14251, B2 => 
                           n12286, ZN => n3974);
   U2512 : AOI221_X1 port map( B1 => n12304, B2 => n11609, C1 => n12298, C2 => 
                           n11429, A => n3955, ZN => n3952);
   U2513 : OAI22_X1 port map( A1 => n14286, A2 => n12292, B1 => n14250, B2 => 
                           n12286, ZN => n3955);
   U2514 : AOI221_X1 port map( B1 => n12304, B2 => n11610, C1 => n12298, C2 => 
                           n11430, A => n3936, ZN => n3933);
   U2515 : OAI22_X1 port map( A1 => n14285, A2 => n12292, B1 => n14249, B2 => 
                           n12286, ZN => n3936);
   U2516 : AOI221_X1 port map( B1 => n12304, B2 => n11611, C1 => n12298, C2 => 
                           n11431, A => n3917, ZN => n3914);
   U2517 : OAI22_X1 port map( A1 => n14284, A2 => n12292, B1 => n14248, B2 => 
                           n12286, ZN => n3917);
   U2518 : AOI221_X1 port map( B1 => n12304, B2 => n11612, C1 => n12298, C2 => 
                           n11432, A => n3898, ZN => n3895);
   U2519 : OAI22_X1 port map( A1 => n14283, A2 => n12292, B1 => n14247, B2 => 
                           n12286, ZN => n3898);
   U2520 : AOI221_X1 port map( B1 => n12304, B2 => n11613, C1 => n12298, C2 => 
                           n11433, A => n3879, ZN => n3876);
   U2521 : OAI22_X1 port map( A1 => n14282, A2 => n12292, B1 => n14246, B2 => 
                           n12286, ZN => n3879);
   U2522 : AOI221_X1 port map( B1 => n12304, B2 => n11614, C1 => n12298, C2 => 
                           n11434, A => n3860, ZN => n3857);
   U2523 : OAI22_X1 port map( A1 => n14281, A2 => n12292, B1 => n14245, B2 => 
                           n12286, ZN => n3860);
   U2524 : AOI221_X1 port map( B1 => n12304, B2 => n11615, C1 => n12298, C2 => 
                           n11435, A => n3841, ZN => n3838);
   U2525 : OAI22_X1 port map( A1 => n14280, A2 => n12292, B1 => n14244, B2 => 
                           n12286, ZN => n3841);
   U2526 : AOI221_X1 port map( B1 => n12304, B2 => n11616, C1 => n12298, C2 => 
                           n11436, A => n3822, ZN => n3819);
   U2527 : OAI22_X1 port map( A1 => n14279, A2 => n12292, B1 => n14243, B2 => 
                           n12286, ZN => n3822);
   U2528 : AOI221_X1 port map( B1 => n12304, B2 => n11617, C1 => n12298, C2 => 
                           n11437, A => n3803, ZN => n3800);
   U2529 : OAI22_X1 port map( A1 => n14278, A2 => n12292, B1 => n14242, B2 => 
                           n12286, ZN => n3803);
   U2530 : AOI221_X1 port map( B1 => n12304, B2 => n11618, C1 => n12298, C2 => 
                           n11438, A => n3784, ZN => n3781);
   U2531 : OAI22_X1 port map( A1 => n14277, A2 => n12292, B1 => n14241, B2 => 
                           n12286, ZN => n3784);
   U2532 : AOI221_X1 port map( B1 => n12305, B2 => n11619, C1 => n12299, C2 => 
                           n11439, A => n3765, ZN => n3762);
   U2533 : OAI22_X1 port map( A1 => n14276, A2 => n12293, B1 => n14240, B2 => 
                           n12287, ZN => n3765);
   U2534 : AOI221_X1 port map( B1 => n12305, B2 => n11620, C1 => n12299, C2 => 
                           n11440, A => n3746, ZN => n3743);
   U2535 : OAI22_X1 port map( A1 => n14275, A2 => n12293, B1 => n14239, B2 => 
                           n12287, ZN => n3746);
   U2536 : AOI221_X1 port map( B1 => n12305, B2 => n11621, C1 => n12299, C2 => 
                           n11441, A => n3727, ZN => n3724);
   U2537 : OAI22_X1 port map( A1 => n14274, A2 => n12293, B1 => n14238, B2 => 
                           n12287, ZN => n3727);
   U2538 : AOI221_X1 port map( B1 => n12305, B2 => n11622, C1 => n12299, C2 => 
                           n11442, A => n3708, ZN => n3705);
   U2539 : OAI22_X1 port map( A1 => n14273, A2 => n12293, B1 => n14237, B2 => 
                           n12287, ZN => n3708);
   U2540 : AOI221_X1 port map( B1 => n12305, B2 => n11623, C1 => n12299, C2 => 
                           n11443, A => n3689, ZN => n3686);
   U2541 : OAI22_X1 port map( A1 => n14272, A2 => n12293, B1 => n14236, B2 => 
                           n12287, ZN => n3689);
   U2542 : AOI221_X1 port map( B1 => n12305, B2 => n11624, C1 => n12299, C2 => 
                           n11444, A => n3670, ZN => n3667);
   U2543 : OAI22_X1 port map( A1 => n14271, A2 => n12293, B1 => n14235, B2 => 
                           n12287, ZN => n3670);
   U2544 : AOI221_X1 port map( B1 => n12305, B2 => n11625, C1 => n12299, C2 => 
                           n11445, A => n3651, ZN => n3648);
   U2545 : OAI22_X1 port map( A1 => n14270, A2 => n12293, B1 => n14234, B2 => 
                           n12287, ZN => n3651);
   U2546 : AOI221_X1 port map( B1 => n12305, B2 => n11626, C1 => n12299, C2 => 
                           n11446, A => n3632, ZN => n3629);
   U2547 : OAI22_X1 port map( A1 => n14269, A2 => n12293, B1 => n14233, B2 => 
                           n12287, ZN => n3632);
   U2548 : AOI221_X1 port map( B1 => n12305, B2 => n11627, C1 => n12299, C2 => 
                           n11447, A => n3613, ZN => n3610);
   U2549 : OAI22_X1 port map( A1 => n14268, A2 => n12293, B1 => n14232, B2 => 
                           n12287, ZN => n3613);
   U2550 : AOI221_X1 port map( B1 => n12305, B2 => n11628, C1 => n12299, C2 => 
                           n11448, A => n3594, ZN => n3591);
   U2551 : OAI22_X1 port map( A1 => n14267, A2 => n12293, B1 => n14231, B2 => 
                           n12287, ZN => n3594);
   U2552 : AOI221_X1 port map( B1 => n12305, B2 => n11629, C1 => n12299, C2 => 
                           n11449, A => n3575, ZN => n3572);
   U2553 : OAI22_X1 port map( A1 => n14266, A2 => n12293, B1 => n14230, B2 => 
                           n12287, ZN => n3575);
   U2554 : AOI221_X1 port map( B1 => n12305, B2 => n11630, C1 => n12299, C2 => 
                           n11450, A => n3556, ZN => n3553);
   U2555 : OAI22_X1 port map( A1 => n14265, A2 => n12293, B1 => n14229, B2 => 
                           n12287, ZN => n3556);
   U2556 : AOI221_X1 port map( B1 => n12306, B2 => n11631, C1 => n12300, C2 => 
                           n11451, A => n3537, ZN => n3534);
   U2557 : OAI22_X1 port map( A1 => n14264, A2 => n12294, B1 => n14228, B2 => 
                           n12288, ZN => n3537);
   U2558 : AOI221_X1 port map( B1 => n12306, B2 => n11632, C1 => n12300, C2 => 
                           n11452, A => n3518, ZN => n3515);
   U2559 : OAI22_X1 port map( A1 => n14263, A2 => n12294, B1 => n14227, B2 => 
                           n12288, ZN => n3518);
   U2560 : AOI221_X1 port map( B1 => n12306, B2 => n11633, C1 => n12300, C2 => 
                           n11453, A => n3499, ZN => n3496);
   U2561 : OAI22_X1 port map( A1 => n14262, A2 => n12294, B1 => n14226, B2 => 
                           n12288, ZN => n3499);
   U2562 : AOI221_X1 port map( B1 => n12306, B2 => n11634, C1 => n12300, C2 => 
                           n11454, A => n3480, ZN => n3477);
   U2563 : OAI22_X1 port map( A1 => n14261, A2 => n12294, B1 => n14225, B2 => 
                           n12288, ZN => n3480);
   U2564 : AOI221_X1 port map( B1 => n12306, B2 => n11635, C1 => n12300, C2 => 
                           n11455, A => n3461, ZN => n3458);
   U2565 : OAI22_X1 port map( A1 => n14260, A2 => n12294, B1 => n14224, B2 => 
                           n12288, ZN => n3461);
   U2566 : AOI221_X1 port map( B1 => n12306, B2 => n11636, C1 => n12300, C2 => 
                           n11456, A => n3442, ZN => n3439);
   U2567 : OAI22_X1 port map( A1 => n14259, A2 => n12294, B1 => n14223, B2 => 
                           n12288, ZN => n3442);
   U2568 : AOI221_X1 port map( B1 => n12306, B2 => n11637, C1 => n12300, C2 => 
                           n11457, A => n3423, ZN => n3420);
   U2569 : OAI22_X1 port map( A1 => n14258, A2 => n12294, B1 => n14222, B2 => 
                           n12288, ZN => n3423);
   U2570 : AOI221_X1 port map( B1 => n12306, B2 => n11638, C1 => n12300, C2 => 
                           n11458, A => n3404, ZN => n3401);
   U2571 : OAI22_X1 port map( A1 => n14257, A2 => n12294, B1 => n14221, B2 => 
                           n12288, ZN => n3404);
   U2572 : AOI221_X1 port map( B1 => n12306, B2 => n11639, C1 => n12300, C2 => 
                           n11459, A => n3385, ZN => n3382);
   U2573 : OAI22_X1 port map( A1 => n14256, A2 => n12294, B1 => n14220, B2 => 
                           n12288, ZN => n3385);
   U2574 : AOI221_X1 port map( B1 => n12306, B2 => n11640, C1 => n12300, C2 => 
                           n11460, A => n3366, ZN => n3363);
   U2575 : OAI22_X1 port map( A1 => n14255, A2 => n12294, B1 => n14219, B2 => 
                           n12288, ZN => n3366);
   U2576 : AOI221_X1 port map( B1 => n12306, B2 => n11641, C1 => n12300, C2 => 
                           n11461, A => n3347, ZN => n3344);
   U2577 : OAI22_X1 port map( A1 => n14254, A2 => n12294, B1 => n14218, B2 => 
                           n12288, ZN => n3347);
   U2578 : AOI221_X1 port map( B1 => n12307, B2 => n13835, C1 => n12301, C2 => 
                           n13839, A => n3309, ZN => n3306);
   U2579 : OAI22_X1 port map( A1 => n13847, A2 => n12295, B1 => n13843, B2 => 
                           n12289, ZN => n3309);
   U2580 : AOI221_X1 port map( B1 => n12307, B2 => n13834, C1 => n12301, C2 => 
                           n13838, A => n3290, ZN => n3287);
   U2581 : OAI22_X1 port map( A1 => n13846, A2 => n12295, B1 => n13842, B2 => 
                           n12289, ZN => n3290);
   U2582 : AOI221_X1 port map( B1 => n12307, B2 => n13833, C1 => n12301, C2 => 
                           n13837, A => n3271, ZN => n3268);
   U2583 : OAI22_X1 port map( A1 => n13845, A2 => n12295, B1 => n13841, B2 => 
                           n12289, ZN => n3271);
   U2584 : AOI221_X1 port map( B1 => n12307, B2 => n13832, C1 => n12301, C2 => 
                           n13836, A => n3226, ZN => n3217);
   U2585 : OAI22_X1 port map( A1 => n13844, A2 => n12295, B1 => n13840, B2 => 
                           n12289, ZN => n3226);
   U2586 : AOI221_X1 port map( B1 => n12278, B2 => n11642, C1 => n12272, C2 => 
                           n11462, A => n4456, ZN => n4445);
   U2587 : OAI22_X1 port map( A1 => n13539, A2 => n12266, B1 => n13494, B2 => 
                           n12260, ZN => n4456);
   U2588 : AOI221_X1 port map( B1 => n12182, B2 => n14153, C1 => n12176, C2 => 
                           n14154, A => n4468, ZN => n4461);
   U2589 : OAI22_X1 port map( A1 => n13746, A2 => n12170, B1 => n13730, B2 => 
                           n12164, ZN => n4468);
   U2590 : AOI221_X1 port map( B1 => n12278, B2 => n11643, C1 => n12272, C2 => 
                           n11463, A => n4431, ZN => n4426);
   U2591 : OAI22_X1 port map( A1 => n13538, A2 => n12266, B1 => n13493, B2 => 
                           n12260, ZN => n4431);
   U2592 : AOI221_X1 port map( B1 => n12182, B2 => n14082, C1 => n12176, C2 => 
                           n14129, A => n4439, ZN => n4434);
   U2593 : OAI22_X1 port map( A1 => n13745, A2 => n12170, B1 => n13729, B2 => 
                           n12164, ZN => n4439);
   U2594 : AOI221_X1 port map( B1 => n12278, B2 => n11644, C1 => n12272, C2 => 
                           n11464, A => n4412, ZN => n4407);
   U2595 : OAI22_X1 port map( A1 => n13537, A2 => n12266, B1 => n13492, B2 => 
                           n12260, ZN => n4412);
   U2596 : AOI221_X1 port map( B1 => n12182, B2 => n14081, C1 => n12176, C2 => 
                           n14128, A => n4420, ZN => n4415);
   U2597 : OAI22_X1 port map( A1 => n13744, A2 => n12170, B1 => n13728, B2 => 
                           n12164, ZN => n4420);
   U2598 : AOI221_X1 port map( B1 => n12278, B2 => n11645, C1 => n12272, C2 => 
                           n11465, A => n4393, ZN => n4388);
   U2599 : OAI22_X1 port map( A1 => n13536, A2 => n12266, B1 => n13491, B2 => 
                           n12260, ZN => n4393);
   U2600 : AOI221_X1 port map( B1 => n12182, B2 => n14079, C1 => n12176, C2 => 
                           n14126, A => n4401, ZN => n4396);
   U2601 : OAI22_X1 port map( A1 => n13743, A2 => n12170, B1 => n13727, B2 => 
                           n12164, ZN => n4401);
   U2602 : AOI221_X1 port map( B1 => n12278, B2 => n11646, C1 => n12272, C2 => 
                           n11466, A => n4374, ZN => n4369);
   U2603 : OAI22_X1 port map( A1 => n14360, A2 => n12266, B1 => n13490, B2 => 
                           n12260, ZN => n4374);
   U2604 : AOI221_X1 port map( B1 => n12182, B2 => n14080, C1 => n12176, C2 => 
                           n14127, A => n4382, ZN => n4377);
   U2605 : OAI22_X1 port map( A1 => n13892, A2 => n12170, B1 => n13726, B2 => 
                           n12164, ZN => n4382);
   U2606 : AOI221_X1 port map( B1 => n12278, B2 => n11647, C1 => n12272, C2 => 
                           n11467, A => n4355, ZN => n4350);
   U2607 : OAI22_X1 port map( A1 => n14359, A2 => n12266, B1 => n13489, B2 => 
                           n12260, ZN => n4355);
   U2608 : AOI221_X1 port map( B1 => n12182, B2 => n14078, C1 => n12176, C2 => 
                           n14125, A => n4363, ZN => n4358);
   U2609 : OAI22_X1 port map( A1 => n13891, A2 => n12170, B1 => n13725, B2 => 
                           n12164, ZN => n4363);
   U2610 : AOI221_X1 port map( B1 => n12278, B2 => n11648, C1 => n12272, C2 => 
                           n11468, A => n4336, ZN => n4331);
   U2611 : OAI22_X1 port map( A1 => n14358, A2 => n12266, B1 => n13488, B2 => 
                           n12260, ZN => n4336);
   U2612 : AOI221_X1 port map( B1 => n12182, B2 => n14077, C1 => n12176, C2 => 
                           n14124, A => n4344, ZN => n4339);
   U2613 : OAI22_X1 port map( A1 => n13890, A2 => n12170, B1 => n13724, B2 => 
                           n12164, ZN => n4344);
   U2614 : AOI221_X1 port map( B1 => n12278, B2 => n11649, C1 => n12272, C2 => 
                           n11469, A => n4317, ZN => n4312);
   U2615 : OAI22_X1 port map( A1 => n14340, A2 => n12266, B1 => n13487, B2 => 
                           n12260, ZN => n4317);
   U2616 : AOI221_X1 port map( B1 => n12182, B2 => n14076, C1 => n12176, C2 => 
                           n14123, A => n4325, ZN => n4320);
   U2617 : OAI22_X1 port map( A1 => n13889, A2 => n12170, B1 => n13723, B2 => 
                           n12164, ZN => n4325);
   U2618 : AOI221_X1 port map( B1 => n12278, B2 => n11650, C1 => n12272, C2 => 
                           n11470, A => n4298, ZN => n4293);
   U2619 : OAI22_X1 port map( A1 => n14339, A2 => n12266, B1 => n13486, B2 => 
                           n12260, ZN => n4298);
   U2620 : AOI221_X1 port map( B1 => n12182, B2 => n14075, C1 => n12176, C2 => 
                           n14122, A => n4306, ZN => n4301);
   U2621 : OAI22_X1 port map( A1 => n13888, A2 => n12170, B1 => n13722, B2 => 
                           n12164, ZN => n4306);
   U2622 : AOI221_X1 port map( B1 => n12278, B2 => n11651, C1 => n12272, C2 => 
                           n11471, A => n4279, ZN => n4274);
   U2623 : OAI22_X1 port map( A1 => n14338, A2 => n12266, B1 => n13485, B2 => 
                           n12260, ZN => n4279);
   U2624 : AOI221_X1 port map( B1 => n12182, B2 => n14074, C1 => n12176, C2 => 
                           n14121, A => n4287, ZN => n4282);
   U2625 : OAI22_X1 port map( A1 => n13887, A2 => n12170, B1 => n13721, B2 => 
                           n12164, ZN => n4287);
   U2626 : AOI221_X1 port map( B1 => n12278, B2 => n11652, C1 => n12272, C2 => 
                           n11472, A => n4260, ZN => n4255);
   U2627 : OAI22_X1 port map( A1 => n14337, A2 => n12266, B1 => n13484, B2 => 
                           n12260, ZN => n4260);
   U2628 : AOI221_X1 port map( B1 => n12182, B2 => n14073, C1 => n12176, C2 => 
                           n14120, A => n4268, ZN => n4263);
   U2629 : OAI22_X1 port map( A1 => n13886, A2 => n12170, B1 => n13720, B2 => 
                           n12164, ZN => n4268);
   U2630 : AOI221_X1 port map( B1 => n12278, B2 => n11653, C1 => n12272, C2 => 
                           n11473, A => n4241, ZN => n4236);
   U2631 : OAI22_X1 port map( A1 => n14336, A2 => n12266, B1 => n13483, B2 => 
                           n12260, ZN => n4241);
   U2632 : AOI221_X1 port map( B1 => n12182, B2 => n14072, C1 => n12176, C2 => 
                           n14119, A => n4249, ZN => n4244);
   U2633 : OAI22_X1 port map( A1 => n13885, A2 => n12170, B1 => n13719, B2 => 
                           n12164, ZN => n4249);
   U2634 : AOI221_X1 port map( B1 => n12279, B2 => n11654, C1 => n12273, C2 => 
                           n11474, A => n4222, ZN => n4217);
   U2635 : OAI22_X1 port map( A1 => n14335, A2 => n12267, B1 => n13482, B2 => 
                           n12261, ZN => n4222);
   U2636 : AOI221_X1 port map( B1 => n12183, B2 => n14071, C1 => n12177, C2 => 
                           n14118, A => n4230, ZN => n4225);
   U2637 : OAI22_X1 port map( A1 => n13884, A2 => n12171, B1 => n13718, B2 => 
                           n12165, ZN => n4230);
   U2638 : AOI221_X1 port map( B1 => n12279, B2 => n11655, C1 => n12273, C2 => 
                           n11475, A => n4203, ZN => n4198);
   U2639 : OAI22_X1 port map( A1 => n14334, A2 => n12267, B1 => n13481, B2 => 
                           n12261, ZN => n4203);
   U2640 : AOI221_X1 port map( B1 => n12183, B2 => n14070, C1 => n12177, C2 => 
                           n14117, A => n4211, ZN => n4206);
   U2641 : OAI22_X1 port map( A1 => n13883, A2 => n12171, B1 => n13717, B2 => 
                           n12165, ZN => n4211);
   U2642 : AOI221_X1 port map( B1 => n12279, B2 => n11656, C1 => n12273, C2 => 
                           n11476, A => n4184, ZN => n4179);
   U2643 : OAI22_X1 port map( A1 => n14333, A2 => n12267, B1 => n13480, B2 => 
                           n12261, ZN => n4184);
   U2644 : AOI221_X1 port map( B1 => n12183, B2 => n14069, C1 => n12177, C2 => 
                           n14116, A => n4192, ZN => n4187);
   U2645 : OAI22_X1 port map( A1 => n13882, A2 => n12171, B1 => n13716, B2 => 
                           n12165, ZN => n4192);
   U2646 : AOI221_X1 port map( B1 => n12279, B2 => n11657, C1 => n12273, C2 => 
                           n11477, A => n4165, ZN => n4160);
   U2647 : OAI22_X1 port map( A1 => n14332, A2 => n12267, B1 => n13479, B2 => 
                           n12261, ZN => n4165);
   U2648 : AOI221_X1 port map( B1 => n12183, B2 => n14068, C1 => n12177, C2 => 
                           n14115, A => n4173, ZN => n4168);
   U2649 : OAI22_X1 port map( A1 => n13881, A2 => n12171, B1 => n13715, B2 => 
                           n12165, ZN => n4173);
   U2650 : AOI221_X1 port map( B1 => n12279, B2 => n11658, C1 => n12273, C2 => 
                           n11478, A => n4146, ZN => n4141);
   U2651 : OAI22_X1 port map( A1 => n13535, A2 => n12267, B1 => n13478, B2 => 
                           n12261, ZN => n4146);
   U2652 : AOI221_X1 port map( B1 => n12183, B2 => n14067, C1 => n12177, C2 => 
                           n14114, A => n4154, ZN => n4149);
   U2653 : OAI22_X1 port map( A1 => n13880, A2 => n12171, B1 => n13714, B2 => 
                           n12165, ZN => n4154);
   U2654 : AOI221_X1 port map( B1 => n12279, B2 => n11659, C1 => n12273, C2 => 
                           n11479, A => n4127, ZN => n4122);
   U2655 : OAI22_X1 port map( A1 => n14331, A2 => n12267, B1 => n13477, B2 => 
                           n12261, ZN => n4127);
   U2656 : AOI221_X1 port map( B1 => n12183, B2 => n14066, C1 => n12177, C2 => 
                           n14113, A => n4135, ZN => n4130);
   U2657 : OAI22_X1 port map( A1 => n13879, A2 => n12171, B1 => n13713, B2 => 
                           n12165, ZN => n4135);
   U2658 : AOI221_X1 port map( B1 => n12279, B2 => n11660, C1 => n12273, C2 => 
                           n11480, A => n4108, ZN => n4103);
   U2659 : OAI22_X1 port map( A1 => n14330, A2 => n12267, B1 => n13476, B2 => 
                           n12261, ZN => n4108);
   U2660 : AOI221_X1 port map( B1 => n12183, B2 => n14065, C1 => n12177, C2 => 
                           n14112, A => n4116, ZN => n4111);
   U2661 : OAI22_X1 port map( A1 => n13878, A2 => n12171, B1 => n13712, B2 => 
                           n12165, ZN => n4116);
   U2662 : AOI221_X1 port map( B1 => n12279, B2 => n11661, C1 => n12273, C2 => 
                           n11481, A => n4089, ZN => n4084);
   U2663 : OAI22_X1 port map( A1 => n14329, A2 => n12267, B1 => n13475, B2 => 
                           n12261, ZN => n4089);
   U2664 : AOI221_X1 port map( B1 => n12183, B2 => n14064, C1 => n12177, C2 => 
                           n14111, A => n4097, ZN => n4092);
   U2665 : OAI22_X1 port map( A1 => n13877, A2 => n12171, B1 => n13711, B2 => 
                           n12165, ZN => n4097);
   U2666 : AOI221_X1 port map( B1 => n12279, B2 => n11662, C1 => n12273, C2 => 
                           n11482, A => n4070, ZN => n4065);
   U2667 : OAI22_X1 port map( A1 => n13534, A2 => n12267, B1 => n13474, B2 => 
                           n12261, ZN => n4070);
   U2668 : AOI221_X1 port map( B1 => n12183, B2 => n14063, C1 => n12177, C2 => 
                           n14110, A => n4078, ZN => n4073);
   U2669 : OAI22_X1 port map( A1 => n13876, A2 => n12171, B1 => n13710, B2 => 
                           n12165, ZN => n4078);
   U2670 : AOI221_X1 port map( B1 => n12279, B2 => n11663, C1 => n12273, C2 => 
                           n11483, A => n4051, ZN => n4046);
   U2671 : OAI22_X1 port map( A1 => n13533, A2 => n12267, B1 => n13473, B2 => 
                           n12261, ZN => n4051);
   U2672 : AOI221_X1 port map( B1 => n12183, B2 => n14062, C1 => n12177, C2 => 
                           n14109, A => n4059, ZN => n4054);
   U2673 : OAI22_X1 port map( A1 => n13875, A2 => n12171, B1 => n13709, B2 => 
                           n12165, ZN => n4059);
   U2674 : AOI221_X1 port map( B1 => n12279, B2 => n11664, C1 => n12273, C2 => 
                           n11484, A => n4032, ZN => n4027);
   U2675 : OAI22_X1 port map( A1 => n13532, A2 => n12267, B1 => n13472, B2 => 
                           n12261, ZN => n4032);
   U2676 : AOI221_X1 port map( B1 => n12183, B2 => n14061, C1 => n12177, C2 => 
                           n14108, A => n4040, ZN => n4035);
   U2677 : OAI22_X1 port map( A1 => n13874, A2 => n12171, B1 => n13708, B2 => 
                           n12165, ZN => n4040);
   U2678 : AOI221_X1 port map( B1 => n12279, B2 => n11665, C1 => n12273, C2 => 
                           n11485, A => n4013, ZN => n4008);
   U2679 : OAI22_X1 port map( A1 => n13531, A2 => n12267, B1 => n13471, B2 => 
                           n12261, ZN => n4013);
   U2680 : AOI221_X1 port map( B1 => n12183, B2 => n14060, C1 => n12177, C2 => 
                           n14107, A => n4021, ZN => n4016);
   U2681 : OAI22_X1 port map( A1 => n13873, A2 => n12171, B1 => n13707, B2 => 
                           n12165, ZN => n4021);
   U2682 : AOI221_X1 port map( B1 => n12280, B2 => n11666, C1 => n12274, C2 => 
                           n11486, A => n3994, ZN => n3989);
   U2683 : OAI22_X1 port map( A1 => n13530, A2 => n12268, B1 => n13470, B2 => 
                           n12262, ZN => n3994);
   U2684 : AOI221_X1 port map( B1 => n12184, B2 => n13928, C1 => n12178, C2 => 
                           n13988, A => n4002, ZN => n3997);
   U2685 : OAI22_X1 port map( A1 => n13872, A2 => n12172, B1 => n13706, B2 => 
                           n12166, ZN => n4002);
   U2686 : AOI221_X1 port map( B1 => n12280, B2 => n11667, C1 => n12274, C2 => 
                           n11487, A => n3975, ZN => n3970);
   U2687 : OAI22_X1 port map( A1 => n13529, A2 => n12268, B1 => n13469, B2 => 
                           n12262, ZN => n3975);
   U2688 : AOI221_X1 port map( B1 => n12184, B2 => n13927, C1 => n12178, C2 => 
                           n13987, A => n3983, ZN => n3978);
   U2689 : OAI22_X1 port map( A1 => n13871, A2 => n12172, B1 => n13705, B2 => 
                           n12166, ZN => n3983);
   U2690 : AOI221_X1 port map( B1 => n12280, B2 => n11668, C1 => n12274, C2 => 
                           n11488, A => n3956, ZN => n3951);
   U2691 : OAI22_X1 port map( A1 => n13528, A2 => n12268, B1 => n13468, B2 => 
                           n12262, ZN => n3956);
   U2692 : AOI221_X1 port map( B1 => n12184, B2 => n13926, C1 => n12178, C2 => 
                           n13986, A => n3964, ZN => n3959);
   U2693 : OAI22_X1 port map( A1 => n13870, A2 => n12172, B1 => n13704, B2 => 
                           n12166, ZN => n3964);
   U2694 : AOI221_X1 port map( B1 => n12280, B2 => n11669, C1 => n12274, C2 => 
                           n11489, A => n3937, ZN => n3932);
   U2695 : OAI22_X1 port map( A1 => n13527, A2 => n12268, B1 => n13467, B2 => 
                           n12262, ZN => n3937);
   U2696 : AOI221_X1 port map( B1 => n12184, B2 => n13925, C1 => n12178, C2 => 
                           n13985, A => n3945, ZN => n3940);
   U2697 : OAI22_X1 port map( A1 => n13869, A2 => n12172, B1 => n13703, B2 => 
                           n12166, ZN => n3945);
   U2698 : AOI221_X1 port map( B1 => n12280, B2 => n11670, C1 => n12274, C2 => 
                           n11490, A => n3918, ZN => n3913);
   U2699 : OAI22_X1 port map( A1 => n13526, A2 => n12268, B1 => n13466, B2 => 
                           n12262, ZN => n3918);
   U2700 : AOI221_X1 port map( B1 => n12184, B2 => n13924, C1 => n12178, C2 => 
                           n13984, A => n3926, ZN => n3921);
   U2701 : OAI22_X1 port map( A1 => n14059, A2 => n12172, B1 => n13702, B2 => 
                           n12166, ZN => n3926);
   U2702 : AOI221_X1 port map( B1 => n12280, B2 => n11671, C1 => n12274, C2 => 
                           n11491, A => n3899, ZN => n3894);
   U2703 : OAI22_X1 port map( A1 => n13525, A2 => n12268, B1 => n13465, B2 => 
                           n12262, ZN => n3899);
   U2704 : AOI221_X1 port map( B1 => n12184, B2 => n13923, C1 => n12178, C2 => 
                           n13983, A => n3907, ZN => n3902);
   U2705 : OAI22_X1 port map( A1 => n14058, A2 => n12172, B1 => n13701, B2 => 
                           n12166, ZN => n3907);
   U2706 : AOI221_X1 port map( B1 => n12280, B2 => n11672, C1 => n12274, C2 => 
                           n11492, A => n3880, ZN => n3875);
   U2707 : OAI22_X1 port map( A1 => n13524, A2 => n12268, B1 => n13464, B2 => 
                           n12262, ZN => n3880);
   U2708 : AOI221_X1 port map( B1 => n12184, B2 => n13922, C1 => n12178, C2 => 
                           n13982, A => n3888, ZN => n3883);
   U2709 : OAI22_X1 port map( A1 => n14057, A2 => n12172, B1 => n13700, B2 => 
                           n12166, ZN => n3888);
   U2710 : AOI221_X1 port map( B1 => n12280, B2 => n11673, C1 => n12274, C2 => 
                           n11493, A => n3861, ZN => n3856);
   U2711 : OAI22_X1 port map( A1 => n13523, A2 => n12268, B1 => n13463, B2 => 
                           n12262, ZN => n3861);
   U2712 : AOI221_X1 port map( B1 => n12184, B2 => n13921, C1 => n12178, C2 => 
                           n13981, A => n3869, ZN => n3864);
   U2713 : OAI22_X1 port map( A1 => n14056, A2 => n12172, B1 => n13699, B2 => 
                           n12166, ZN => n3869);
   U2714 : AOI221_X1 port map( B1 => n12280, B2 => n11674, C1 => n12274, C2 => 
                           n11494, A => n3842, ZN => n3837);
   U2715 : OAI22_X1 port map( A1 => n13522, A2 => n12268, B1 => n13462, B2 => 
                           n12262, ZN => n3842);
   U2716 : AOI221_X1 port map( B1 => n12184, B2 => n13920, C1 => n12178, C2 => 
                           n13980, A => n3850, ZN => n3845);
   U2717 : OAI22_X1 port map( A1 => n14055, A2 => n12172, B1 => n13698, B2 => 
                           n12166, ZN => n3850);
   U2718 : AOI221_X1 port map( B1 => n12280, B2 => n11675, C1 => n12274, C2 => 
                           n11495, A => n3823, ZN => n3818);
   U2719 : OAI22_X1 port map( A1 => n13521, A2 => n12268, B1 => n13461, B2 => 
                           n12262, ZN => n3823);
   U2720 : AOI221_X1 port map( B1 => n12184, B2 => n13919, C1 => n12178, C2 => 
                           n13979, A => n3831, ZN => n3826);
   U2721 : OAI22_X1 port map( A1 => n14054, A2 => n12172, B1 => n13697, B2 => 
                           n12166, ZN => n3831);
   U2722 : AOI221_X1 port map( B1 => n12280, B2 => n11676, C1 => n12274, C2 => 
                           n11496, A => n3804, ZN => n3799);
   U2723 : OAI22_X1 port map( A1 => n13520, A2 => n12268, B1 => n13460, B2 => 
                           n12262, ZN => n3804);
   U2724 : AOI221_X1 port map( B1 => n12184, B2 => n13918, C1 => n12178, C2 => 
                           n13978, A => n3812, ZN => n3807);
   U2725 : OAI22_X1 port map( A1 => n14053, A2 => n12172, B1 => n13696, B2 => 
                           n12166, ZN => n3812);
   U2726 : AOI221_X1 port map( B1 => n12280, B2 => n11677, C1 => n12274, C2 => 
                           n11497, A => n3785, ZN => n3780);
   U2727 : OAI22_X1 port map( A1 => n13519, A2 => n12268, B1 => n13459, B2 => 
                           n12262, ZN => n3785);
   U2728 : AOI221_X1 port map( B1 => n12184, B2 => n13917, C1 => n12178, C2 => 
                           n13977, A => n3793, ZN => n3788);
   U2729 : OAI22_X1 port map( A1 => n14052, A2 => n12172, B1 => n13695, B2 => 
                           n12166, ZN => n3793);
   U2730 : AOI221_X1 port map( B1 => n12281, B2 => n11678, C1 => n12275, C2 => 
                           n11498, A => n3766, ZN => n3761);
   U2731 : OAI22_X1 port map( A1 => n13518, A2 => n12269, B1 => n13458, B2 => 
                           n12263, ZN => n3766);
   U2732 : AOI221_X1 port map( B1 => n12185, B2 => n13916, C1 => n12179, C2 => 
                           n13976, A => n3774, ZN => n3769);
   U2733 : OAI22_X1 port map( A1 => n14051, A2 => n12173, B1 => n13694, B2 => 
                           n12167, ZN => n3774);
   U2734 : AOI221_X1 port map( B1 => n12281, B2 => n11679, C1 => n12275, C2 => 
                           n11499, A => n3747, ZN => n3742);
   U2735 : OAI22_X1 port map( A1 => n13517, A2 => n12269, B1 => n13457, B2 => 
                           n12263, ZN => n3747);
   U2736 : AOI221_X1 port map( B1 => n12185, B2 => n13915, C1 => n12179, C2 => 
                           n13975, A => n3755, ZN => n3750);
   U2737 : OAI22_X1 port map( A1 => n14050, A2 => n12173, B1 => n13693, B2 => 
                           n12167, ZN => n3755);
   U2738 : AOI221_X1 port map( B1 => n12281, B2 => n11680, C1 => n12275, C2 => 
                           n11500, A => n3728, ZN => n3723);
   U2739 : OAI22_X1 port map( A1 => n13516, A2 => n12269, B1 => n13456, B2 => 
                           n12263, ZN => n3728);
   U2740 : AOI221_X1 port map( B1 => n12185, B2 => n13914, C1 => n12179, C2 => 
                           n13974, A => n3736, ZN => n3731);
   U2741 : OAI22_X1 port map( A1 => n14049, A2 => n12173, B1 => n13692, B2 => 
                           n12167, ZN => n3736);
   U2742 : AOI221_X1 port map( B1 => n12281, B2 => n11681, C1 => n12275, C2 => 
                           n11501, A => n3709, ZN => n3704);
   U2743 : OAI22_X1 port map( A1 => n14460, A2 => n12269, B1 => n13455, B2 => 
                           n12263, ZN => n3709);
   U2744 : AOI221_X1 port map( B1 => n12185, B2 => n13913, C1 => n12179, C2 => 
                           n13973, A => n3717, ZN => n3712);
   U2745 : OAI22_X1 port map( A1 => n14048, A2 => n12173, B1 => n13691, B2 => 
                           n12167, ZN => n3717);
   U2746 : AOI221_X1 port map( B1 => n12281, B2 => n11682, C1 => n12275, C2 => 
                           n11502, A => n3690, ZN => n3685);
   U2747 : OAI22_X1 port map( A1 => n14459, A2 => n12269, B1 => n13454, B2 => 
                           n12263, ZN => n3690);
   U2748 : AOI221_X1 port map( B1 => n12185, B2 => n13912, C1 => n12179, C2 => 
                           n13972, A => n3698, ZN => n3693);
   U2749 : OAI22_X1 port map( A1 => n14047, A2 => n12173, B1 => n13690, B2 => 
                           n12167, ZN => n3698);
   U2750 : AOI221_X1 port map( B1 => n12281, B2 => n11683, C1 => n12275, C2 => 
                           n11503, A => n3671, ZN => n3666);
   U2751 : OAI22_X1 port map( A1 => n14458, A2 => n12269, B1 => n13453, B2 => 
                           n12263, ZN => n3671);
   U2752 : AOI221_X1 port map( B1 => n12185, B2 => n13911, C1 => n12179, C2 => 
                           n13971, A => n3679, ZN => n3674);
   U2753 : OAI22_X1 port map( A1 => n14046, A2 => n12173, B1 => n13689, B2 => 
                           n12167, ZN => n3679);
   U2754 : AOI221_X1 port map( B1 => n12281, B2 => n11684, C1 => n12275, C2 => 
                           n11504, A => n3652, ZN => n3647);
   U2755 : OAI22_X1 port map( A1 => n14457, A2 => n12269, B1 => n13452, B2 => 
                           n12263, ZN => n3652);
   U2756 : AOI221_X1 port map( B1 => n12185, B2 => n13910, C1 => n12179, C2 => 
                           n13970, A => n3660, ZN => n3655);
   U2757 : OAI22_X1 port map( A1 => n14045, A2 => n12173, B1 => n13688, B2 => 
                           n12167, ZN => n3660);
   U2758 : AOI221_X1 port map( B1 => n12281, B2 => n11685, C1 => n12275, C2 => 
                           n11505, A => n3633, ZN => n3628);
   U2759 : OAI22_X1 port map( A1 => n13515, A2 => n12269, B1 => n13451, B2 => 
                           n12263, ZN => n3633);
   U2760 : AOI221_X1 port map( B1 => n12185, B2 => n13909, C1 => n12179, C2 => 
                           n13969, A => n3641, ZN => n3636);
   U2761 : OAI22_X1 port map( A1 => n14044, A2 => n12173, B1 => n13687, B2 => 
                           n12167, ZN => n3641);
   U2762 : AOI221_X1 port map( B1 => n12281, B2 => n11686, C1 => n12275, C2 => 
                           n11506, A => n3614, ZN => n3609);
   U2763 : OAI22_X1 port map( A1 => n13514, A2 => n12269, B1 => n13450, B2 => 
                           n12263, ZN => n3614);
   U2764 : AOI221_X1 port map( B1 => n12185, B2 => n13908, C1 => n12179, C2 => 
                           n13968, A => n3622, ZN => n3617);
   U2765 : OAI22_X1 port map( A1 => n14043, A2 => n12173, B1 => n13686, B2 => 
                           n12167, ZN => n3622);
   U2766 : AOI221_X1 port map( B1 => n12281, B2 => n11687, C1 => n12275, C2 => 
                           n11507, A => n3595, ZN => n3590);
   U2767 : OAI22_X1 port map( A1 => n13513, A2 => n12269, B1 => n13449, B2 => 
                           n12263, ZN => n3595);
   U2768 : AOI221_X1 port map( B1 => n12185, B2 => n13907, C1 => n12179, C2 => 
                           n13967, A => n3603, ZN => n3598);
   U2769 : OAI22_X1 port map( A1 => n14042, A2 => n12173, B1 => n13685, B2 => 
                           n12167, ZN => n3603);
   U2770 : AOI221_X1 port map( B1 => n12281, B2 => n11688, C1 => n12275, C2 => 
                           n11508, A => n3576, ZN => n3571);
   U2771 : OAI22_X1 port map( A1 => n13512, A2 => n12269, B1 => n13448, B2 => 
                           n12263, ZN => n3576);
   U2772 : AOI221_X1 port map( B1 => n12185, B2 => n13906, C1 => n12179, C2 => 
                           n13966, A => n3584, ZN => n3579);
   U2773 : OAI22_X1 port map( A1 => n14041, A2 => n12173, B1 => n13684, B2 => 
                           n12167, ZN => n3584);
   U2774 : AOI221_X1 port map( B1 => n12281, B2 => n11689, C1 => n12275, C2 => 
                           n11509, A => n3557, ZN => n3552);
   U2775 : OAI22_X1 port map( A1 => n13511, A2 => n12269, B1 => n13447, B2 => 
                           n12263, ZN => n3557);
   U2776 : AOI221_X1 port map( B1 => n12185, B2 => n13905, C1 => n12179, C2 => 
                           n13965, A => n3565, ZN => n3560);
   U2777 : OAI22_X1 port map( A1 => n14040, A2 => n12173, B1 => n13683, B2 => 
                           n12167, ZN => n3565);
   U2778 : AOI221_X1 port map( B1 => n12282, B2 => n11690, C1 => n12276, C2 => 
                           n11510, A => n3538, ZN => n3533);
   U2779 : OAI22_X1 port map( A1 => n13510, A2 => n12270, B1 => n13446, B2 => 
                           n12264, ZN => n3538);
   U2780 : AOI221_X1 port map( B1 => n12186, B2 => n13904, C1 => n12180, C2 => 
                           n13964, A => n3546, ZN => n3541);
   U2781 : OAI22_X1 port map( A1 => n14039, A2 => n12174, B1 => n13682, B2 => 
                           n12168, ZN => n3546);
   U2782 : AOI221_X1 port map( B1 => n12282, B2 => n11691, C1 => n12276, C2 => 
                           n11511, A => n3519, ZN => n3514);
   U2783 : OAI22_X1 port map( A1 => n13509, A2 => n12270, B1 => n13445, B2 => 
                           n12264, ZN => n3519);
   U2784 : AOI221_X1 port map( B1 => n12186, B2 => n13903, C1 => n12180, C2 => 
                           n13963, A => n3527, ZN => n3522);
   U2785 : OAI22_X1 port map( A1 => n14038, A2 => n12174, B1 => n13681, B2 => 
                           n12168, ZN => n3527);
   U2786 : AOI221_X1 port map( B1 => n12282, B2 => n11692, C1 => n12276, C2 => 
                           n11512, A => n3500, ZN => n3495);
   U2787 : OAI22_X1 port map( A1 => n13508, A2 => n12270, B1 => n13444, B2 => 
                           n12264, ZN => n3500);
   U2788 : AOI221_X1 port map( B1 => n12186, B2 => n13902, C1 => n12180, C2 => 
                           n13962, A => n3508, ZN => n3503);
   U2789 : OAI22_X1 port map( A1 => n14037, A2 => n12174, B1 => n13680, B2 => 
                           n12168, ZN => n3508);
   U2790 : AOI221_X1 port map( B1 => n12282, B2 => n11693, C1 => n12276, C2 => 
                           n11513, A => n3481, ZN => n3476);
   U2791 : OAI22_X1 port map( A1 => n13507, A2 => n12270, B1 => n13443, B2 => 
                           n12264, ZN => n3481);
   U2792 : AOI221_X1 port map( B1 => n12186, B2 => n13901, C1 => n12180, C2 => 
                           n13961, A => n3489, ZN => n3484);
   U2793 : OAI22_X1 port map( A1 => n14036, A2 => n12174, B1 => n13679, B2 => 
                           n12168, ZN => n3489);
   U2794 : AOI221_X1 port map( B1 => n12282, B2 => n11694, C1 => n12276, C2 => 
                           n11514, A => n3462, ZN => n3457);
   U2795 : OAI22_X1 port map( A1 => n13506, A2 => n12270, B1 => n13442, B2 => 
                           n12264, ZN => n3462);
   U2796 : AOI221_X1 port map( B1 => n12186, B2 => n13900, C1 => n12180, C2 => 
                           n13960, A => n3470, ZN => n3465);
   U2797 : OAI22_X1 port map( A1 => n13742, A2 => n12174, B1 => n13678, B2 => 
                           n12168, ZN => n3470);
   U2798 : AOI221_X1 port map( B1 => n12282, B2 => n11695, C1 => n12276, C2 => 
                           n11515, A => n3443, ZN => n3438);
   U2799 : OAI22_X1 port map( A1 => n13505, A2 => n12270, B1 => n13441, B2 => 
                           n12264, ZN => n3443);
   U2800 : AOI221_X1 port map( B1 => n12186, B2 => n13899, C1 => n12180, C2 => 
                           n13959, A => n3451, ZN => n3446);
   U2801 : OAI22_X1 port map( A1 => n13741, A2 => n12174, B1 => n13677, B2 => 
                           n12168, ZN => n3451);
   U2802 : AOI221_X1 port map( B1 => n12282, B2 => n11696, C1 => n12276, C2 => 
                           n11516, A => n3424, ZN => n3419);
   U2803 : OAI22_X1 port map( A1 => n13504, A2 => n12270, B1 => n13440, B2 => 
                           n12264, ZN => n3424);
   U2804 : AOI221_X1 port map( B1 => n12186, B2 => n13898, C1 => n12180, C2 => 
                           n13958, A => n3432, ZN => n3427);
   U2805 : OAI22_X1 port map( A1 => n13740, A2 => n12174, B1 => n13676, B2 => 
                           n12168, ZN => n3432);
   U2806 : AOI221_X1 port map( B1 => n12282, B2 => n11697, C1 => n12276, C2 => 
                           n11517, A => n3405, ZN => n3400);
   U2807 : OAI22_X1 port map( A1 => n13503, A2 => n12270, B1 => n13439, B2 => 
                           n12264, ZN => n3405);
   U2808 : AOI221_X1 port map( B1 => n12186, B2 => n13897, C1 => n12180, C2 => 
                           n13957, A => n3413, ZN => n3408);
   U2809 : OAI22_X1 port map( A1 => n13739, A2 => n12174, B1 => n13675, B2 => 
                           n12168, ZN => n3413);
   U2810 : AOI221_X1 port map( B1 => n12282, B2 => n11698, C1 => n12276, C2 => 
                           n11518, A => n3386, ZN => n3381);
   U2811 : OAI22_X1 port map( A1 => n13502, A2 => n12270, B1 => n13438, B2 => 
                           n12264, ZN => n3386);
   U2812 : AOI221_X1 port map( B1 => n12186, B2 => n13896, C1 => n12180, C2 => 
                           n13956, A => n3394, ZN => n3389);
   U2813 : OAI22_X1 port map( A1 => n13738, A2 => n12174, B1 => n13674, B2 => 
                           n12168, ZN => n3394);
   U2814 : AOI221_X1 port map( B1 => n12282, B2 => n11699, C1 => n12276, C2 => 
                           n11519, A => n3367, ZN => n3362);
   U2815 : OAI22_X1 port map( A1 => n13501, A2 => n12270, B1 => n13437, B2 => 
                           n12264, ZN => n3367);
   U2816 : AOI221_X1 port map( B1 => n12186, B2 => n13895, C1 => n12180, C2 => 
                           n13955, A => n3375, ZN => n3370);
   U2817 : OAI22_X1 port map( A1 => n13737, A2 => n12174, B1 => n13673, B2 => 
                           n12168, ZN => n3375);
   U2818 : AOI221_X1 port map( B1 => n12282, B2 => n11700, C1 => n12276, C2 => 
                           n11520, A => n3348, ZN => n3343);
   U2819 : OAI22_X1 port map( A1 => n13500, A2 => n12270, B1 => n13436, B2 => 
                           n12264, ZN => n3348);
   U2820 : AOI221_X1 port map( B1 => n12186, B2 => n13894, C1 => n12180, C2 => 
                           n13954, A => n3356, ZN => n3351);
   U2821 : OAI22_X1 port map( A1 => n13736, A2 => n12174, B1 => n13672, B2 => 
                           n12168, ZN => n3356);
   U2822 : AOI221_X1 port map( B1 => n12282, B2 => n11701, C1 => n12276, C2 => 
                           n11521, A => n3329, ZN => n3324);
   U2823 : OAI22_X1 port map( A1 => n13499, A2 => n12270, B1 => n13435, B2 => 
                           n12264, ZN => n3329);
   U2824 : AOI221_X1 port map( B1 => n12186, B2 => n13893, C1 => n12180, C2 => 
                           n13953, A => n3337, ZN => n3332);
   U2825 : OAI22_X1 port map( A1 => n13735, A2 => n12174, B1 => n13671, B2 => 
                           n12168, ZN => n3337);
   U2826 : AOI221_X1 port map( B1 => n12187, B2 => n13819, C1 => n12181, C2 => 
                           n13823, A => n3318, ZN => n3313);
   U2827 : OAI22_X1 port map( A1 => n13734, A2 => n12175, B1 => n13670, B2 => 
                           n12169, ZN => n3318);
   U2828 : AOI221_X1 port map( B1 => n12283, B2 => n13860, C1 => n12277, C2 => 
                           n13856, A => n3310, ZN => n3305);
   U2829 : OAI22_X1 port map( A1 => n13498, A2 => n12271, B1 => n13434, B2 => 
                           n12265, ZN => n3310);
   U2830 : AOI221_X1 port map( B1 => n12187, B2 => n13818, C1 => n12181, C2 => 
                           n13822, A => n3299, ZN => n3294);
   U2831 : OAI22_X1 port map( A1 => n13733, A2 => n12175, B1 => n13669, B2 => 
                           n12169, ZN => n3299);
   U2832 : AOI221_X1 port map( B1 => n12283, B2 => n13859, C1 => n12277, C2 => 
                           n13855, A => n3291, ZN => n3286);
   U2833 : OAI22_X1 port map( A1 => n13497, A2 => n12271, B1 => n13433, B2 => 
                           n12265, ZN => n3291);
   U2834 : AOI221_X1 port map( B1 => n12187, B2 => n13817, C1 => n12181, C2 => 
                           n13821, A => n3280, ZN => n3275);
   U2835 : OAI22_X1 port map( A1 => n13732, A2 => n12175, B1 => n13668, B2 => 
                           n12169, ZN => n3280);
   U2836 : AOI221_X1 port map( B1 => n12283, B2 => n13858, C1 => n12277, C2 => 
                           n13854, A => n3272, ZN => n3267);
   U2837 : OAI22_X1 port map( A1 => n13496, A2 => n12271, B1 => n13432, B2 => 
                           n12265, ZN => n3272);
   U2838 : AOI221_X1 port map( B1 => n12187, B2 => n13816, C1 => n12181, C2 => 
                           n13820, A => n3255, ZN => n3240);
   U2839 : OAI22_X1 port map( A1 => n13731, A2 => n12175, B1 => n13667, B2 => 
                           n12169, ZN => n3255);
   U2840 : AOI221_X1 port map( B1 => n12283, B2 => n13857, C1 => n12277, C2 => 
                           n13853, A => n3231, ZN => n3216);
   U2841 : OAI22_X1 port map( A1 => n13495, A2 => n12271, B1 => n13431, B2 => 
                           n12265, ZN => n3231);
   U2842 : AOI221_X1 port map( B1 => n12254, B2 => n11702, C1 => n12248, C2 => 
                           n11522, A => n4459, ZN => n4444);
   U2843 : OAI22_X1 port map( A1 => n13650, A2 => n12242, B1 => n13603, B2 => 
                           n12236, ZN => n4459);
   U2844 : AOI221_X1 port map( B1 => n12158, B2 => n14155, C1 => n12152, C2 => 
                           n13831, A => n4471, ZN => n4460);
   U2845 : OAI22_X1 port map( A1 => n13815, A2 => n12146, B1 => n13810, B2 => 
                           n12140, ZN => n4471);
   U2846 : AOI221_X1 port map( B1 => n12254, B2 => n11703, C1 => n12248, C2 => 
                           n11523, A => n4432, ZN => n4425);
   U2847 : OAI22_X1 port map( A1 => n13649, A2 => n12242, B1 => n13602, B2 => 
                           n12236, ZN => n4432);
   U2848 : AOI221_X1 port map( B1 => n12158, B2 => n14152, C1 => n12152, C2 => 
                           n13830, A => n4440, ZN => n4433);
   U2849 : OAI22_X1 port map( A1 => n13814, A2 => n12146, B1 => n13809, B2 => 
                           n12140, ZN => n4440);
   U2850 : AOI221_X1 port map( B1 => n12254, B2 => n11704, C1 => n12248, C2 => 
                           n11524, A => n4413, ZN => n4406);
   U2851 : OAI22_X1 port map( A1 => n13648, A2 => n12242, B1 => n13601, B2 => 
                           n12236, ZN => n4413);
   U2852 : AOI221_X1 port map( B1 => n12158, B2 => n14151, C1 => n12152, C2 => 
                           n13829, A => n4421, ZN => n4414);
   U2853 : OAI22_X1 port map( A1 => n13813, A2 => n12146, B1 => n13808, B2 => 
                           n12140, ZN => n4421);
   U2854 : AOI221_X1 port map( B1 => n12254, B2 => n11705, C1 => n12248, C2 => 
                           n11525, A => n4394, ZN => n4387);
   U2855 : OAI22_X1 port map( A1 => n13647, A2 => n12242, B1 => n13600, B2 => 
                           n12236, ZN => n4394);
   U2856 : AOI221_X1 port map( B1 => n12158, B2 => n14149, C1 => n12152, C2 => 
                           n13828, A => n4402, ZN => n4395);
   U2857 : OAI22_X1 port map( A1 => n13812, A2 => n12146, B1 => n13807, B2 => 
                           n12140, ZN => n4402);
   U2858 : AOI221_X1 port map( B1 => n12254, B2 => n11706, C1 => n12248, C2 => 
                           n11526, A => n4375, ZN => n4368);
   U2859 : OAI22_X1 port map( A1 => n14357, A2 => n12242, B1 => n13599, B2 => 
                           n12236, ZN => n4375);
   U2860 : AOI221_X1 port map( B1 => n12158, B2 => n14150, C1 => n12152, C2 => 
                           n14215, A => n4383, ZN => n4376);
   U2861 : OAI22_X1 port map( A1 => n13811, A2 => n12146, B1 => n13806, B2 => 
                           n12140, ZN => n4383);
   U2862 : AOI221_X1 port map( B1 => n12254, B2 => n11707, C1 => n12248, C2 => 
                           n11527, A => n4356, ZN => n4349);
   U2863 : OAI22_X1 port map( A1 => n14356, A2 => n12242, B1 => n13598, B2 => 
                           n12236, ZN => n4356);
   U2864 : AOI221_X1 port map( B1 => n12158, B2 => n14148, C1 => n12152, C2 => 
                           n14214, A => n4364, ZN => n4357);
   U2865 : OAI22_X1 port map( A1 => n14035, A2 => n12146, B1 => n13805, B2 => 
                           n12140, ZN => n4364);
   U2866 : AOI221_X1 port map( B1 => n12254, B2 => n11708, C1 => n12248, C2 => 
                           n11528, A => n4337, ZN => n4330);
   U2867 : OAI22_X1 port map( A1 => n14355, A2 => n12242, B1 => n13597, B2 => 
                           n12236, ZN => n4337);
   U2868 : AOI221_X1 port map( B1 => n12158, B2 => n14147, C1 => n12152, C2 => 
                           n14213, A => n4345, ZN => n4338);
   U2869 : OAI22_X1 port map( A1 => n14034, A2 => n12146, B1 => n13804, B2 => 
                           n12140, ZN => n4345);
   U2870 : AOI221_X1 port map( B1 => n12254, B2 => n11709, C1 => n12248, C2 => 
                           n11529, A => n4318, ZN => n4311);
   U2871 : OAI22_X1 port map( A1 => n14354, A2 => n12242, B1 => n13596, B2 => 
                           n12236, ZN => n4318);
   U2872 : AOI221_X1 port map( B1 => n12158, B2 => n14146, C1 => n12152, C2 => 
                           n14212, A => n4326, ZN => n4319);
   U2873 : OAI22_X1 port map( A1 => n14033, A2 => n12146, B1 => n13803, B2 => 
                           n12140, ZN => n4326);
   U2874 : AOI221_X1 port map( B1 => n12254, B2 => n11710, C1 => n12248, C2 => 
                           n11530, A => n4299, ZN => n4292);
   U2875 : OAI22_X1 port map( A1 => n14353, A2 => n12242, B1 => n13595, B2 => 
                           n12236, ZN => n4299);
   U2876 : AOI221_X1 port map( B1 => n12158, B2 => n14145, C1 => n12152, C2 => 
                           n14211, A => n4307, ZN => n4300);
   U2877 : OAI22_X1 port map( A1 => n14032, A2 => n12146, B1 => n13802, B2 => 
                           n12140, ZN => n4307);
   U2878 : AOI221_X1 port map( B1 => n12254, B2 => n11711, C1 => n12248, C2 => 
                           n11531, A => n4280, ZN => n4273);
   U2879 : OAI22_X1 port map( A1 => n14352, A2 => n12242, B1 => n13594, B2 => 
                           n12236, ZN => n4280);
   U2880 : AOI221_X1 port map( B1 => n12158, B2 => n14144, C1 => n12152, C2 => 
                           n14210, A => n4288, ZN => n4281);
   U2881 : OAI22_X1 port map( A1 => n14031, A2 => n12146, B1 => n13801, B2 => 
                           n12140, ZN => n4288);
   U2882 : AOI221_X1 port map( B1 => n12254, B2 => n11712, C1 => n12248, C2 => 
                           n11532, A => n4261, ZN => n4254);
   U2883 : OAI22_X1 port map( A1 => n14351, A2 => n12242, B1 => n13593, B2 => 
                           n12236, ZN => n4261);
   U2884 : AOI221_X1 port map( B1 => n12158, B2 => n14143, C1 => n12152, C2 => 
                           n14209, A => n4269, ZN => n4262);
   U2885 : OAI22_X1 port map( A1 => n14030, A2 => n12146, B1 => n13800, B2 => 
                           n12140, ZN => n4269);
   U2886 : AOI221_X1 port map( B1 => n12254, B2 => n11713, C1 => n12248, C2 => 
                           n11533, A => n4242, ZN => n4235);
   U2887 : OAI22_X1 port map( A1 => n14350, A2 => n12242, B1 => n13592, B2 => 
                           n12236, ZN => n4242);
   U2888 : AOI221_X1 port map( B1 => n12158, B2 => n14142, C1 => n12152, C2 => 
                           n14208, A => n4250, ZN => n4243);
   U2889 : OAI22_X1 port map( A1 => n14029, A2 => n12146, B1 => n13799, B2 => 
                           n12140, ZN => n4250);
   U2890 : AOI221_X1 port map( B1 => n12255, B2 => n11714, C1 => n12249, C2 => 
                           n11534, A => n4223, ZN => n4216);
   U2891 : OAI22_X1 port map( A1 => n14349, A2 => n12243, B1 => n13591, B2 => 
                           n12237, ZN => n4223);
   U2892 : AOI221_X1 port map( B1 => n12159, B2 => n14141, C1 => n12153, C2 => 
                           n14207, A => n4231, ZN => n4224);
   U2893 : OAI22_X1 port map( A1 => n14028, A2 => n12147, B1 => n13798, B2 => 
                           n12141, ZN => n4231);
   U2894 : AOI221_X1 port map( B1 => n12255, B2 => n11715, C1 => n12249, C2 => 
                           n11535, A => n4204, ZN => n4197);
   U2895 : OAI22_X1 port map( A1 => n14348, A2 => n12243, B1 => n13590, B2 => 
                           n12237, ZN => n4204);
   U2896 : AOI221_X1 port map( B1 => n12159, B2 => n14140, C1 => n12153, C2 => 
                           n14206, A => n4212, ZN => n4205);
   U2897 : OAI22_X1 port map( A1 => n14027, A2 => n12147, B1 => n13797, B2 => 
                           n12141, ZN => n4212);
   U2898 : AOI221_X1 port map( B1 => n12255, B2 => n11716, C1 => n12249, C2 => 
                           n11536, A => n4185, ZN => n4178);
   U2899 : OAI22_X1 port map( A1 => n14347, A2 => n12243, B1 => n13589, B2 => 
                           n12237, ZN => n4185);
   U2900 : AOI221_X1 port map( B1 => n12159, B2 => n14139, C1 => n12153, C2 => 
                           n14205, A => n4193, ZN => n4186);
   U2901 : OAI22_X1 port map( A1 => n14026, A2 => n12147, B1 => n13796, B2 => 
                           n12141, ZN => n4193);
   U2902 : AOI221_X1 port map( B1 => n12255, B2 => n11717, C1 => n12249, C2 => 
                           n11537, A => n4166, ZN => n4159);
   U2903 : OAI22_X1 port map( A1 => n14346, A2 => n12243, B1 => n13588, B2 => 
                           n12237, ZN => n4166);
   U2904 : AOI221_X1 port map( B1 => n12159, B2 => n14138, C1 => n12153, C2 => 
                           n14204, A => n4174, ZN => n4167);
   U2905 : OAI22_X1 port map( A1 => n14025, A2 => n12147, B1 => n13795, B2 => 
                           n12141, ZN => n4174);
   U2906 : AOI221_X1 port map( B1 => n12255, B2 => n11718, C1 => n12249, C2 => 
                           n11538, A => n4147, ZN => n4140);
   U2907 : OAI22_X1 port map( A1 => n13646, A2 => n12243, B1 => n13587, B2 => 
                           n12237, ZN => n4147);
   U2908 : AOI221_X1 port map( B1 => n12159, B2 => n14137, C1 => n12153, C2 => 
                           n14203, A => n4155, ZN => n4148);
   U2909 : OAI22_X1 port map( A1 => n13952, A2 => n12147, B1 => n13794, B2 => 
                           n12141, ZN => n4155);
   U2910 : AOI221_X1 port map( B1 => n12255, B2 => n11719, C1 => n12249, C2 => 
                           n11539, A => n4128, ZN => n4121);
   U2911 : OAI22_X1 port map( A1 => n14345, A2 => n12243, B1 => n13586, B2 => 
                           n12237, ZN => n4128);
   U2912 : AOI221_X1 port map( B1 => n12159, B2 => n14136, C1 => n12153, C2 => 
                           n14202, A => n4136, ZN => n4129);
   U2913 : OAI22_X1 port map( A1 => n13951, A2 => n12147, B1 => n13793, B2 => 
                           n12141, ZN => n4136);
   U2914 : AOI221_X1 port map( B1 => n12255, B2 => n11720, C1 => n12249, C2 => 
                           n11540, A => n4109, ZN => n4102);
   U2915 : OAI22_X1 port map( A1 => n14344, A2 => n12243, B1 => n13585, B2 => 
                           n12237, ZN => n4109);
   U2916 : AOI221_X1 port map( B1 => n12159, B2 => n14135, C1 => n12153, C2 => 
                           n14201, A => n4117, ZN => n4110);
   U2917 : OAI22_X1 port map( A1 => n13950, A2 => n12147, B1 => n13792, B2 => 
                           n12141, ZN => n4117);
   U2918 : AOI221_X1 port map( B1 => n12255, B2 => n11721, C1 => n12249, C2 => 
                           n11541, A => n4090, ZN => n4083);
   U2919 : OAI22_X1 port map( A1 => n14343, A2 => n12243, B1 => n13584, B2 => 
                           n12237, ZN => n4090);
   U2920 : AOI221_X1 port map( B1 => n12159, B2 => n14134, C1 => n12153, C2 => 
                           n14200, A => n4098, ZN => n4091);
   U2921 : OAI22_X1 port map( A1 => n13949, A2 => n12147, B1 => n13791, B2 => 
                           n12141, ZN => n4098);
   U2922 : AOI221_X1 port map( B1 => n12255, B2 => n11722, C1 => n12249, C2 => 
                           n11542, A => n4071, ZN => n4064);
   U2923 : OAI22_X1 port map( A1 => n14342, A2 => n12243, B1 => n13583, B2 => 
                           n12237, ZN => n4071);
   U2924 : AOI221_X1 port map( B1 => n12159, B2 => n14133, C1 => n12153, C2 => 
                           n14199, A => n4079, ZN => n4072);
   U2925 : OAI22_X1 port map( A1 => n13948, A2 => n12147, B1 => n13790, B2 => 
                           n12141, ZN => n4079);
   U2926 : AOI221_X1 port map( B1 => n12255, B2 => n11723, C1 => n12249, C2 => 
                           n11543, A => n4052, ZN => n4045);
   U2927 : OAI22_X1 port map( A1 => n14341, A2 => n12243, B1 => n13582, B2 => 
                           n12237, ZN => n4052);
   U2928 : AOI221_X1 port map( B1 => n12159, B2 => n14132, C1 => n12153, C2 => 
                           n14198, A => n4060, ZN => n4053);
   U2929 : OAI22_X1 port map( A1 => n13947, A2 => n12147, B1 => n13789, B2 => 
                           n12141, ZN => n4060);
   U2930 : AOI221_X1 port map( B1 => n12255, B2 => n11724, C1 => n12249, C2 => 
                           n11544, A => n4033, ZN => n4026);
   U2931 : OAI22_X1 port map( A1 => n13645, A2 => n12243, B1 => n13581, B2 => 
                           n12237, ZN => n4033);
   U2932 : AOI221_X1 port map( B1 => n12159, B2 => n14131, C1 => n12153, C2 => 
                           n14197, A => n4041, ZN => n4034);
   U2933 : OAI22_X1 port map( A1 => n13946, A2 => n12147, B1 => n13788, B2 => 
                           n12141, ZN => n4041);
   U2934 : AOI221_X1 port map( B1 => n12255, B2 => n11725, C1 => n12249, C2 => 
                           n11545, A => n4014, ZN => n4007);
   U2935 : OAI22_X1 port map( A1 => n13644, A2 => n12243, B1 => n13580, B2 => 
                           n12237, ZN => n4014);
   U2936 : AOI221_X1 port map( B1 => n12159, B2 => n14130, C1 => n12153, C2 => 
                           n14196, A => n4022, ZN => n4015);
   U2937 : OAI22_X1 port map( A1 => n13945, A2 => n12147, B1 => n13787, B2 => 
                           n12141, ZN => n4022);
   U2938 : AOI221_X1 port map( B1 => n12256, B2 => n11726, C1 => n12250, C2 => 
                           n11546, A => n3995, ZN => n3988);
   U2939 : OAI22_X1 port map( A1 => n13643, A2 => n12244, B1 => n13579, B2 => 
                           n12238, ZN => n3995);
   U2940 : AOI221_X1 port map( B1 => n12160, B2 => n14024, C1 => n12154, C2 => 
                           n14195, A => n4003, ZN => n3996);
   U2941 : OAI22_X1 port map( A1 => n13944, A2 => n12148, B1 => n13786, B2 => 
                           n12142, ZN => n4003);
   U2942 : AOI221_X1 port map( B1 => n12256, B2 => n11727, C1 => n12250, C2 => 
                           n11547, A => n3976, ZN => n3969);
   U2943 : OAI22_X1 port map( A1 => n13642, A2 => n12244, B1 => n13578, B2 => 
                           n12238, ZN => n3976);
   U2944 : AOI221_X1 port map( B1 => n12160, B2 => n14023, C1 => n12154, C2 => 
                           n14194, A => n3984, ZN => n3977);
   U2945 : OAI22_X1 port map( A1 => n13943, A2 => n12148, B1 => n13785, B2 => 
                           n12142, ZN => n3984);
   U2946 : AOI221_X1 port map( B1 => n12256, B2 => n11728, C1 => n12250, C2 => 
                           n11548, A => n3957, ZN => n3950);
   U2947 : OAI22_X1 port map( A1 => n13641, A2 => n12244, B1 => n13577, B2 => 
                           n12238, ZN => n3957);
   U2948 : AOI221_X1 port map( B1 => n12160, B2 => n14022, C1 => n12154, C2 => 
                           n14193, A => n3965, ZN => n3958);
   U2949 : OAI22_X1 port map( A1 => n13942, A2 => n12148, B1 => n13784, B2 => 
                           n12142, ZN => n3965);
   U2950 : AOI221_X1 port map( B1 => n12256, B2 => n11729, C1 => n12250, C2 => 
                           n11549, A => n3938, ZN => n3931);
   U2951 : OAI22_X1 port map( A1 => n13640, A2 => n12244, B1 => n13576, B2 => 
                           n12238, ZN => n3938);
   U2952 : AOI221_X1 port map( B1 => n12160, B2 => n14021, C1 => n12154, C2 => 
                           n14192, A => n3946, ZN => n3939);
   U2953 : OAI22_X1 port map( A1 => n13941, A2 => n12148, B1 => n13783, B2 => 
                           n12142, ZN => n3946);
   U2954 : AOI221_X1 port map( B1 => n12256, B2 => n11730, C1 => n12250, C2 => 
                           n11550, A => n3919, ZN => n3912);
   U2955 : OAI22_X1 port map( A1 => n13639, A2 => n12244, B1 => n13575, B2 => 
                           n12238, ZN => n3919);
   U2956 : AOI221_X1 port map( B1 => n12160, B2 => n14020, C1 => n12154, C2 => 
                           n14191, A => n3927, ZN => n3920);
   U2957 : OAI22_X1 port map( A1 => n13940, A2 => n12148, B1 => n13782, B2 => 
                           n12142, ZN => n3927);
   U2958 : AOI221_X1 port map( B1 => n12256, B2 => n11731, C1 => n12250, C2 => 
                           n11551, A => n3900, ZN => n3893);
   U2959 : OAI22_X1 port map( A1 => n13638, A2 => n12244, B1 => n13574, B2 => 
                           n12238, ZN => n3900);
   U2960 : AOI221_X1 port map( B1 => n12160, B2 => n14019, C1 => n12154, C2 => 
                           n14190, A => n3908, ZN => n3901);
   U2961 : OAI22_X1 port map( A1 => n13939, A2 => n12148, B1 => n13781, B2 => 
                           n12142, ZN => n3908);
   U2962 : AOI221_X1 port map( B1 => n12256, B2 => n11732, C1 => n12250, C2 => 
                           n11552, A => n3881, ZN => n3874);
   U2963 : OAI22_X1 port map( A1 => n13637, A2 => n12244, B1 => n13573, B2 => 
                           n12238, ZN => n3881);
   U2964 : AOI221_X1 port map( B1 => n12160, B2 => n14018, C1 => n12154, C2 => 
                           n14189, A => n3889, ZN => n3882);
   U2965 : OAI22_X1 port map( A1 => n13938, A2 => n12148, B1 => n13780, B2 => 
                           n12142, ZN => n3889);
   U2966 : AOI221_X1 port map( B1 => n12256, B2 => n11733, C1 => n12250, C2 => 
                           n11553, A => n3862, ZN => n3855);
   U2967 : OAI22_X1 port map( A1 => n13636, A2 => n12244, B1 => n13572, B2 => 
                           n12238, ZN => n3862);
   U2968 : AOI221_X1 port map( B1 => n12160, B2 => n14017, C1 => n12154, C2 => 
                           n14188, A => n3870, ZN => n3863);
   U2969 : OAI22_X1 port map( A1 => n13937, A2 => n12148, B1 => n13779, B2 => 
                           n12142, ZN => n3870);
   U2970 : AOI221_X1 port map( B1 => n12256, B2 => n11734, C1 => n12250, C2 => 
                           n11554, A => n3843, ZN => n3836);
   U2971 : OAI22_X1 port map( A1 => n13635, A2 => n12244, B1 => n13571, B2 => 
                           n12238, ZN => n3843);
   U2972 : AOI221_X1 port map( B1 => n12160, B2 => n14016, C1 => n12154, C2 => 
                           n14187, A => n3851, ZN => n3844);
   U2973 : OAI22_X1 port map( A1 => n13936, A2 => n12148, B1 => n13778, B2 => 
                           n12142, ZN => n3851);
   U2974 : AOI221_X1 port map( B1 => n12256, B2 => n11735, C1 => n12250, C2 => 
                           n11555, A => n3824, ZN => n3817);
   U2975 : OAI22_X1 port map( A1 => n13634, A2 => n12244, B1 => n13570, B2 => 
                           n12238, ZN => n3824);
   U2976 : AOI221_X1 port map( B1 => n12160, B2 => n14015, C1 => n12154, C2 => 
                           n14186, A => n3832, ZN => n3825);
   U2977 : OAI22_X1 port map( A1 => n13935, A2 => n12148, B1 => n13777, B2 => 
                           n12142, ZN => n3832);
   U2978 : AOI221_X1 port map( B1 => n12256, B2 => n11736, C1 => n12250, C2 => 
                           n11556, A => n3805, ZN => n3798);
   U2979 : OAI22_X1 port map( A1 => n13633, A2 => n12244, B1 => n13569, B2 => 
                           n12238, ZN => n3805);
   U2980 : AOI221_X1 port map( B1 => n12160, B2 => n14014, C1 => n12154, C2 => 
                           n14185, A => n3813, ZN => n3806);
   U2981 : OAI22_X1 port map( A1 => n13934, A2 => n12148, B1 => n13776, B2 => 
                           n12142, ZN => n3813);
   U2982 : AOI221_X1 port map( B1 => n12256, B2 => n11737, C1 => n12250, C2 => 
                           n11557, A => n3786, ZN => n3779);
   U2983 : OAI22_X1 port map( A1 => n13632, A2 => n12244, B1 => n13568, B2 => 
                           n12238, ZN => n3786);
   U2984 : AOI221_X1 port map( B1 => n12160, B2 => n14013, C1 => n12154, C2 => 
                           n14184, A => n3794, ZN => n3787);
   U2985 : OAI22_X1 port map( A1 => n13933, A2 => n12148, B1 => n13775, B2 => 
                           n12142, ZN => n3794);
   U2986 : AOI221_X1 port map( B1 => n12257, B2 => n11738, C1 => n12251, C2 => 
                           n11558, A => n3767, ZN => n3760);
   U2987 : OAI22_X1 port map( A1 => n13631, A2 => n12245, B1 => n13567, B2 => 
                           n12239, ZN => n3767);
   U2988 : AOI221_X1 port map( B1 => n12161, B2 => n14012, C1 => n12155, C2 => 
                           n14183, A => n3775, ZN => n3768);
   U2989 : OAI22_X1 port map( A1 => n13932, A2 => n12149, B1 => n13774, B2 => 
                           n12143, ZN => n3775);
   U2990 : AOI221_X1 port map( B1 => n12257, B2 => n11739, C1 => n12251, C2 => 
                           n11559, A => n3748, ZN => n3741);
   U2991 : OAI22_X1 port map( A1 => n13630, A2 => n12245, B1 => n13566, B2 => 
                           n12239, ZN => n3748);
   U2992 : AOI221_X1 port map( B1 => n12161, B2 => n14011, C1 => n12155, C2 => 
                           n14182, A => n3756, ZN => n3749);
   U2993 : OAI22_X1 port map( A1 => n13931, A2 => n12149, B1 => n13773, B2 => 
                           n12143, ZN => n3756);
   U2994 : AOI221_X1 port map( B1 => n12257, B2 => n11740, C1 => n12251, C2 => 
                           n11560, A => n3729, ZN => n3722);
   U2995 : OAI22_X1 port map( A1 => n13629, A2 => n12245, B1 => n13565, B2 => 
                           n12239, ZN => n3729);
   U2996 : AOI221_X1 port map( B1 => n12161, B2 => n14010, C1 => n12155, C2 => 
                           n14181, A => n3737, ZN => n3730);
   U2997 : OAI22_X1 port map( A1 => n13930, A2 => n12149, B1 => n13772, B2 => 
                           n12143, ZN => n3737);
   U2998 : AOI221_X1 port map( B1 => n12257, B2 => n11741, C1 => n12251, C2 => 
                           n11561, A => n3710, ZN => n3703);
   U2999 : OAI22_X1 port map( A1 => n13628, A2 => n12245, B1 => n13564, B2 => 
                           n12239, ZN => n3710);
   U3000 : AOI221_X1 port map( B1 => n12161, B2 => n14009, C1 => n12155, C2 => 
                           n14180, A => n3718, ZN => n3711);
   U3001 : OAI22_X1 port map( A1 => n13929, A2 => n12149, B1 => n13771, B2 => 
                           n12143, ZN => n3718);
   U3002 : AOI221_X1 port map( B1 => n12257, B2 => n11742, C1 => n12251, C2 => 
                           n11562, A => n3691, ZN => n3684);
   U3003 : OAI22_X1 port map( A1 => n13627, A2 => n12245, B1 => n13563, B2 => 
                           n12239, ZN => n3691);
   U3004 : AOI221_X1 port map( B1 => n12161, B2 => n14008, C1 => n12155, C2 => 
                           n14179, A => n3699, ZN => n3692);
   U3005 : OAI22_X1 port map( A1 => n14106, A2 => n12149, B1 => n13770, B2 => 
                           n12143, ZN => n3699);
   U3006 : AOI221_X1 port map( B1 => n12257, B2 => n11743, C1 => n12251, C2 => 
                           n11563, A => n3672, ZN => n3665);
   U3007 : OAI22_X1 port map( A1 => n13626, A2 => n12245, B1 => n13562, B2 => 
                           n12239, ZN => n3672);
   U3008 : AOI221_X1 port map( B1 => n12161, B2 => n14007, C1 => n12155, C2 => 
                           n14178, A => n3680, ZN => n3673);
   U3009 : OAI22_X1 port map( A1 => n14105, A2 => n12149, B1 => n13769, B2 => 
                           n12143, ZN => n3680);
   U3010 : AOI221_X1 port map( B1 => n12257, B2 => n11744, C1 => n12251, C2 => 
                           n11564, A => n3653, ZN => n3646);
   U3011 : OAI22_X1 port map( A1 => n13625, A2 => n12245, B1 => n13561, B2 => 
                           n12239, ZN => n3653);
   U3012 : AOI221_X1 port map( B1 => n12161, B2 => n14006, C1 => n12155, C2 => 
                           n14177, A => n3661, ZN => n3654);
   U3013 : OAI22_X1 port map( A1 => n14104, A2 => n12149, B1 => n13768, B2 => 
                           n12143, ZN => n3661);
   U3014 : AOI221_X1 port map( B1 => n12257, B2 => n11745, C1 => n12251, C2 => 
                           n11565, A => n3634, ZN => n3627);
   U3015 : OAI22_X1 port map( A1 => n13624, A2 => n12245, B1 => n13560, B2 => 
                           n12239, ZN => n3634);
   U3016 : AOI221_X1 port map( B1 => n12161, B2 => n14005, C1 => n12155, C2 => 
                           n14176, A => n3642, ZN => n3635);
   U3017 : OAI22_X1 port map( A1 => n14103, A2 => n12149, B1 => n13767, B2 => 
                           n12143, ZN => n3642);
   U3018 : AOI221_X1 port map( B1 => n12257, B2 => n11746, C1 => n12251, C2 => 
                           n11566, A => n3615, ZN => n3608);
   U3019 : OAI22_X1 port map( A1 => n13623, A2 => n12245, B1 => n13559, B2 => 
                           n12239, ZN => n3615);
   U3020 : AOI221_X1 port map( B1 => n12161, B2 => n14004, C1 => n12155, C2 => 
                           n14175, A => n3623, ZN => n3616);
   U3021 : OAI22_X1 port map( A1 => n14102, A2 => n12149, B1 => n13766, B2 => 
                           n12143, ZN => n3623);
   U3022 : AOI221_X1 port map( B1 => n12257, B2 => n11747, C1 => n12251, C2 => 
                           n11567, A => n3596, ZN => n3589);
   U3023 : OAI22_X1 port map( A1 => n13622, A2 => n12245, B1 => n13558, B2 => 
                           n12239, ZN => n3596);
   U3024 : AOI221_X1 port map( B1 => n12161, B2 => n14003, C1 => n12155, C2 => 
                           n14174, A => n3604, ZN => n3597);
   U3025 : OAI22_X1 port map( A1 => n14101, A2 => n12149, B1 => n13765, B2 => 
                           n12143, ZN => n3604);
   U3026 : AOI221_X1 port map( B1 => n12257, B2 => n11748, C1 => n12251, C2 => 
                           n11568, A => n3577, ZN => n3570);
   U3027 : OAI22_X1 port map( A1 => n13621, A2 => n12245, B1 => n13557, B2 => 
                           n12239, ZN => n3577);
   U3028 : AOI221_X1 port map( B1 => n12161, B2 => n14002, C1 => n12155, C2 => 
                           n14173, A => n3585, ZN => n3578);
   U3029 : OAI22_X1 port map( A1 => n14100, A2 => n12149, B1 => n13764, B2 => 
                           n12143, ZN => n3585);
   U3030 : AOI221_X1 port map( B1 => n12257, B2 => n11749, C1 => n12251, C2 => 
                           n11569, A => n3558, ZN => n3551);
   U3031 : OAI22_X1 port map( A1 => n13620, A2 => n12245, B1 => n13556, B2 => 
                           n12239, ZN => n3558);
   U3032 : AOI221_X1 port map( B1 => n12161, B2 => n14001, C1 => n12155, C2 => 
                           n14172, A => n3566, ZN => n3559);
   U3033 : OAI22_X1 port map( A1 => n14099, A2 => n12149, B1 => n13763, B2 => 
                           n12143, ZN => n3566);
   U3034 : AOI221_X1 port map( B1 => n12258, B2 => n11750, C1 => n12252, C2 => 
                           n11570, A => n3539, ZN => n3532);
   U3035 : OAI22_X1 port map( A1 => n13619, A2 => n12246, B1 => n13555, B2 => 
                           n12240, ZN => n3539);
   U3036 : AOI221_X1 port map( B1 => n12162, B2 => n14000, C1 => n12156, C2 => 
                           n14171, A => n3547, ZN => n3540);
   U3037 : OAI22_X1 port map( A1 => n14098, A2 => n12150, B1 => n13762, B2 => 
                           n12144, ZN => n3547);
   U3038 : AOI221_X1 port map( B1 => n12258, B2 => n11751, C1 => n12252, C2 => 
                           n11571, A => n3520, ZN => n3513);
   U3039 : OAI22_X1 port map( A1 => n13618, A2 => n12246, B1 => n13554, B2 => 
                           n12240, ZN => n3520);
   U3040 : AOI221_X1 port map( B1 => n12162, B2 => n13999, C1 => n12156, C2 => 
                           n14170, A => n3528, ZN => n3521);
   U3041 : OAI22_X1 port map( A1 => n14097, A2 => n12150, B1 => n13761, B2 => 
                           n12144, ZN => n3528);
   U3042 : AOI221_X1 port map( B1 => n12258, B2 => n11752, C1 => n12252, C2 => 
                           n11572, A => n3501, ZN => n3494);
   U3043 : OAI22_X1 port map( A1 => n13617, A2 => n12246, B1 => n13553, B2 => 
                           n12240, ZN => n3501);
   U3044 : AOI221_X1 port map( B1 => n12162, B2 => n13998, C1 => n12156, C2 => 
                           n14169, A => n3509, ZN => n3502);
   U3045 : OAI22_X1 port map( A1 => n14096, A2 => n12150, B1 => n13760, B2 => 
                           n12144, ZN => n3509);
   U3046 : AOI221_X1 port map( B1 => n12258, B2 => n11753, C1 => n12252, C2 => 
                           n11573, A => n3482, ZN => n3475);
   U3047 : OAI22_X1 port map( A1 => n13616, A2 => n12246, B1 => n13552, B2 => 
                           n12240, ZN => n3482);
   U3048 : AOI221_X1 port map( B1 => n12162, B2 => n13997, C1 => n12156, C2 => 
                           n14168, A => n3490, ZN => n3483);
   U3049 : OAI22_X1 port map( A1 => n14095, A2 => n12150, B1 => n13759, B2 => 
                           n12144, ZN => n3490);
   U3050 : AOI221_X1 port map( B1 => n12258, B2 => n11754, C1 => n12252, C2 => 
                           n11574, A => n3463, ZN => n3456);
   U3051 : OAI22_X1 port map( A1 => n13615, A2 => n12246, B1 => n13551, B2 => 
                           n12240, ZN => n3463);
   U3052 : AOI221_X1 port map( B1 => n12162, B2 => n13996, C1 => n12156, C2 => 
                           n14167, A => n3471, ZN => n3464);
   U3053 : OAI22_X1 port map( A1 => n14094, A2 => n12150, B1 => n13758, B2 => 
                           n12144, ZN => n3471);
   U3054 : AOI221_X1 port map( B1 => n12258, B2 => n11755, C1 => n12252, C2 => 
                           n11575, A => n3444, ZN => n3437);
   U3055 : OAI22_X1 port map( A1 => n13614, A2 => n12246, B1 => n13550, B2 => 
                           n12240, ZN => n3444);
   U3056 : AOI221_X1 port map( B1 => n12162, B2 => n13995, C1 => n12156, C2 => 
                           n14166, A => n3452, ZN => n3445);
   U3057 : OAI22_X1 port map( A1 => n14093, A2 => n12150, B1 => n13757, B2 => 
                           n12144, ZN => n3452);
   U3058 : AOI221_X1 port map( B1 => n12258, B2 => n11756, C1 => n12252, C2 => 
                           n11576, A => n3425, ZN => n3418);
   U3059 : OAI22_X1 port map( A1 => n13613, A2 => n12246, B1 => n13549, B2 => 
                           n12240, ZN => n3425);
   U3060 : AOI221_X1 port map( B1 => n12162, B2 => n13994, C1 => n12156, C2 => 
                           n14165, A => n3433, ZN => n3426);
   U3061 : OAI22_X1 port map( A1 => n14092, A2 => n12150, B1 => n13756, B2 => 
                           n12144, ZN => n3433);
   U3062 : AOI221_X1 port map( B1 => n12258, B2 => n11757, C1 => n12252, C2 => 
                           n11577, A => n3406, ZN => n3399);
   U3063 : OAI22_X1 port map( A1 => n13612, A2 => n12246, B1 => n13548, B2 => 
                           n12240, ZN => n3406);
   U3064 : AOI221_X1 port map( B1 => n12162, B2 => n13993, C1 => n12156, C2 => 
                           n14164, A => n3414, ZN => n3407);
   U3065 : OAI22_X1 port map( A1 => n14091, A2 => n12150, B1 => n13755, B2 => 
                           n12144, ZN => n3414);
   U3066 : AOI221_X1 port map( B1 => n12258, B2 => n11758, C1 => n12252, C2 => 
                           n11578, A => n3387, ZN => n3380);
   U3067 : OAI22_X1 port map( A1 => n13611, A2 => n12246, B1 => n13547, B2 => 
                           n12240, ZN => n3387);
   U3068 : AOI221_X1 port map( B1 => n12162, B2 => n13992, C1 => n12156, C2 => 
                           n14163, A => n3395, ZN => n3388);
   U3069 : OAI22_X1 port map( A1 => n14090, A2 => n12150, B1 => n13754, B2 => 
                           n12144, ZN => n3395);
   U3070 : AOI221_X1 port map( B1 => n12258, B2 => n11759, C1 => n12252, C2 => 
                           n11579, A => n3368, ZN => n3361);
   U3071 : OAI22_X1 port map( A1 => n13610, A2 => n12246, B1 => n13546, B2 => 
                           n12240, ZN => n3368);
   U3072 : AOI221_X1 port map( B1 => n12162, B2 => n13991, C1 => n12156, C2 => 
                           n14162, A => n3376, ZN => n3369);
   U3073 : OAI22_X1 port map( A1 => n14089, A2 => n12150, B1 => n13753, B2 => 
                           n12144, ZN => n3376);
   U3074 : AOI221_X1 port map( B1 => n12258, B2 => n11760, C1 => n12252, C2 => 
                           n11580, A => n3349, ZN => n3342);
   U3075 : OAI22_X1 port map( A1 => n13609, A2 => n12246, B1 => n13545, B2 => 
                           n12240, ZN => n3349);
   U3076 : AOI221_X1 port map( B1 => n12162, B2 => n13990, C1 => n12156, C2 => 
                           n14161, A => n3357, ZN => n3350);
   U3077 : OAI22_X1 port map( A1 => n14088, A2 => n12150, B1 => n13752, B2 => 
                           n12144, ZN => n3357);
   U3078 : AOI221_X1 port map( B1 => n12258, B2 => n11761, C1 => n12252, C2 => 
                           n11581, A => n3330, ZN => n3323);
   U3079 : OAI22_X1 port map( A1 => n13608, A2 => n12246, B1 => n13544, B2 => 
                           n12240, ZN => n3330);
   U3080 : AOI221_X1 port map( B1 => n12162, B2 => n13989, C1 => n12156, C2 => 
                           n14160, A => n3338, ZN => n3331);
   U3081 : OAI22_X1 port map( A1 => n14087, A2 => n12150, B1 => n13751, B2 => 
                           n12144, ZN => n3338);
   U3082 : AOI221_X1 port map( B1 => n12163, B2 => n13827, C1 => n12157, C2 => 
                           n14159, A => n3319, ZN => n3312);
   U3083 : OAI22_X1 port map( A1 => n14086, A2 => n12151, B1 => n13750, B2 => 
                           n12145, ZN => n3319);
   U3084 : AOI221_X1 port map( B1 => n12259, B2 => n13864, C1 => n12253, C2 => 
                           n13868, A => n3311, ZN => n3304);
   U3085 : OAI22_X1 port map( A1 => n13607, A2 => n12247, B1 => n13543, B2 => 
                           n12241, ZN => n3311);
   U3086 : AOI221_X1 port map( B1 => n12163, B2 => n13826, C1 => n12157, C2 => 
                           n14158, A => n3300, ZN => n3293);
   U3087 : OAI22_X1 port map( A1 => n14085, A2 => n12151, B1 => n13749, B2 => 
                           n12145, ZN => n3300);
   U3088 : AOI221_X1 port map( B1 => n12259, B2 => n13863, C1 => n12253, C2 => 
                           n13867, A => n3292, ZN => n3285);
   U3089 : OAI22_X1 port map( A1 => n13606, A2 => n12247, B1 => n13542, B2 => 
                           n12241, ZN => n3292);
   U3090 : AOI221_X1 port map( B1 => n12163, B2 => n13825, C1 => n12157, C2 => 
                           n14157, A => n3281, ZN => n3274);
   U3091 : OAI22_X1 port map( A1 => n14084, A2 => n12151, B1 => n13748, B2 => 
                           n12145, ZN => n3281);
   U3092 : AOI221_X1 port map( B1 => n12259, B2 => n13862, C1 => n12253, C2 => 
                           n13866, A => n3273, ZN => n3266);
   U3093 : OAI22_X1 port map( A1 => n13605, A2 => n12247, B1 => n13541, B2 => 
                           n12241, ZN => n3273);
   U3094 : AOI221_X1 port map( B1 => n12163, B2 => n13824, C1 => n12157, C2 => 
                           n14156, A => n3260, ZN => n3239);
   U3095 : OAI22_X1 port map( A1 => n14083, A2 => n12151, B1 => n13747, B2 => 
                           n12145, ZN => n3260);
   U3096 : AOI221_X1 port map( B1 => n12259, B2 => n13861, C1 => n12253, C2 => 
                           n13865, A => n3236, ZN => n3215);
   U3097 : OAI22_X1 port map( A1 => n13604, A2 => n12247, B1 => n13540, B2 => 
                           n12241, ZN => n3236);
   U3098 : NAND2_X1 port map( A1 => n4450, A2 => n4466, ZN => n3246);
   U3099 : NAND2_X1 port map( A1 => n4450, A2 => n4465, ZN => n3247);
   U3100 : NAND2_X1 port map( A1 => n4454, A2 => n4466, ZN => n3251);
   U3101 : NAND2_X1 port map( A1 => n4454, A2 => n4465, ZN => n3252);
   U3102 : AOI221_X1 port map( B1 => n12302, B2 => n11762, C1 => n12296, C2 => 
                           n11582, A => n4430, ZN => n4427);
   U3103 : OAI22_X1 port map( A1 => n14408, A2 => n12290, B1 => n14385, B2 => 
                           n12284, ZN => n4430);
   U3104 : AOI221_X1 port map( B1 => n12302, B2 => n11763, C1 => n12296, C2 => 
                           n11583, A => n4354, ZN => n4351);
   U3105 : OAI22_X1 port map( A1 => n14404, A2 => n12290, B1 => n14381, B2 => 
                           n12284, ZN => n4354);
   U3106 : AOI221_X1 port map( B1 => n12302, B2 => n11764, C1 => n12296, C2 => 
                           n11584, A => n4335, ZN => n4332);
   U3107 : OAI22_X1 port map( A1 => n14403, A2 => n12290, B1 => n14380, B2 => 
                           n12284, ZN => n4335);
   U3108 : AOI221_X1 port map( B1 => n12306, B2 => n11765, C1 => n12300, C2 => 
                           n11585, A => n3328, ZN => n3325);
   U3109 : OAI22_X1 port map( A1 => n14253, A2 => n12294, B1 => n14217, B2 => 
                           n12288, ZN => n3328);
   U3110 : BUF_X1 port map( A => n1892, Z => n13210);
   U3111 : BUF_X1 port map( A => n1891, Z => n13213);
   U3112 : BUF_X1 port map( A => n1890, Z => n13216);
   U3113 : BUF_X1 port map( A => n1889, Z => n13219);
   U3114 : BUF_X1 port map( A => n1888, Z => n13222);
   U3115 : BUF_X1 port map( A => n1887, Z => n13225);
   U3116 : BUF_X1 port map( A => n1881, Z => n13243);
   U3117 : BUF_X1 port map( A => n1880, Z => n13246);
   U3118 : BUF_X1 port map( A => n1879, Z => n13249);
   U3119 : BUF_X1 port map( A => n1878, Z => n13252);
   U3120 : BUF_X1 port map( A => n1877, Z => n13255);
   U3121 : BUF_X1 port map( A => n1876, Z => n13258);
   U3122 : BUF_X1 port map( A => n1875, Z => n13261);
   U3123 : BUF_X1 port map( A => n1874, Z => n13264);
   U3124 : BUF_X1 port map( A => n1873, Z => n13267);
   U3125 : BUF_X1 port map( A => n1872, Z => n13270);
   U3126 : BUF_X1 port map( A => n1871, Z => n13273);
   U3127 : BUF_X1 port map( A => n1870, Z => n13276);
   U3128 : BUF_X1 port map( A => n1869, Z => n13279);
   U3129 : BUF_X1 port map( A => n1868, Z => n13282);
   U3130 : BUF_X1 port map( A => n1867, Z => n13285);
   U3131 : BUF_X1 port map( A => n1866, Z => n13288);
   U3132 : BUF_X1 port map( A => n1865, Z => n13291);
   U3133 : BUF_X1 port map( A => n1864, Z => n13294);
   U3134 : BUF_X1 port map( A => n1863, Z => n13297);
   U3135 : BUF_X1 port map( A => n1862, Z => n13300);
   U3136 : BUF_X1 port map( A => n1861, Z => n13303);
   U3137 : BUF_X1 port map( A => n1860, Z => n13306);
   U3138 : BUF_X1 port map( A => n1859, Z => n13309);
   U3139 : BUF_X1 port map( A => n1858, Z => n13312);
   U3140 : BUF_X1 port map( A => n1857, Z => n13315);
   U3141 : BUF_X1 port map( A => n1856, Z => n13318);
   U3142 : BUF_X1 port map( A => n1855, Z => n13321);
   U3143 : BUF_X1 port map( A => n1854, Z => n13324);
   U3144 : BUF_X1 port map( A => n1853, Z => n13327);
   U3145 : BUF_X1 port map( A => n1852, Z => n13330);
   U3146 : BUF_X1 port map( A => n1851, Z => n13333);
   U3147 : BUF_X1 port map( A => n1850, Z => n13336);
   U3148 : BUF_X1 port map( A => n1849, Z => n13339);
   U3149 : BUF_X1 port map( A => n1848, Z => n13342);
   U3150 : BUF_X1 port map( A => n1847, Z => n13345);
   U3151 : BUF_X1 port map( A => n1846, Z => n13348);
   U3152 : BUF_X1 port map( A => n1845, Z => n13351);
   U3153 : BUF_X1 port map( A => n1844, Z => n13354);
   U3154 : BUF_X1 port map( A => n1843, Z => n13357);
   U3155 : BUF_X1 port map( A => n1841, Z => n13380);
   U3156 : BUF_X1 port map( A => n1876, Z => n13257);
   U3157 : BUF_X1 port map( A => n1875, Z => n13260);
   U3158 : BUF_X1 port map( A => n1874, Z => n13263);
   U3159 : BUF_X1 port map( A => n1873, Z => n13266);
   U3160 : BUF_X1 port map( A => n1872, Z => n13269);
   U3161 : BUF_X1 port map( A => n1871, Z => n13272);
   U3162 : BUF_X1 port map( A => n1870, Z => n13275);
   U3163 : BUF_X1 port map( A => n1869, Z => n13278);
   U3164 : BUF_X1 port map( A => n1868, Z => n13281);
   U3165 : BUF_X1 port map( A => n1867, Z => n13284);
   U3166 : BUF_X1 port map( A => n1866, Z => n13287);
   U3167 : BUF_X1 port map( A => n1865, Z => n13290);
   U3168 : BUF_X1 port map( A => n1864, Z => n13293);
   U3169 : BUF_X1 port map( A => n1863, Z => n13296);
   U3170 : BUF_X1 port map( A => n1862, Z => n13299);
   U3171 : BUF_X1 port map( A => n1861, Z => n13302);
   U3172 : BUF_X1 port map( A => n1860, Z => n13305);
   U3173 : BUF_X1 port map( A => n1850, Z => n13335);
   U3174 : BUF_X1 port map( A => n1849, Z => n13338);
   U3175 : BUF_X1 port map( A => n1848, Z => n13341);
   U3176 : BUF_X1 port map( A => n1847, Z => n13344);
   U3177 : BUF_X1 port map( A => n1846, Z => n13347);
   U3178 : BUF_X1 port map( A => n1845, Z => n13350);
   U3179 : BUF_X1 port map( A => n1844, Z => n13353);
   U3180 : BUF_X1 port map( A => n1843, Z => n13356);
   U3181 : BUF_X1 port map( A => n1893, Z => n13206);
   U3182 : BUF_X1 port map( A => n1892, Z => n13209);
   U3183 : BUF_X1 port map( A => n1891, Z => n13212);
   U3184 : BUF_X1 port map( A => n1890, Z => n13215);
   U3185 : BUF_X1 port map( A => n1889, Z => n13218);
   U3186 : BUF_X1 port map( A => n1888, Z => n13221);
   U3187 : BUF_X1 port map( A => n1887, Z => n13224);
   U3188 : BUF_X1 port map( A => n1886, Z => n13227);
   U3189 : BUF_X1 port map( A => n1885, Z => n13230);
   U3190 : BUF_X1 port map( A => n1884, Z => n13233);
   U3191 : BUF_X1 port map( A => n1883, Z => n13236);
   U3192 : BUF_X1 port map( A => n1882, Z => n13239);
   U3193 : BUF_X1 port map( A => n1881, Z => n13242);
   U3194 : BUF_X1 port map( A => n1880, Z => n13245);
   U3195 : BUF_X1 port map( A => n1879, Z => n13248);
   U3196 : BUF_X1 port map( A => n1878, Z => n13251);
   U3197 : BUF_X1 port map( A => n1877, Z => n13254);
   U3198 : BUF_X1 port map( A => n1859, Z => n13308);
   U3199 : BUF_X1 port map( A => n1858, Z => n13311);
   U3200 : BUF_X1 port map( A => n1857, Z => n13314);
   U3201 : BUF_X1 port map( A => n1856, Z => n13317);
   U3202 : BUF_X1 port map( A => n1855, Z => n13320);
   U3203 : BUF_X1 port map( A => n1854, Z => n13323);
   U3204 : BUF_X1 port map( A => n1853, Z => n13326);
   U3205 : BUF_X1 port map( A => n1852, Z => n13329);
   U3206 : BUF_X1 port map( A => n1851, Z => n13332);
   U3207 : BUF_X1 port map( A => n1841, Z => n13379);
   U3208 : NAND2_X1 port map( A1 => n4469, A2 => n4450, ZN => n3257);
   U3209 : NAND2_X1 port map( A1 => n4470, A2 => n4450, ZN => n3256);
   U3210 : NAND2_X1 port map( A1 => n4449, A2 => n4450, ZN => n3223);
   U3211 : NAND2_X1 port map( A1 => n4451, A2 => n4450, ZN => n3222);
   U3212 : NAND2_X1 port map( A1 => n4469, A2 => n4454, ZN => n3262);
   U3213 : NAND2_X1 port map( A1 => n4470, A2 => n4454, ZN => n3261);
   U3214 : NAND2_X1 port map( A1 => n4449, A2 => n4454, ZN => n3228);
   U3215 : NAND2_X1 port map( A1 => n4451, A2 => n4454, ZN => n3227);
   U3216 : NAND2_X1 port map( A1 => n4458, A2 => n4452, ZN => n3232);
   U3217 : NAND2_X1 port map( A1 => n4457, A2 => n4452, ZN => n3233);
   U3218 : NAND2_X1 port map( A1 => n4458, A2 => n4455, ZN => n3237);
   U3219 : NAND2_X1 port map( A1 => n4457, A2 => n4455, ZN => n3238);
   U3220 : BUF_X1 port map( A => n1905, Z => n13171);
   U3221 : BUF_X1 port map( A => n1904, Z => n13174);
   U3222 : BUF_X1 port map( A => n1903, Z => n13177);
   U3223 : BUF_X1 port map( A => n1902, Z => n13180);
   U3224 : BUF_X1 port map( A => n1901, Z => n13183);
   U3225 : BUF_X1 port map( A => n1900, Z => n13186);
   U3226 : BUF_X1 port map( A => n1893, Z => n13207);
   U3227 : BUF_X1 port map( A => n1886, Z => n13228);
   U3228 : BUF_X1 port map( A => n1885, Z => n13231);
   U3229 : BUF_X1 port map( A => n1884, Z => n13234);
   U3230 : BUF_X1 port map( A => n1883, Z => n13237);
   U3231 : BUF_X1 port map( A => n1882, Z => n13240);
   U3232 : BUF_X1 port map( A => n1899, Z => n13189);
   U3233 : BUF_X1 port map( A => n1898, Z => n13192);
   U3234 : BUF_X1 port map( A => n1897, Z => n13195);
   U3235 : BUF_X1 port map( A => n1896, Z => n13198);
   U3236 : BUF_X1 port map( A => n1895, Z => n13201);
   U3237 : BUF_X1 port map( A => n1894, Z => n13204);
   U3238 : BUF_X1 port map( A => n1905, Z => n13172);
   U3239 : BUF_X1 port map( A => n1904, Z => n13175);
   U3240 : BUF_X1 port map( A => n1903, Z => n13178);
   U3241 : BUF_X1 port map( A => n1902, Z => n13181);
   U3242 : BUF_X1 port map( A => n1901, Z => n13184);
   U3243 : BUF_X1 port map( A => n1900, Z => n13187);
   U3244 : BUF_X1 port map( A => n1899, Z => n13190);
   U3245 : BUF_X1 port map( A => n1898, Z => n13193);
   U3246 : BUF_X1 port map( A => n1897, Z => n13196);
   U3247 : BUF_X1 port map( A => n1896, Z => n13199);
   U3248 : BUF_X1 port map( A => n1895, Z => n13202);
   U3249 : BUF_X1 port map( A => n1894, Z => n13205);
   U3250 : BUF_X1 port map( A => n1893, Z => n13208);
   U3251 : BUF_X1 port map( A => n1892, Z => n13211);
   U3252 : BUF_X1 port map( A => n1891, Z => n13214);
   U3253 : BUF_X1 port map( A => n1890, Z => n13217);
   U3254 : BUF_X1 port map( A => n1889, Z => n13220);
   U3255 : BUF_X1 port map( A => n1888, Z => n13223);
   U3256 : BUF_X1 port map( A => n1887, Z => n13226);
   U3257 : BUF_X1 port map( A => n1886, Z => n13229);
   U3258 : BUF_X1 port map( A => n1885, Z => n13232);
   U3259 : BUF_X1 port map( A => n1884, Z => n13235);
   U3260 : BUF_X1 port map( A => n1883, Z => n13238);
   U3261 : BUF_X1 port map( A => n1882, Z => n13241);
   U3262 : BUF_X1 port map( A => n1881, Z => n13244);
   U3263 : BUF_X1 port map( A => n1880, Z => n13247);
   U3264 : BUF_X1 port map( A => n1879, Z => n13250);
   U3265 : BUF_X1 port map( A => n1878, Z => n13253);
   U3266 : BUF_X1 port map( A => n1877, Z => n13256);
   U3267 : BUF_X1 port map( A => n1876, Z => n13259);
   U3268 : BUF_X1 port map( A => n1875, Z => n13262);
   U3269 : BUF_X1 port map( A => n1874, Z => n13265);
   U3270 : BUF_X1 port map( A => n1873, Z => n13268);
   U3271 : BUF_X1 port map( A => n1872, Z => n13271);
   U3272 : BUF_X1 port map( A => n1871, Z => n13274);
   U3273 : BUF_X1 port map( A => n1870, Z => n13277);
   U3274 : BUF_X1 port map( A => n1869, Z => n13280);
   U3275 : BUF_X1 port map( A => n1868, Z => n13283);
   U3276 : BUF_X1 port map( A => n1867, Z => n13286);
   U3277 : BUF_X1 port map( A => n1866, Z => n13289);
   U3278 : BUF_X1 port map( A => n1865, Z => n13292);
   U3279 : BUF_X1 port map( A => n1864, Z => n13295);
   U3280 : BUF_X1 port map( A => n1863, Z => n13298);
   U3281 : BUF_X1 port map( A => n1862, Z => n13301);
   U3282 : BUF_X1 port map( A => n1861, Z => n13304);
   U3283 : BUF_X1 port map( A => n1860, Z => n13307);
   U3284 : BUF_X1 port map( A => n1859, Z => n13310);
   U3285 : BUF_X1 port map( A => n1858, Z => n13313);
   U3286 : BUF_X1 port map( A => n1857, Z => n13316);
   U3287 : BUF_X1 port map( A => n1856, Z => n13319);
   U3288 : BUF_X1 port map( A => n1855, Z => n13322);
   U3289 : BUF_X1 port map( A => n1854, Z => n13325);
   U3290 : BUF_X1 port map( A => n1853, Z => n13328);
   U3291 : BUF_X1 port map( A => n1852, Z => n13331);
   U3292 : BUF_X1 port map( A => n1851, Z => n13334);
   U3293 : BUF_X1 port map( A => n1850, Z => n13337);
   U3294 : BUF_X1 port map( A => n1849, Z => n13340);
   U3295 : BUF_X1 port map( A => n1848, Z => n13343);
   U3296 : BUF_X1 port map( A => n1847, Z => n13346);
   U3297 : BUF_X1 port map( A => n1846, Z => n13349);
   U3298 : BUF_X1 port map( A => n1845, Z => n13352);
   U3299 : BUF_X1 port map( A => n1844, Z => n13355);
   U3300 : BUF_X1 port map( A => n1843, Z => n13358);
   U3301 : BUF_X1 port map( A => n1841, Z => n13381);
   U3302 : BUF_X1 port map( A => n1905, Z => n13170);
   U3303 : BUF_X1 port map( A => n1904, Z => n13173);
   U3304 : BUF_X1 port map( A => n1903, Z => n13176);
   U3305 : BUF_X1 port map( A => n1902, Z => n13179);
   U3306 : BUF_X1 port map( A => n1901, Z => n13182);
   U3307 : BUF_X1 port map( A => n1900, Z => n13185);
   U3308 : BUF_X1 port map( A => n1899, Z => n13188);
   U3309 : BUF_X1 port map( A => n1898, Z => n13191);
   U3310 : BUF_X1 port map( A => n1897, Z => n13194);
   U3311 : BUF_X1 port map( A => n1896, Z => n13197);
   U3312 : BUF_X1 port map( A => n1895, Z => n13200);
   U3313 : BUF_X1 port map( A => n1894, Z => n13203);
   U3314 : BUF_X1 port map( A => n3211, Z => n12332);
   U3315 : AND2_X1 port map( A1 => n4466, A2 => n4452, ZN => n3244);
   U3316 : AND2_X1 port map( A1 => n4452, A2 => n4465, ZN => n3243);
   U3317 : AND2_X1 port map( A1 => n4455, A2 => n4465, ZN => n3248);
   U3318 : AND2_X1 port map( A1 => n4455, A2 => n4466, ZN => n3249);
   U3319 : AND2_X1 port map( A1 => n4457, A2 => n4450, ZN => n3229);
   U3320 : AND2_X1 port map( A1 => n4458, A2 => n4450, ZN => n3230);
   U3321 : AND2_X1 port map( A1 => n4457, A2 => n4454, ZN => n3234);
   U3322 : AND2_X1 port map( A1 => n4458, A2 => n4454, ZN => n3235);
   U3323 : AND2_X1 port map( A1 => n4469, A2 => n4452, ZN => n3253);
   U3324 : AND2_X1 port map( A1 => n4469, A2 => n4455, ZN => n3258);
   U3325 : AND2_X1 port map( A1 => n4449, A2 => n4452, ZN => n3219);
   U3326 : AND2_X1 port map( A1 => n4451, A2 => n4452, ZN => n3220);
   U3327 : AND2_X1 port map( A1 => n4449, A2 => n4455, ZN => n3224);
   U3328 : AND2_X1 port map( A1 => n4451, A2 => n4455, ZN => n3225);
   U3329 : AND2_X1 port map( A1 => n4470, A2 => n4452, ZN => n3254);
   U3330 : BUF_X1 port map( A => n3211, Z => n12333);
   U3331 : BUF_X1 port map( A => n1950, Z => n12537);
   U3332 : BUF_X1 port map( A => n1950, Z => n12538);
   U3333 : AOI221_X1 port map( B1 => n12435, B2 => n4642, C1 => n12429, C2 => 
                           n4643, A => n3203, ZN => n3202);
   U3334 : OAI22_X1 port map( A1 => n8577, A2 => n12423, B1 => n8578, B2 => 
                           n12417, ZN => n3203);
   U3335 : AOI221_X1 port map( B1 => n12435, B2 => n4646, C1 => n12429, C2 => 
                           n4647, A => n3176, ZN => n3175);
   U3336 : OAI22_X1 port map( A1 => n8560, A2 => n12423, B1 => n8561, B2 => 
                           n12417, ZN => n3176);
   U3337 : AOI221_X1 port map( B1 => n12435, B2 => n4652, C1 => n12429, C2 => 
                           n4653, A => n3157, ZN => n3156);
   U3338 : OAI22_X1 port map( A1 => n8543, A2 => n12423, B1 => n8544, B2 => 
                           n12417, ZN => n3157);
   U3339 : AOI221_X1 port map( B1 => n12435, B2 => n4654, C1 => n12429, C2 => 
                           n4655, A => n3138, ZN => n3137);
   U3340 : OAI22_X1 port map( A1 => n8526, A2 => n12423, B1 => n8527, B2 => 
                           n12417, ZN => n3138);
   U3341 : AOI221_X1 port map( B1 => n12435, B2 => n8599, C1 => n12429, C2 => 
                           n8600, A => n3119, ZN => n3118);
   U3342 : OAI22_X1 port map( A1 => n8509, A2 => n12423, B1 => n8510, B2 => 
                           n12417, ZN => n3119);
   U3343 : AOI221_X1 port map( B1 => n12435, B2 => n8603, C1 => n12429, C2 => 
                           n8604, A => n3100, ZN => n3099);
   U3344 : OAI22_X1 port map( A1 => n8492, A2 => n12423, B1 => n8493, B2 => 
                           n12417, ZN => n3100);
   U3345 : AOI221_X1 port map( B1 => n12435, B2 => n8611, C1 => n12429, C2 => 
                           n8612, A => n3081, ZN => n3080);
   U3346 : OAI22_X1 port map( A1 => n8475, A2 => n12423, B1 => n8476, B2 => 
                           n12417, ZN => n3081);
   U3347 : AOI221_X1 port map( B1 => n12435, B2 => n8617, C1 => n12429, C2 => 
                           n8618, A => n3062, ZN => n3061);
   U3348 : OAI22_X1 port map( A1 => n8458, A2 => n12423, B1 => n8459, B2 => 
                           n12417, ZN => n3062);
   U3349 : AOI221_X1 port map( B1 => n12435, B2 => n8619, C1 => n12429, C2 => 
                           n8620, A => n3043, ZN => n3042);
   U3350 : OAI22_X1 port map( A1 => n8441, A2 => n12423, B1 => n8442, B2 => 
                           n12417, ZN => n3043);
   U3351 : AOI221_X1 port map( B1 => n12435, B2 => n8621, C1 => n12429, C2 => 
                           n8622, A => n3024, ZN => n3023);
   U3352 : OAI22_X1 port map( A1 => n8424, A2 => n12423, B1 => n8425, B2 => 
                           n12417, ZN => n3024);
   U3353 : AOI221_X1 port map( B1 => n12435, B2 => n8623, C1 => n12429, C2 => 
                           n8624, A => n3005, ZN => n3004);
   U3354 : OAI22_X1 port map( A1 => n8407, A2 => n12423, B1 => n8408, B2 => 
                           n12417, ZN => n3005);
   U3355 : AOI221_X1 port map( B1 => n12435, B2 => n8625, C1 => n12429, C2 => 
                           n8626, A => n2986, ZN => n2985);
   U3356 : OAI22_X1 port map( A1 => n8390, A2 => n12423, B1 => n8391, B2 => 
                           n12417, ZN => n2986);
   U3357 : AOI221_X1 port map( B1 => n12436, B2 => n8627, C1 => n12430, C2 => 
                           n8628, A => n2967, ZN => n2966);
   U3358 : OAI22_X1 port map( A1 => n8373, A2 => n12424, B1 => n8374, B2 => 
                           n12418, ZN => n2967);
   U3359 : AOI221_X1 port map( B1 => n12436, B2 => n8629, C1 => n12430, C2 => 
                           n8630, A => n2948, ZN => n2947);
   U3360 : OAI22_X1 port map( A1 => n8356, A2 => n12424, B1 => n8357, B2 => 
                           n12418, ZN => n2948);
   U3361 : AOI221_X1 port map( B1 => n12436, B2 => n8631, C1 => n12430, C2 => 
                           n8632, A => n2929, ZN => n2928);
   U3362 : OAI22_X1 port map( A1 => n8339, A2 => n12424, B1 => n8340, B2 => 
                           n12418, ZN => n2929);
   U3363 : AOI221_X1 port map( B1 => n12436, B2 => n8633, C1 => n12430, C2 => 
                           n8634, A => n2910, ZN => n2909);
   U3364 : OAI22_X1 port map( A1 => n8322, A2 => n12424, B1 => n8323, B2 => 
                           n12418, ZN => n2910);
   U3365 : AOI221_X1 port map( B1 => n12436, B2 => n8635, C1 => n12430, C2 => 
                           n8636, A => n2891, ZN => n2890);
   U3366 : OAI22_X1 port map( A1 => n8305, A2 => n12424, B1 => n8306, B2 => 
                           n12418, ZN => n2891);
   U3367 : AOI221_X1 port map( B1 => n12436, B2 => n8637, C1 => n12430, C2 => 
                           n8638, A => n2872, ZN => n2871);
   U3368 : OAI22_X1 port map( A1 => n8288, A2 => n12424, B1 => n8289, B2 => 
                           n12418, ZN => n2872);
   U3369 : AOI221_X1 port map( B1 => n12436, B2 => n8639, C1 => n12430, C2 => 
                           n8640, A => n2853, ZN => n2852);
   U3370 : OAI22_X1 port map( A1 => n8271, A2 => n12424, B1 => n8272, B2 => 
                           n12418, ZN => n2853);
   U3371 : AOI221_X1 port map( B1 => n12436, B2 => n8641, C1 => n12430, C2 => 
                           n8642, A => n2834, ZN => n2833);
   U3372 : OAI22_X1 port map( A1 => n8254, A2 => n12424, B1 => n8255, B2 => 
                           n12418, ZN => n2834);
   U3373 : AOI221_X1 port map( B1 => n12436, B2 => n8643, C1 => n12430, C2 => 
                           n8644, A => n2815, ZN => n2814);
   U3374 : OAI22_X1 port map( A1 => n8237, A2 => n12424, B1 => n8238, B2 => 
                           n12418, ZN => n2815);
   U3375 : AOI221_X1 port map( B1 => n12436, B2 => n8645, C1 => n12430, C2 => 
                           n8646, A => n2796, ZN => n2795);
   U3376 : OAI22_X1 port map( A1 => n8220, A2 => n12424, B1 => n8221, B2 => 
                           n12418, ZN => n2796);
   U3377 : AOI221_X1 port map( B1 => n12436, B2 => n8647, C1 => n12430, C2 => 
                           n8648, A => n2777, ZN => n2776);
   U3378 : OAI22_X1 port map( A1 => n8203, A2 => n12424, B1 => n8204, B2 => 
                           n12418, ZN => n2777);
   U3379 : AOI221_X1 port map( B1 => n12436, B2 => n8649, C1 => n12430, C2 => 
                           n8650, A => n2758, ZN => n2757);
   U3380 : OAI22_X1 port map( A1 => n8186, A2 => n12424, B1 => n8187, B2 => 
                           n12418, ZN => n2758);
   U3381 : AOI221_X1 port map( B1 => n12437, B2 => n8651, C1 => n12431, C2 => 
                           n8652, A => n2739, ZN => n2738);
   U3382 : OAI22_X1 port map( A1 => n8169, A2 => n12425, B1 => n8170, B2 => 
                           n12419, ZN => n2739);
   U3383 : AOI221_X1 port map( B1 => n12437, B2 => n8653, C1 => n12431, C2 => 
                           n8654, A => n2720, ZN => n2719);
   U3384 : OAI22_X1 port map( A1 => n8152, A2 => n12425, B1 => n8153, B2 => 
                           n12419, ZN => n2720);
   U3385 : AOI221_X1 port map( B1 => n12437, B2 => n8655, C1 => n12431, C2 => 
                           n8656, A => n2701, ZN => n2700);
   U3386 : OAI22_X1 port map( A1 => n8135, A2 => n12425, B1 => n8136, B2 => 
                           n12419, ZN => n2701);
   U3387 : AOI221_X1 port map( B1 => n12437, B2 => n8657, C1 => n12431, C2 => 
                           n8658, A => n2682, ZN => n2681);
   U3388 : OAI22_X1 port map( A1 => n8118, A2 => n12425, B1 => n8119, B2 => 
                           n12419, ZN => n2682);
   U3389 : AOI221_X1 port map( B1 => n12437, B2 => n8659, C1 => n12431, C2 => 
                           n8660, A => n2663, ZN => n2662);
   U3390 : OAI22_X1 port map( A1 => n8101, A2 => n12425, B1 => n8102, B2 => 
                           n12419, ZN => n2663);
   U3391 : AOI221_X1 port map( B1 => n12437, B2 => n8661, C1 => n12431, C2 => 
                           n8662, A => n2644, ZN => n2643);
   U3392 : OAI22_X1 port map( A1 => n8084, A2 => n12425, B1 => n8085, B2 => 
                           n12419, ZN => n2644);
   U3393 : AOI221_X1 port map( B1 => n12437, B2 => n8663, C1 => n12431, C2 => 
                           n8664, A => n2625, ZN => n2624);
   U3394 : OAI22_X1 port map( A1 => n8067, A2 => n12425, B1 => n8068, B2 => 
                           n12419, ZN => n2625);
   U3395 : AOI221_X1 port map( B1 => n12437, B2 => n8665, C1 => n12431, C2 => 
                           n8666, A => n2606, ZN => n2605);
   U3396 : OAI22_X1 port map( A1 => n8050, A2 => n12425, B1 => n8051, B2 => 
                           n12419, ZN => n2606);
   U3397 : AOI221_X1 port map( B1 => n12437, B2 => n8667, C1 => n12431, C2 => 
                           n8668, A => n2587, ZN => n2586);
   U3398 : OAI22_X1 port map( A1 => n8033, A2 => n12425, B1 => n8034, B2 => 
                           n12419, ZN => n2587);
   U3399 : AOI221_X1 port map( B1 => n12437, B2 => n8669, C1 => n12431, C2 => 
                           n8670, A => n2568, ZN => n2567);
   U3400 : OAI22_X1 port map( A1 => n8016, A2 => n12425, B1 => n8017, B2 => 
                           n12419, ZN => n2568);
   U3401 : AOI221_X1 port map( B1 => n12437, B2 => n8671, C1 => n12431, C2 => 
                           n8672, A => n2549, ZN => n2548);
   U3402 : OAI22_X1 port map( A1 => n7999, A2 => n12425, B1 => n8000, B2 => 
                           n12419, ZN => n2549);
   U3403 : AOI221_X1 port map( B1 => n12437, B2 => n8673, C1 => n12431, C2 => 
                           n8674, A => n2530, ZN => n2529);
   U3404 : OAI22_X1 port map( A1 => n7982, A2 => n12425, B1 => n7983, B2 => 
                           n12419, ZN => n2530);
   U3405 : AOI221_X1 port map( B1 => n12438, B2 => n8675, C1 => n12432, C2 => 
                           n8676, A => n2511, ZN => n2510);
   U3406 : OAI22_X1 port map( A1 => n7965, A2 => n12426, B1 => n7966, B2 => 
                           n12420, ZN => n2511);
   U3407 : AOI221_X1 port map( B1 => n12438, B2 => n8677, C1 => n12432, C2 => 
                           n8678, A => n2492, ZN => n2491);
   U3408 : OAI22_X1 port map( A1 => n7948, A2 => n12426, B1 => n7949, B2 => 
                           n12420, ZN => n2492);
   U3409 : AOI221_X1 port map( B1 => n12438, B2 => n8679, C1 => n12432, C2 => 
                           n8680, A => n2473, ZN => n2472);
   U3410 : OAI22_X1 port map( A1 => n7931, A2 => n12426, B1 => n7932, B2 => 
                           n12420, ZN => n2473);
   U3411 : AOI221_X1 port map( B1 => n12438, B2 => n8681, C1 => n12432, C2 => 
                           n8682, A => n2454, ZN => n2453);
   U3412 : OAI22_X1 port map( A1 => n7914, A2 => n12426, B1 => n7915, B2 => 
                           n12420, ZN => n2454);
   U3413 : AOI221_X1 port map( B1 => n12438, B2 => n8683, C1 => n12432, C2 => 
                           n8684, A => n2435, ZN => n2434);
   U3414 : OAI22_X1 port map( A1 => n7897, A2 => n12426, B1 => n7898, B2 => 
                           n12420, ZN => n2435);
   U3415 : AOI221_X1 port map( B1 => n12438, B2 => n8685, C1 => n12432, C2 => 
                           n8686, A => n2416, ZN => n2415);
   U3416 : OAI22_X1 port map( A1 => n7880, A2 => n12426, B1 => n7881, B2 => 
                           n12420, ZN => n2416);
   U3417 : AOI221_X1 port map( B1 => n12438, B2 => n8687, C1 => n12432, C2 => 
                           n8688, A => n2397, ZN => n2396);
   U3418 : OAI22_X1 port map( A1 => n7863, A2 => n12426, B1 => n7864, B2 => 
                           n12420, ZN => n2397);
   U3419 : AOI221_X1 port map( B1 => n12438, B2 => n8689, C1 => n12432, C2 => 
                           n8690, A => n2378, ZN => n2377);
   U3420 : OAI22_X1 port map( A1 => n7846, A2 => n12426, B1 => n7847, B2 => 
                           n12420, ZN => n2378);
   U3421 : AOI221_X1 port map( B1 => n12438, B2 => n8691, C1 => n12432, C2 => 
                           n8692, A => n2359, ZN => n2358);
   U3422 : OAI22_X1 port map( A1 => n7829, A2 => n12426, B1 => n7830, B2 => 
                           n12420, ZN => n2359);
   U3423 : AOI221_X1 port map( B1 => n12438, B2 => n8693, C1 => n12432, C2 => 
                           n8694, A => n2340, ZN => n2339);
   U3424 : OAI22_X1 port map( A1 => n7812, A2 => n12426, B1 => n7813, B2 => 
                           n12420, ZN => n2340);
   U3425 : AOI221_X1 port map( B1 => n12438, B2 => n8695, C1 => n12432, C2 => 
                           n8696, A => n2321, ZN => n2320);
   U3426 : OAI22_X1 port map( A1 => n7795, A2 => n12426, B1 => n7796, B2 => 
                           n12420, ZN => n2321);
   U3427 : AOI221_X1 port map( B1 => n12438, B2 => n4656, C1 => n12432, C2 => 
                           n4657, A => n2302, ZN => n2301);
   U3428 : OAI22_X1 port map( A1 => n7778, A2 => n12426, B1 => n7779, B2 => 
                           n12420, ZN => n2302);
   U3429 : AOI221_X1 port map( B1 => n12439, B2 => n4658, C1 => n12433, C2 => 
                           n4659, A => n2283, ZN => n2282);
   U3430 : OAI22_X1 port map( A1 => n7761, A2 => n12427, B1 => n7762, B2 => 
                           n12421, ZN => n2283);
   U3431 : AOI221_X1 port map( B1 => n12439, B2 => n4660, C1 => n12433, C2 => 
                           n4661, A => n2264, ZN => n2263);
   U3432 : OAI22_X1 port map( A1 => n7744, A2 => n12427, B1 => n7745, B2 => 
                           n12421, ZN => n2264);
   U3433 : AOI221_X1 port map( B1 => n12439, B2 => n4662, C1 => n12433, C2 => 
                           n4663, A => n2245, ZN => n2244);
   U3434 : OAI22_X1 port map( A1 => n7642, A2 => n12427, B1 => n7643, B2 => 
                           n12421, ZN => n2245);
   U3435 : AOI221_X1 port map( B1 => n12439, B2 => n4664, C1 => n12433, C2 => 
                           n4665, A => n2226, ZN => n2225);
   U3436 : OAI22_X1 port map( A1 => n7625, A2 => n12427, B1 => n7626, B2 => 
                           n12421, ZN => n2226);
   U3437 : AOI221_X1 port map( B1 => n12439, B2 => n4666, C1 => n12433, C2 => 
                           n4667, A => n2207, ZN => n2206);
   U3438 : OAI22_X1 port map( A1 => n7521, A2 => n12427, B1 => n7522, B2 => 
                           n12421, ZN => n2207);
   U3439 : AOI221_X1 port map( B1 => n12439, B2 => n4668, C1 => n12433, C2 => 
                           n4669, A => n2188, ZN => n2187);
   U3440 : OAI22_X1 port map( A1 => n7504, A2 => n12427, B1 => n7505, B2 => 
                           n12421, ZN => n2188);
   U3441 : AOI221_X1 port map( B1 => n12439, B2 => n4670, C1 => n12433, C2 => 
                           n4671, A => n2169, ZN => n2168);
   U3442 : OAI22_X1 port map( A1 => n7402, A2 => n12427, B1 => n7403, B2 => 
                           n12421, ZN => n2169);
   U3443 : AOI221_X1 port map( B1 => n12439, B2 => n4672, C1 => n12433, C2 => 
                           n4673, A => n2150, ZN => n2149);
   U3444 : OAI22_X1 port map( A1 => n7385, A2 => n12427, B1 => n7386, B2 => 
                           n12421, ZN => n2150);
   U3445 : AOI221_X1 port map( B1 => n12439, B2 => n4674, C1 => n12433, C2 => 
                           n4675, A => n2131, ZN => n2130);
   U3446 : OAI22_X1 port map( A1 => n7368, A2 => n12427, B1 => n7369, B2 => 
                           n12421, ZN => n2131);
   U3447 : AOI221_X1 port map( B1 => n12439, B2 => n4676, C1 => n12433, C2 => 
                           n4677, A => n2112, ZN => n2111);
   U3448 : OAI22_X1 port map( A1 => n7269, A2 => n12427, B1 => n7270, B2 => 
                           n12421, ZN => n2112);
   U3449 : AOI221_X1 port map( B1 => n12439, B2 => n4678, C1 => n12433, C2 => 
                           n4679, A => n2093, ZN => n2092);
   U3450 : OAI22_X1 port map( A1 => n7252, A2 => n12427, B1 => n7253, B2 => 
                           n12421, ZN => n2093);
   U3451 : AOI221_X1 port map( B1 => n12439, B2 => n4682, C1 => n12433, C2 => 
                           n4683, A => n2074, ZN => n2073);
   U3452 : OAI22_X1 port map( A1 => n7235, A2 => n12427, B1 => n7236, B2 => 
                           n12421, ZN => n2074);
   U3453 : AOI221_X1 port map( B1 => n12440, B2 => n4472, C1 => n12434, C2 => 
                           n4473, A => n2055, ZN => n2054);
   U3454 : OAI22_X1 port map( A1 => n7138, A2 => n12428, B1 => n7139, B2 => 
                           n12422, ZN => n2055);
   U3455 : AOI221_X1 port map( B1 => n12536, B2 => n9952, C1 => n12530, C2 => 
                           n9888, A => n2047, ZN => n2046);
   U3456 : OAI22_X1 port map( A1 => n14435, A2 => n12524, B1 => n14412, B2 => 
                           n12518, ZN => n2047);
   U3457 : AOI221_X1 port map( B1 => n12440, B2 => n4474, C1 => n12434, C2 => 
                           n4475, A => n2036, ZN => n2035);
   U3458 : OAI22_X1 port map( A1 => n7121, A2 => n12428, B1 => n7122, B2 => 
                           n12422, ZN => n2036);
   U3459 : AOI221_X1 port map( B1 => n12536, B2 => n9951, C1 => n12530, C2 => 
                           n9887, A => n2028, ZN => n2027);
   U3460 : OAI22_X1 port map( A1 => n14434, A2 => n12524, B1 => n14411, B2 => 
                           n12518, ZN => n2028);
   U3461 : AOI221_X1 port map( B1 => n12440, B2 => n4476, C1 => n12434, C2 => 
                           n4477, A => n2017, ZN => n2016);
   U3462 : OAI22_X1 port map( A1 => n4860, A2 => n12428, B1 => n4861, B2 => 
                           n12422, ZN => n2017);
   U3463 : AOI221_X1 port map( B1 => n12536, B2 => n9950, C1 => n12530, C2 => 
                           n9886, A => n2009, ZN => n2008);
   U3464 : OAI22_X1 port map( A1 => n14433, A2 => n12524, B1 => n14410, B2 => 
                           n12518, ZN => n2009);
   U3465 : AOI221_X1 port map( B1 => n12440, B2 => n4478, C1 => n12434, C2 => 
                           n4479, A => n1984, ZN => n1981);
   U3466 : OAI22_X1 port map( A1 => n4843, A2 => n12428, B1 => n4844, B2 => 
                           n12422, ZN => n1984);
   U3467 : AOI221_X1 port map( B1 => n12536, B2 => n9949, C1 => n12530, C2 => 
                           n9885, A => n1960, ZN => n1957);
   U3468 : OAI22_X1 port map( A1 => n13392, A2 => n12524, B1 => n14409, B2 => 
                           n12518, ZN => n1960);
   U3469 : AOI221_X1 port map( B1 => n12411, B2 => n4480, C1 => n12405, C2 => 
                           n4481, A => n3206, ZN => n3201);
   U3470 : OAI22_X1 port map( A1 => n8579, A2 => n12399, B1 => n8580, B2 => 
                           n12393, ZN => n3206);
   U3471 : AOI221_X1 port map( B1 => n12411, B2 => n4648, C1 => n12405, C2 => 
                           n4649, A => n3177, ZN => n3174);
   U3472 : OAI22_X1 port map( A1 => n8562, A2 => n12399, B1 => n8563, B2 => 
                           n12393, ZN => n3177);
   U3473 : AOI221_X1 port map( B1 => n12411, B2 => n4482, C1 => n12405, C2 => 
                           n4483, A => n3158, ZN => n3155);
   U3474 : OAI22_X1 port map( A1 => n8545, A2 => n12399, B1 => n8546, B2 => 
                           n12393, ZN => n3158);
   U3475 : AOI221_X1 port map( B1 => n12411, B2 => n4484, C1 => n12405, C2 => 
                           n4485, A => n3139, ZN => n3136);
   U3476 : OAI22_X1 port map( A1 => n8528, A2 => n12399, B1 => n8529, B2 => 
                           n12393, ZN => n3139);
   U3477 : AOI221_X1 port map( B1 => n12411, B2 => n7080, C1 => n12405, C2 => 
                           n7081, A => n3120, ZN => n3117);
   U3478 : OAI22_X1 port map( A1 => n8511, A2 => n12399, B1 => n8512, B2 => 
                           n12393, ZN => n3120);
   U3479 : AOI221_X1 port map( B1 => n12411, B2 => n8605, C1 => n12405, C2 => 
                           n8606, A => n3101, ZN => n3098);
   U3480 : OAI22_X1 port map( A1 => n8494, A2 => n12399, B1 => n8495, B2 => 
                           n12393, ZN => n3101);
   U3481 : AOI221_X1 port map( B1 => n12411, B2 => n8613, C1 => n12405, C2 => 
                           n8614, A => n3082, ZN => n3079);
   U3482 : OAI22_X1 port map( A1 => n8477, A2 => n12399, B1 => n8478, B2 => 
                           n12393, ZN => n3082);
   U3483 : AOI221_X1 port map( B1 => n12411, B2 => n7084, C1 => n12405, C2 => 
                           n7085, A => n3063, ZN => n3060);
   U3484 : OAI22_X1 port map( A1 => n8460, A2 => n12399, B1 => n8461, B2 => 
                           n12393, ZN => n3063);
   U3485 : AOI221_X1 port map( B1 => n12411, B2 => n7088, C1 => n12405, C2 => 
                           n7089, A => n3044, ZN => n3041);
   U3486 : OAI22_X1 port map( A1 => n8443, A2 => n12399, B1 => n8444, B2 => 
                           n12393, ZN => n3044);
   U3487 : AOI221_X1 port map( B1 => n12411, B2 => n7092, C1 => n12405, C2 => 
                           n7093, A => n3025, ZN => n3022);
   U3488 : OAI22_X1 port map( A1 => n8426, A2 => n12399, B1 => n8427, B2 => 
                           n12393, ZN => n3025);
   U3489 : AOI221_X1 port map( B1 => n12411, B2 => n7096, C1 => n12405, C2 => 
                           n7097, A => n3006, ZN => n3003);
   U3490 : OAI22_X1 port map( A1 => n8409, A2 => n12399, B1 => n8410, B2 => 
                           n12393, ZN => n3006);
   U3491 : AOI221_X1 port map( B1 => n12411, B2 => n7100, C1 => n12405, C2 => 
                           n7101, A => n2987, ZN => n2984);
   U3492 : OAI22_X1 port map( A1 => n8392, A2 => n12399, B1 => n8393, B2 => 
                           n12393, ZN => n2987);
   U3493 : AOI221_X1 port map( B1 => n12412, B2 => n7104, C1 => n12406, C2 => 
                           n7105, A => n2968, ZN => n2965);
   U3494 : OAI22_X1 port map( A1 => n8375, A2 => n12400, B1 => n8376, B2 => 
                           n12394, ZN => n2968);
   U3495 : AOI221_X1 port map( B1 => n12412, B2 => n7130, C1 => n12406, C2 => 
                           n7131, A => n2949, ZN => n2946);
   U3496 : OAI22_X1 port map( A1 => n8358, A2 => n12400, B1 => n8359, B2 => 
                           n12394, ZN => n2949);
   U3497 : AOI221_X1 port map( B1 => n12412, B2 => n7154, C1 => n12406, C2 => 
                           n7155, A => n2930, ZN => n2927);
   U3498 : OAI22_X1 port map( A1 => n8341, A2 => n12400, B1 => n8342, B2 => 
                           n12394, ZN => n2930);
   U3499 : AOI221_X1 port map( B1 => n12412, B2 => n7158, C1 => n12406, C2 => 
                           n7159, A => n2911, ZN => n2908);
   U3500 : OAI22_X1 port map( A1 => n8324, A2 => n12400, B1 => n8325, B2 => 
                           n12394, ZN => n2911);
   U3501 : AOI221_X1 port map( B1 => n12412, B2 => n7162, C1 => n12406, C2 => 
                           n7163, A => n2892, ZN => n2889);
   U3502 : OAI22_X1 port map( A1 => n8307, A2 => n12400, B1 => n8308, B2 => 
                           n12394, ZN => n2892);
   U3503 : AOI221_X1 port map( B1 => n12412, B2 => n7166, C1 => n12406, C2 => 
                           n7167, A => n2873, ZN => n2870);
   U3504 : OAI22_X1 port map( A1 => n8290, A2 => n12400, B1 => n8291, B2 => 
                           n12394, ZN => n2873);
   U3505 : AOI221_X1 port map( B1 => n12412, B2 => n7170, C1 => n12406, C2 => 
                           n7171, A => n2854, ZN => n2851);
   U3506 : OAI22_X1 port map( A1 => n8273, A2 => n12400, B1 => n8274, B2 => 
                           n12394, ZN => n2854);
   U3507 : AOI221_X1 port map( B1 => n12412, B2 => n7174, C1 => n12406, C2 => 
                           n7175, A => n2835, ZN => n2832);
   U3508 : OAI22_X1 port map( A1 => n8256, A2 => n12400, B1 => n8257, B2 => 
                           n12394, ZN => n2835);
   U3509 : AOI221_X1 port map( B1 => n12412, B2 => n7178, C1 => n12406, C2 => 
                           n7179, A => n2816, ZN => n2813);
   U3510 : OAI22_X1 port map( A1 => n8239, A2 => n12400, B1 => n8240, B2 => 
                           n12394, ZN => n2816);
   U3511 : AOI221_X1 port map( B1 => n12412, B2 => n7182, C1 => n12406, C2 => 
                           n7183, A => n2797, ZN => n2794);
   U3512 : OAI22_X1 port map( A1 => n8222, A2 => n12400, B1 => n8223, B2 => 
                           n12394, ZN => n2797);
   U3513 : AOI221_X1 port map( B1 => n12412, B2 => n7186, C1 => n12406, C2 => 
                           n7187, A => n2778, ZN => n2775);
   U3514 : OAI22_X1 port map( A1 => n8205, A2 => n12400, B1 => n8206, B2 => 
                           n12394, ZN => n2778);
   U3515 : AOI221_X1 port map( B1 => n12412, B2 => n7190, C1 => n12406, C2 => 
                           n7191, A => n2759, ZN => n2756);
   U3516 : OAI22_X1 port map( A1 => n8188, A2 => n12400, B1 => n8189, B2 => 
                           n12394, ZN => n2759);
   U3517 : AOI221_X1 port map( B1 => n12413, B2 => n7194, C1 => n12407, C2 => 
                           n7195, A => n2740, ZN => n2737);
   U3518 : OAI22_X1 port map( A1 => n8171, A2 => n12401, B1 => n8172, B2 => 
                           n12395, ZN => n2740);
   U3519 : AOI221_X1 port map( B1 => n12413, B2 => n7198, C1 => n12407, C2 => 
                           n7199, A => n2721, ZN => n2718);
   U3520 : OAI22_X1 port map( A1 => n8154, A2 => n12401, B1 => n8155, B2 => 
                           n12395, ZN => n2721);
   U3521 : AOI221_X1 port map( B1 => n12413, B2 => n7202, C1 => n12407, C2 => 
                           n8708, A => n2702, ZN => n2699);
   U3522 : OAI22_X1 port map( A1 => n8137, A2 => n12401, B1 => n8138, B2 => 
                           n12395, ZN => n2702);
   U3523 : AOI221_X1 port map( B1 => n12413, B2 => n7205, C1 => n12407, C2 => 
                           n8707, A => n2683, ZN => n2680);
   U3524 : OAI22_X1 port map( A1 => n8120, A2 => n12401, B1 => n8121, B2 => 
                           n12395, ZN => n2683);
   U3525 : AOI221_X1 port map( B1 => n12413, B2 => n7208, C1 => n12407, C2 => 
                           n8706, A => n2664, ZN => n2661);
   U3526 : OAI22_X1 port map( A1 => n8103, A2 => n12401, B1 => n8104, B2 => 
                           n12395, ZN => n2664);
   U3527 : AOI221_X1 port map( B1 => n12413, B2 => n7211, C1 => n12407, C2 => 
                           n8705, A => n2645, ZN => n2642);
   U3528 : OAI22_X1 port map( A1 => n8086, A2 => n12401, B1 => n8087, B2 => 
                           n12395, ZN => n2645);
   U3529 : AOI221_X1 port map( B1 => n12413, B2 => n7214, C1 => n12407, C2 => 
                           n8704, A => n2626, ZN => n2623);
   U3530 : OAI22_X1 port map( A1 => n8069, A2 => n12401, B1 => n8070, B2 => 
                           n12395, ZN => n2626);
   U3531 : AOI221_X1 port map( B1 => n12413, B2 => n7217, C1 => n12407, C2 => 
                           n8703, A => n2607, ZN => n2604);
   U3532 : OAI22_X1 port map( A1 => n8052, A2 => n12401, B1 => n8053, B2 => 
                           n12395, ZN => n2607);
   U3533 : AOI221_X1 port map( B1 => n12413, B2 => n7220, C1 => n12407, C2 => 
                           n8702, A => n2588, ZN => n2585);
   U3534 : OAI22_X1 port map( A1 => n8035, A2 => n12401, B1 => n8036, B2 => 
                           n12395, ZN => n2588);
   U3535 : AOI221_X1 port map( B1 => n12413, B2 => n7223, C1 => n12407, C2 => 
                           n8701, A => n2569, ZN => n2566);
   U3536 : OAI22_X1 port map( A1 => n8018, A2 => n12401, B1 => n8019, B2 => 
                           n12395, ZN => n2569);
   U3537 : AOI221_X1 port map( B1 => n12413, B2 => n7226, C1 => n12407, C2 => 
                           n8700, A => n2550, ZN => n2547);
   U3538 : OAI22_X1 port map( A1 => n8001, A2 => n12401, B1 => n8002, B2 => 
                           n12395, ZN => n2550);
   U3539 : AOI221_X1 port map( B1 => n12413, B2 => n7229, C1 => n12407, C2 => 
                           n8699, A => n2531, ZN => n2528);
   U3540 : OAI22_X1 port map( A1 => n7984, A2 => n12401, B1 => n7985, B2 => 
                           n12395, ZN => n2531);
   U3541 : AOI221_X1 port map( B1 => n12414, B2 => n7232, C1 => n12408, C2 => 
                           n8698, A => n2512, ZN => n2509);
   U3542 : OAI22_X1 port map( A1 => n7967, A2 => n12402, B1 => n7968, B2 => 
                           n12396, ZN => n2512);
   U3543 : AOI221_X1 port map( B1 => n12414, B2 => n7245, C1 => n12408, C2 => 
                           n8697, A => n2493, ZN => n2490);
   U3544 : OAI22_X1 port map( A1 => n7950, A2 => n12402, B1 => n7951, B2 => 
                           n12396, ZN => n2493);
   U3545 : AOI221_X1 port map( B1 => n12414, B2 => n7278, C1 => n12408, C2 => 
                           n7279, A => n2474, ZN => n2471);
   U3546 : OAI22_X1 port map( A1 => n7933, A2 => n12402, B1 => n7934, B2 => 
                           n12396, ZN => n2474);
   U3547 : AOI221_X1 port map( B1 => n12414, B2 => n7282, C1 => n12408, C2 => 
                           n7283, A => n2455, ZN => n2452);
   U3548 : OAI22_X1 port map( A1 => n7916, A2 => n12402, B1 => n7917, B2 => 
                           n12396, ZN => n2455);
   U3549 : AOI221_X1 port map( B1 => n12414, B2 => n7286, C1 => n12408, C2 => 
                           n7287, A => n2436, ZN => n2433);
   U3550 : OAI22_X1 port map( A1 => n7899, A2 => n12402, B1 => n7900, B2 => 
                           n12396, ZN => n2436);
   U3551 : AOI221_X1 port map( B1 => n12414, B2 => n7290, C1 => n12408, C2 => 
                           n7291, A => n2417, ZN => n2414);
   U3552 : OAI22_X1 port map( A1 => n7882, A2 => n12402, B1 => n7883, B2 => 
                           n12396, ZN => n2417);
   U3553 : AOI221_X1 port map( B1 => n12414, B2 => n7294, C1 => n12408, C2 => 
                           n7295, A => n2398, ZN => n2395);
   U3554 : OAI22_X1 port map( A1 => n7865, A2 => n12402, B1 => n7866, B2 => 
                           n12396, ZN => n2398);
   U3555 : AOI221_X1 port map( B1 => n12414, B2 => n7298, C1 => n12408, C2 => 
                           n7299, A => n2379, ZN => n2376);
   U3556 : OAI22_X1 port map( A1 => n7848, A2 => n12402, B1 => n7849, B2 => 
                           n12396, ZN => n2379);
   U3557 : AOI221_X1 port map( B1 => n12414, B2 => n7302, C1 => n12408, C2 => 
                           n7303, A => n2360, ZN => n2357);
   U3558 : OAI22_X1 port map( A1 => n7831, A2 => n12402, B1 => n7832, B2 => 
                           n12396, ZN => n2360);
   U3559 : AOI221_X1 port map( B1 => n12414, B2 => n7306, C1 => n12408, C2 => 
                           n7307, A => n2341, ZN => n2338);
   U3560 : OAI22_X1 port map( A1 => n7814, A2 => n12402, B1 => n7815, B2 => 
                           n12396, ZN => n2341);
   U3561 : AOI221_X1 port map( B1 => n12414, B2 => n7310, C1 => n12408, C2 => 
                           n7311, A => n2322, ZN => n2319);
   U3562 : OAI22_X1 port map( A1 => n7797, A2 => n12402, B1 => n7798, B2 => 
                           n12396, ZN => n2322);
   U3563 : AOI221_X1 port map( B1 => n12414, B2 => n7314, C1 => n12408, C2 => 
                           n7315, A => n2303, ZN => n2300);
   U3564 : OAI22_X1 port map( A1 => n7780, A2 => n12402, B1 => n7781, B2 => 
                           n12396, ZN => n2303);
   U3565 : AOI221_X1 port map( B1 => n12415, B2 => n7318, C1 => n12409, C2 => 
                           n7319, A => n2284, ZN => n2281);
   U3566 : OAI22_X1 port map( A1 => n7763, A2 => n12403, B1 => n7764, B2 => 
                           n12397, ZN => n2284);
   U3567 : AOI221_X1 port map( B1 => n12415, B2 => n7322, C1 => n12409, C2 => 
                           n7323, A => n2265, ZN => n2262);
   U3568 : OAI22_X1 port map( A1 => n7746, A2 => n12403, B1 => n7747, B2 => 
                           n12397, ZN => n2265);
   U3569 : AOI221_X1 port map( B1 => n12415, B2 => n4486, C1 => n12409, C2 => 
                           n4487, A => n2246, ZN => n2243);
   U3570 : OAI22_X1 port map( A1 => n7644, A2 => n12403, B1 => n7645, B2 => 
                           n12397, ZN => n2246);
   U3571 : AOI221_X1 port map( B1 => n12415, B2 => n4488, C1 => n12409, C2 => 
                           n4489, A => n2227, ZN => n2224);
   U3572 : OAI22_X1 port map( A1 => n7627, A2 => n12403, B1 => n7628, B2 => 
                           n12397, ZN => n2227);
   U3573 : AOI221_X1 port map( B1 => n12415, B2 => n4490, C1 => n12409, C2 => 
                           n4491, A => n2208, ZN => n2205);
   U3574 : OAI22_X1 port map( A1 => n7523, A2 => n12403, B1 => n7524, B2 => 
                           n12397, ZN => n2208);
   U3575 : AOI221_X1 port map( B1 => n12415, B2 => n4492, C1 => n12409, C2 => 
                           n4493, A => n2189, ZN => n2186);
   U3576 : OAI22_X1 port map( A1 => n7506, A2 => n12403, B1 => n7507, B2 => 
                           n12397, ZN => n2189);
   U3577 : AOI221_X1 port map( B1 => n12415, B2 => n4494, C1 => n12409, C2 => 
                           n4495, A => n2170, ZN => n2167);
   U3578 : OAI22_X1 port map( A1 => n7404, A2 => n12403, B1 => n7490, B2 => 
                           n12397, ZN => n2170);
   U3579 : AOI221_X1 port map( B1 => n12415, B2 => n4496, C1 => n12409, C2 => 
                           n4497, A => n2151, ZN => n2148);
   U3580 : OAI22_X1 port map( A1 => n7387, A2 => n12403, B1 => n7388, B2 => 
                           n12397, ZN => n2151);
   U3581 : AOI221_X1 port map( B1 => n12415, B2 => n4498, C1 => n12409, C2 => 
                           n4499, A => n2132, ZN => n2129);
   U3582 : OAI22_X1 port map( A1 => n7370, A2 => n12403, B1 => n7371, B2 => 
                           n12397, ZN => n2132);
   U3583 : AOI221_X1 port map( B1 => n12415, B2 => n4500, C1 => n12409, C2 => 
                           n4501, A => n2113, ZN => n2110);
   U3584 : OAI22_X1 port map( A1 => n7271, A2 => n12403, B1 => n7272, B2 => 
                           n12397, ZN => n2113);
   U3585 : AOI221_X1 port map( B1 => n12415, B2 => n4502, C1 => n12409, C2 => 
                           n4503, A => n2094, ZN => n2091);
   U3586 : OAI22_X1 port map( A1 => n7254, A2 => n12403, B1 => n7255, B2 => 
                           n12397, ZN => n2094);
   U3587 : AOI221_X1 port map( B1 => n12415, B2 => n4684, C1 => n12409, C2 => 
                           n4685, A => n2075, ZN => n2072);
   U3588 : OAI22_X1 port map( A1 => n7237, A2 => n12403, B1 => n7238, B2 => 
                           n12397, ZN => n2075);
   U3589 : AOI221_X1 port map( B1 => n12416, B2 => n4504, C1 => n12410, C2 => 
                           n4505, A => n2056, ZN => n2053);
   U3590 : OAI22_X1 port map( A1 => n7140, A2 => n12404, B1 => n7141, B2 => 
                           n12398, ZN => n2056);
   U3591 : AOI221_X1 port map( B1 => n12416, B2 => n4506, C1 => n12410, C2 => 
                           n4507, A => n2037, ZN => n2034);
   U3592 : OAI22_X1 port map( A1 => n7123, A2 => n12404, B1 => n7124, B2 => 
                           n12398, ZN => n2037);
   U3593 : AOI221_X1 port map( B1 => n12416, B2 => n4508, C1 => n12410, C2 => 
                           n4509, A => n2018, ZN => n2015);
   U3594 : OAI22_X1 port map( A1 => n7106, A2 => n12404, B1 => n7107, B2 => 
                           n12398, ZN => n2018);
   U3595 : AOI221_X1 port map( B1 => n12416, B2 => n4510, C1 => n12410, C2 => 
                           n4511, A => n1989, ZN => n1980);
   U3596 : OAI22_X1 port map( A1 => n4845, A2 => n12404, B1 => n4846, B2 => 
                           n12398, ZN => n1989);
   U3597 : AOI221_X1 port map( B1 => n12531, B2 => n11766, C1 => n12525, C2 => 
                           n9948, A => n3187, ZN => n3186);
   U3598 : OAI22_X1 port map( A1 => n14216, A2 => n12519, B1 => n13430, B2 => 
                           n12513, ZN => n3187);
   U3599 : AOI221_X1 port map( B1 => n12531, B2 => n11767, C1 => n12525, C2 => 
                           n9947, A => n3168, ZN => n3167);
   U3600 : OAI22_X1 port map( A1 => n14328, A2 => n12519, B1 => n13429, B2 => 
                           n12513, ZN => n3168);
   U3601 : AOI221_X1 port map( B1 => n12531, B2 => n11768, C1 => n12525, C2 => 
                           n9946, A => n3149, ZN => n3148);
   U3602 : OAI22_X1 port map( A1 => n14327, A2 => n12519, B1 => n13428, B2 => 
                           n12513, ZN => n3149);
   U3603 : AOI221_X1 port map( B1 => n12531, B2 => n11769, C1 => n12525, C2 => 
                           n9945, A => n3130, ZN => n3129);
   U3604 : OAI22_X1 port map( A1 => n14326, A2 => n12519, B1 => n13427, B2 => 
                           n12513, ZN => n3130);
   U3605 : AOI221_X1 port map( B1 => n12531, B2 => n11770, C1 => n12525, C2 => 
                           n9944, A => n3111, ZN => n3110);
   U3606 : OAI22_X1 port map( A1 => n14325, A2 => n12519, B1 => n13426, B2 => 
                           n12513, ZN => n3111);
   U3607 : AOI221_X1 port map( B1 => n12531, B2 => n11771, C1 => n12525, C2 => 
                           n9943, A => n3092, ZN => n3091);
   U3608 : OAI22_X1 port map( A1 => n14324, A2 => n12519, B1 => n13425, B2 => 
                           n12513, ZN => n3092);
   U3609 : AOI221_X1 port map( B1 => n12531, B2 => n11772, C1 => n12525, C2 => 
                           n9942, A => n3073, ZN => n3072);
   U3610 : OAI22_X1 port map( A1 => n14311, A2 => n12519, B1 => n13424, B2 => 
                           n12513, ZN => n3073);
   U3611 : AOI221_X1 port map( B1 => n12531, B2 => n11773, C1 => n12525, C2 => 
                           n9941, A => n3054, ZN => n3053);
   U3612 : OAI22_X1 port map( A1 => n14310, A2 => n12519, B1 => n13423, B2 => 
                           n12513, ZN => n3054);
   U3613 : AOI221_X1 port map( B1 => n12531, B2 => n11774, C1 => n12525, C2 => 
                           n9940, A => n3035, ZN => n3034);
   U3614 : OAI22_X1 port map( A1 => n14323, A2 => n12519, B1 => n13422, B2 => 
                           n12513, ZN => n3035);
   U3615 : AOI221_X1 port map( B1 => n12531, B2 => n11775, C1 => n12525, C2 => 
                           n9939, A => n3016, ZN => n3015);
   U3616 : OAI22_X1 port map( A1 => n14309, A2 => n12519, B1 => n13421, B2 => 
                           n12513, ZN => n3016);
   U3617 : AOI221_X1 port map( B1 => n12531, B2 => n11776, C1 => n12525, C2 => 
                           n9938, A => n2997, ZN => n2996);
   U3618 : OAI22_X1 port map( A1 => n14308, A2 => n12519, B1 => n13420, B2 => 
                           n12513, ZN => n2997);
   U3619 : AOI221_X1 port map( B1 => n12531, B2 => n11777, C1 => n12525, C2 => 
                           n9937, A => n2978, ZN => n2977);
   U3620 : OAI22_X1 port map( A1 => n14307, A2 => n12519, B1 => n13419, B2 => 
                           n12513, ZN => n2978);
   U3621 : AOI221_X1 port map( B1 => n12532, B2 => n11778, C1 => n12526, C2 => 
                           n9936, A => n2959, ZN => n2958);
   U3622 : OAI22_X1 port map( A1 => n14306, A2 => n12520, B1 => n13418, B2 => 
                           n12514, ZN => n2959);
   U3623 : AOI221_X1 port map( B1 => n12532, B2 => n9999, C1 => n12526, C2 => 
                           n9935, A => n2940, ZN => n2939);
   U3624 : OAI22_X1 port map( A1 => n14305, A2 => n12520, B1 => n13417, B2 => 
                           n12514, ZN => n2940);
   U3625 : AOI221_X1 port map( B1 => n12532, B2 => n9998, C1 => n12526, C2 => 
                           n9934, A => n2921, ZN => n2920);
   U3626 : OAI22_X1 port map( A1 => n14304, A2 => n12520, B1 => n13416, B2 => 
                           n12514, ZN => n2921);
   U3627 : AOI221_X1 port map( B1 => n12532, B2 => n9997, C1 => n12526, C2 => 
                           n9933, A => n2902, ZN => n2901);
   U3628 : OAI22_X1 port map( A1 => n14303, A2 => n12520, B1 => n13415, B2 => 
                           n12514, ZN => n2902);
   U3629 : AOI221_X1 port map( B1 => n12532, B2 => n9996, C1 => n12526, C2 => 
                           n9932, A => n2883, ZN => n2882);
   U3630 : OAI22_X1 port map( A1 => n14302, A2 => n12520, B1 => n13414, B2 => 
                           n12514, ZN => n2883);
   U3631 : AOI221_X1 port map( B1 => n12532, B2 => n9995, C1 => n12526, C2 => 
                           n9931, A => n2864, ZN => n2863);
   U3632 : OAI22_X1 port map( A1 => n14301, A2 => n12520, B1 => n13413, B2 => 
                           n12514, ZN => n2864);
   U3633 : AOI221_X1 port map( B1 => n12532, B2 => n9994, C1 => n12526, C2 => 
                           n9930, A => n2845, ZN => n2844);
   U3634 : OAI22_X1 port map( A1 => n14300, A2 => n12520, B1 => n13412, B2 => 
                           n12514, ZN => n2845);
   U3635 : AOI221_X1 port map( B1 => n12532, B2 => n9993, C1 => n12526, C2 => 
                           n9929, A => n2826, ZN => n2825);
   U3636 : OAI22_X1 port map( A1 => n14299, A2 => n12520, B1 => n13411, B2 => 
                           n12514, ZN => n2826);
   U3637 : AOI221_X1 port map( B1 => n12532, B2 => n9992, C1 => n12526, C2 => 
                           n9928, A => n2807, ZN => n2806);
   U3638 : OAI22_X1 port map( A1 => n14298, A2 => n12520, B1 => n13410, B2 => 
                           n12514, ZN => n2807);
   U3639 : AOI221_X1 port map( B1 => n12532, B2 => n9991, C1 => n12526, C2 => 
                           n9927, A => n2788, ZN => n2787);
   U3640 : OAI22_X1 port map( A1 => n14297, A2 => n12520, B1 => n13409, B2 => 
                           n12514, ZN => n2788);
   U3641 : AOI221_X1 port map( B1 => n12532, B2 => n9990, C1 => n12526, C2 => 
                           n9926, A => n2769, ZN => n2768);
   U3642 : OAI22_X1 port map( A1 => n14296, A2 => n12520, B1 => n13408, B2 => 
                           n12514, ZN => n2769);
   U3643 : AOI221_X1 port map( B1 => n12532, B2 => n9989, C1 => n12526, C2 => 
                           n9925, A => n2750, ZN => n2749);
   U3644 : OAI22_X1 port map( A1 => n14295, A2 => n12520, B1 => n13407, B2 => 
                           n12514, ZN => n2750);
   U3645 : AOI221_X1 port map( B1 => n12533, B2 => n9988, C1 => n12527, C2 => 
                           n9924, A => n2731, ZN => n2730);
   U3646 : OAI22_X1 port map( A1 => n14294, A2 => n12521, B1 => n13406, B2 => 
                           n12515, ZN => n2731);
   U3647 : AOI221_X1 port map( B1 => n12533, B2 => n9987, C1 => n12527, C2 => 
                           n9923, A => n2712, ZN => n2711);
   U3648 : OAI22_X1 port map( A1 => n14293, A2 => n12521, B1 => n13405, B2 => 
                           n12515, ZN => n2712);
   U3649 : AOI221_X1 port map( B1 => n12533, B2 => n9986, C1 => n12527, C2 => 
                           n9922, A => n2693, ZN => n2692);
   U3650 : OAI22_X1 port map( A1 => n14292, A2 => n12521, B1 => n13404, B2 => 
                           n12515, ZN => n2693);
   U3651 : AOI221_X1 port map( B1 => n12533, B2 => n9985, C1 => n12527, C2 => 
                           n9921, A => n2674, ZN => n2673);
   U3652 : OAI22_X1 port map( A1 => n14291, A2 => n12521, B1 => n13403, B2 => 
                           n12515, ZN => n2674);
   U3653 : AOI221_X1 port map( B1 => n12533, B2 => n9984, C1 => n12527, C2 => 
                           n9920, A => n2655, ZN => n2654);
   U3654 : OAI22_X1 port map( A1 => n14290, A2 => n12521, B1 => n13402, B2 => 
                           n12515, ZN => n2655);
   U3655 : AOI221_X1 port map( B1 => n12533, B2 => n9983, C1 => n12527, C2 => 
                           n9919, A => n2636, ZN => n2635);
   U3656 : OAI22_X1 port map( A1 => n14289, A2 => n12521, B1 => n14322, B2 => 
                           n12515, ZN => n2636);
   U3657 : AOI221_X1 port map( B1 => n12533, B2 => n9982, C1 => n12527, C2 => 
                           n9918, A => n2617, ZN => n2616);
   U3658 : OAI22_X1 port map( A1 => n14456, A2 => n12521, B1 => n14321, B2 => 
                           n12515, ZN => n2617);
   U3659 : AOI221_X1 port map( B1 => n12533, B2 => n9981, C1 => n12527, C2 => 
                           n9917, A => n2598, ZN => n2597);
   U3660 : OAI22_X1 port map( A1 => n14455, A2 => n12521, B1 => n14320, B2 => 
                           n12515, ZN => n2598);
   U3661 : AOI221_X1 port map( B1 => n12533, B2 => n9980, C1 => n12527, C2 => 
                           n9916, A => n2579, ZN => n2578);
   U3662 : OAI22_X1 port map( A1 => n14454, A2 => n12521, B1 => n14319, B2 => 
                           n12515, ZN => n2579);
   U3663 : AOI221_X1 port map( B1 => n12533, B2 => n9979, C1 => n12527, C2 => 
                           n9915, A => n2560, ZN => n2559);
   U3664 : OAI22_X1 port map( A1 => n14453, A2 => n12521, B1 => n14318, B2 => 
                           n12515, ZN => n2560);
   U3665 : AOI221_X1 port map( B1 => n12533, B2 => n9978, C1 => n12527, C2 => 
                           n9914, A => n2541, ZN => n2540);
   U3666 : OAI22_X1 port map( A1 => n14452, A2 => n12521, B1 => n14317, B2 => 
                           n12515, ZN => n2541);
   U3667 : AOI221_X1 port map( B1 => n12533, B2 => n9977, C1 => n12527, C2 => 
                           n9913, A => n2522, ZN => n2521);
   U3668 : OAI22_X1 port map( A1 => n14451, A2 => n12521, B1 => n14316, B2 => 
                           n12515, ZN => n2522);
   U3669 : AOI221_X1 port map( B1 => n12534, B2 => n9976, C1 => n12528, C2 => 
                           n9912, A => n2503, ZN => n2502);
   U3670 : OAI22_X1 port map( A1 => n14450, A2 => n12522, B1 => n14315, B2 => 
                           n12516, ZN => n2503);
   U3671 : AOI221_X1 port map( B1 => n12534, B2 => n9975, C1 => n12528, C2 => 
                           n9911, A => n2484, ZN => n2483);
   U3672 : OAI22_X1 port map( A1 => n14449, A2 => n12522, B1 => n14314, B2 => 
                           n12516, ZN => n2484);
   U3673 : AOI221_X1 port map( B1 => n12534, B2 => n9974, C1 => n12528, C2 => 
                           n9910, A => n2465, ZN => n2464);
   U3674 : OAI22_X1 port map( A1 => n14448, A2 => n12522, B1 => n14313, B2 => 
                           n12516, ZN => n2465);
   U3675 : AOI221_X1 port map( B1 => n12534, B2 => n9973, C1 => n12528, C2 => 
                           n9909, A => n2446, ZN => n2445);
   U3676 : OAI22_X1 port map( A1 => n14447, A2 => n12522, B1 => n14312, B2 => 
                           n12516, ZN => n2446);
   U3677 : AOI221_X1 port map( B1 => n12534, B2 => n9972, C1 => n12528, C2 => 
                           n9908, A => n2427, ZN => n2426);
   U3678 : OAI22_X1 port map( A1 => n14446, A2 => n12522, B1 => n14432, B2 => 
                           n12516, ZN => n2427);
   U3679 : AOI221_X1 port map( B1 => n12534, B2 => n9971, C1 => n12528, C2 => 
                           n9907, A => n2408, ZN => n2407);
   U3680 : OAI22_X1 port map( A1 => n14445, A2 => n12522, B1 => n14431, B2 => 
                           n12516, ZN => n2408);
   U3681 : AOI221_X1 port map( B1 => n12534, B2 => n9970, C1 => n12528, C2 => 
                           n9906, A => n2389, ZN => n2388);
   U3682 : OAI22_X1 port map( A1 => n14444, A2 => n12522, B1 => n14430, B2 => 
                           n12516, ZN => n2389);
   U3683 : AOI221_X1 port map( B1 => n12534, B2 => n9969, C1 => n12528, C2 => 
                           n9905, A => n2370, ZN => n2369);
   U3684 : OAI22_X1 port map( A1 => n14443, A2 => n12522, B1 => n14429, B2 => 
                           n12516, ZN => n2370);
   U3685 : AOI221_X1 port map( B1 => n12534, B2 => n9968, C1 => n12528, C2 => 
                           n9904, A => n2351, ZN => n2350);
   U3686 : OAI22_X1 port map( A1 => n14442, A2 => n12522, B1 => n14428, B2 => 
                           n12516, ZN => n2351);
   U3687 : AOI221_X1 port map( B1 => n12534, B2 => n9967, C1 => n12528, C2 => 
                           n9903, A => n2332, ZN => n2331);
   U3688 : OAI22_X1 port map( A1 => n14441, A2 => n12522, B1 => n14427, B2 => 
                           n12516, ZN => n2332);
   U3689 : AOI221_X1 port map( B1 => n12534, B2 => n9966, C1 => n12528, C2 => 
                           n9902, A => n2313, ZN => n2312);
   U3690 : OAI22_X1 port map( A1 => n13401, A2 => n12522, B1 => n14426, B2 => 
                           n12516, ZN => n2313);
   U3691 : AOI221_X1 port map( B1 => n12534, B2 => n9965, C1 => n12528, C2 => 
                           n9901, A => n2294, ZN => n2293);
   U3692 : OAI22_X1 port map( A1 => n13400, A2 => n12522, B1 => n14425, B2 => 
                           n12516, ZN => n2294);
   U3693 : AOI221_X1 port map( B1 => n12535, B2 => n9964, C1 => n12529, C2 => 
                           n9900, A => n2275, ZN => n2274);
   U3694 : OAI22_X1 port map( A1 => n13399, A2 => n12523, B1 => n14424, B2 => 
                           n12517, ZN => n2275);
   U3695 : AOI221_X1 port map( B1 => n12535, B2 => n9963, C1 => n12529, C2 => 
                           n9899, A => n2256, ZN => n2255);
   U3696 : OAI22_X1 port map( A1 => n13398, A2 => n12523, B1 => n14423, B2 => 
                           n12517, ZN => n2256);
   U3697 : AOI221_X1 port map( B1 => n12535, B2 => n9962, C1 => n12529, C2 => 
                           n9898, A => n2237, ZN => n2236);
   U3698 : OAI22_X1 port map( A1 => n13397, A2 => n12523, B1 => n14422, B2 => 
                           n12517, ZN => n2237);
   U3699 : AOI221_X1 port map( B1 => n12535, B2 => n9961, C1 => n12529, C2 => 
                           n9897, A => n2218, ZN => n2217);
   U3700 : OAI22_X1 port map( A1 => n13396, A2 => n12523, B1 => n14421, B2 => 
                           n12517, ZN => n2218);
   U3701 : AOI221_X1 port map( B1 => n12535, B2 => n9960, C1 => n12529, C2 => 
                           n9896, A => n2199, ZN => n2198);
   U3702 : OAI22_X1 port map( A1 => n13395, A2 => n12523, B1 => n14420, B2 => 
                           n12517, ZN => n2199);
   U3703 : AOI221_X1 port map( B1 => n12535, B2 => n9959, C1 => n12529, C2 => 
                           n9895, A => n2180, ZN => n2179);
   U3704 : OAI22_X1 port map( A1 => n13394, A2 => n12523, B1 => n14419, B2 => 
                           n12517, ZN => n2180);
   U3705 : AOI221_X1 port map( B1 => n12535, B2 => n9958, C1 => n12529, C2 => 
                           n9894, A => n2161, ZN => n2160);
   U3706 : OAI22_X1 port map( A1 => n13393, A2 => n12523, B1 => n14418, B2 => 
                           n12517, ZN => n2161);
   U3707 : AOI221_X1 port map( B1 => n12535, B2 => n9957, C1 => n12529, C2 => 
                           n9893, A => n2142, ZN => n2141);
   U3708 : OAI22_X1 port map( A1 => n14440, A2 => n12523, B1 => n14417, B2 => 
                           n12517, ZN => n2142);
   U3709 : AOI221_X1 port map( B1 => n12535, B2 => n9956, C1 => n12529, C2 => 
                           n9892, A => n2123, ZN => n2122);
   U3710 : OAI22_X1 port map( A1 => n14439, A2 => n12523, B1 => n14416, B2 => 
                           n12517, ZN => n2123);
   U3711 : AOI221_X1 port map( B1 => n12535, B2 => n9955, C1 => n12529, C2 => 
                           n9891, A => n2104, ZN => n2103);
   U3712 : OAI22_X1 port map( A1 => n14438, A2 => n12523, B1 => n14415, B2 => 
                           n12517, ZN => n2104);
   U3713 : AOI221_X1 port map( B1 => n12535, B2 => n9954, C1 => n12529, C2 => 
                           n9890, A => n2085, ZN => n2084);
   U3714 : OAI22_X1 port map( A1 => n14437, A2 => n12523, B1 => n14414, B2 => 
                           n12517, ZN => n2085);
   U3715 : AOI221_X1 port map( B1 => n12535, B2 => n9953, C1 => n12529, C2 => 
                           n9889, A => n2066, ZN => n2065);
   U3716 : OAI22_X1 port map( A1 => n14436, A2 => n12523, B1 => n14413, B2 => 
                           n12517, ZN => n2066);
   U3717 : OAI22_X1 port map( A1 => n13122, A2 => n13242, B1 => n13112, B2 => 
                           n11959, ZN => n6806);
   U3718 : OAI22_X1 port map( A1 => n13122, A2 => n13245, B1 => n13112, B2 => 
                           n11960, ZN => n6807);
   U3719 : OAI22_X1 port map( A1 => n13122, A2 => n13248, B1 => n13112, B2 => 
                           n11961, ZN => n6808);
   U3720 : OAI22_X1 port map( A1 => n13122, A2 => n13251, B1 => n13112, B2 => 
                           n11962, ZN => n6809);
   U3721 : OAI22_X1 port map( A1 => n13122, A2 => n13254, B1 => n13112, B2 => 
                           n11963, ZN => n6810);
   U3722 : OAI22_X1 port map( A1 => n13121, A2 => n13257, B1 => n13112, B2 => 
                           n11964, ZN => n6811);
   U3723 : OAI22_X1 port map( A1 => n13121, A2 => n13260, B1 => n13112, B2 => 
                           n11965, ZN => n6812);
   U3724 : OAI22_X1 port map( A1 => n13121, A2 => n13263, B1 => n13112, B2 => 
                           n11966, ZN => n6813);
   U3725 : OAI22_X1 port map( A1 => n13121, A2 => n13266, B1 => n13112, B2 => 
                           n11967, ZN => n6814);
   U3726 : OAI22_X1 port map( A1 => n13121, A2 => n13269, B1 => n13112, B2 => 
                           n11968, ZN => n6815);
   U3727 : OAI22_X1 port map( A1 => n13120, A2 => n13272, B1 => n13112, B2 => 
                           n11969, ZN => n6816);
   U3728 : OAI22_X1 port map( A1 => n13120, A2 => n13275, B1 => n13112, B2 => 
                           n11970, ZN => n6817);
   U3729 : OAI22_X1 port map( A1 => n13120, A2 => n13278, B1 => n13112, B2 => 
                           n11971, ZN => n6818);
   U3730 : OAI22_X1 port map( A1 => n13120, A2 => n13281, B1 => n13113, B2 => 
                           n11972, ZN => n6819);
   U3731 : OAI22_X1 port map( A1 => n13120, A2 => n13284, B1 => n13113, B2 => 
                           n11973, ZN => n6820);
   U3732 : OAI22_X1 port map( A1 => n13119, A2 => n13287, B1 => n13113, B2 => 
                           n11974, ZN => n6821);
   U3733 : OAI22_X1 port map( A1 => n13119, A2 => n13290, B1 => n13113, B2 => 
                           n11975, ZN => n6822);
   U3734 : OAI22_X1 port map( A1 => n13119, A2 => n13293, B1 => n13113, B2 => 
                           n11976, ZN => n6823);
   U3735 : OAI22_X1 port map( A1 => n13119, A2 => n13296, B1 => n13113, B2 => 
                           n11977, ZN => n6824);
   U3736 : OAI22_X1 port map( A1 => n13119, A2 => n13299, B1 => n13113, B2 => 
                           n11978, ZN => n6825);
   U3737 : OAI22_X1 port map( A1 => n13118, A2 => n13302, B1 => n13113, B2 => 
                           n11979, ZN => n6826);
   U3738 : OAI22_X1 port map( A1 => n13118, A2 => n13305, B1 => n13113, B2 => 
                           n11980, ZN => n6827);
   U3739 : OAI22_X1 port map( A1 => n13118, A2 => n13308, B1 => n13113, B2 => 
                           n11981, ZN => n6828);
   U3740 : OAI22_X1 port map( A1 => n13118, A2 => n13311, B1 => n13113, B2 => 
                           n11982, ZN => n6829);
   U3741 : OAI22_X1 port map( A1 => n13118, A2 => n13314, B1 => n13113, B2 => 
                           n11983, ZN => n6830);
   U3742 : OAI22_X1 port map( A1 => n13117, A2 => n13317, B1 => n13113, B2 => 
                           n11984, ZN => n6831);
   U3743 : OAI22_X1 port map( A1 => n13117, A2 => n13320, B1 => n13114, B2 => 
                           n11985, ZN => n6832);
   U3744 : OAI22_X1 port map( A1 => n13117, A2 => n13323, B1 => n13114, B2 => 
                           n11986, ZN => n6833);
   U3745 : OAI22_X1 port map( A1 => n13117, A2 => n13326, B1 => n13114, B2 => 
                           n11987, ZN => n6834);
   U3746 : OAI22_X1 port map( A1 => n13117, A2 => n13329, B1 => n13114, B2 => 
                           n11988, ZN => n6835);
   U3747 : OAI22_X1 port map( A1 => n13116, A2 => n13332, B1 => n13114, B2 => 
                           n11989, ZN => n6836);
   U3748 : OAI22_X1 port map( A1 => n13116, A2 => n13335, B1 => n13114, B2 => 
                           n11990, ZN => n6837);
   U3749 : OAI22_X1 port map( A1 => n13116, A2 => n13338, B1 => n13114, B2 => 
                           n11991, ZN => n6838);
   U3750 : OAI22_X1 port map( A1 => n13116, A2 => n13341, B1 => n13114, B2 => 
                           n11992, ZN => n6839);
   U3751 : OAI22_X1 port map( A1 => n13116, A2 => n13344, B1 => n13114, B2 => 
                           n11993, ZN => n6840);
   U3752 : OAI22_X1 port map( A1 => n13115, A2 => n13347, B1 => n13114, B2 => 
                           n11994, ZN => n6841);
   U3753 : OAI22_X1 port map( A1 => n13115, A2 => n13350, B1 => n13114, B2 => 
                           n11995, ZN => n6842);
   U3754 : OAI22_X1 port map( A1 => n13115, A2 => n13353, B1 => n13114, B2 => 
                           n11996, ZN => n6843);
   U3755 : OAI22_X1 port map( A1 => n13115, A2 => n13356, B1 => n13114, B2 => 
                           n11997, ZN => n6844);
   U3756 : OAI22_X1 port map( A1 => n13147, A2 => n13173, B1 => n13133, B2 => 
                           n11779, ZN => n6847);
   U3757 : OAI22_X1 port map( A1 => n13147, A2 => n13176, B1 => n13134, B2 => 
                           n11780, ZN => n6848);
   U3758 : OAI22_X1 port map( A1 => n13147, A2 => n13179, B1 => n13131, B2 => 
                           n11781, ZN => n6849);
   U3759 : OAI22_X1 port map( A1 => n13146, A2 => n13182, B1 => n13133, B2 => 
                           n11782, ZN => n6850);
   U3760 : OAI22_X1 port map( A1 => n13146, A2 => n13185, B1 => n13134, B2 => 
                           n11783, ZN => n6851);
   U3761 : OAI22_X1 port map( A1 => n13146, A2 => n13188, B1 => n13130, B2 => 
                           n11784, ZN => n6852);
   U3762 : OAI22_X1 port map( A1 => n13146, A2 => n13191, B1 => n1910, B2 => 
                           n11785, ZN => n6853);
   U3763 : OAI22_X1 port map( A1 => n13146, A2 => n13194, B1 => n1910, B2 => 
                           n11786, ZN => n6854);
   U3764 : OAI22_X1 port map( A1 => n13145, A2 => n13197, B1 => n1910, B2 => 
                           n11787, ZN => n6855);
   U3765 : OAI22_X1 port map( A1 => n13145, A2 => n13200, B1 => n1910, B2 => 
                           n11788, ZN => n6856);
   U3766 : OAI22_X1 port map( A1 => n13145, A2 => n13203, B1 => n1910, B2 => 
                           n11789, ZN => n6857);
   U3767 : OAI22_X1 port map( A1 => n13145, A2 => n13206, B1 => n13131, B2 => 
                           n11790, ZN => n6858);
   U3768 : OAI22_X1 port map( A1 => n13145, A2 => n13209, B1 => n13131, B2 => 
                           n11791, ZN => n6859);
   U3769 : OAI22_X1 port map( A1 => n13144, A2 => n13212, B1 => n13131, B2 => 
                           n11792, ZN => n6860);
   U3770 : OAI22_X1 port map( A1 => n13144, A2 => n13215, B1 => n13131, B2 => 
                           n11793, ZN => n6861);
   U3771 : OAI22_X1 port map( A1 => n13144, A2 => n13218, B1 => n13131, B2 => 
                           n11794, ZN => n6862);
   U3772 : OAI22_X1 port map( A1 => n13144, A2 => n13221, B1 => n13131, B2 => 
                           n11795, ZN => n6863);
   U3773 : OAI22_X1 port map( A1 => n13144, A2 => n13224, B1 => n13131, B2 => 
                           n11796, ZN => n6864);
   U3774 : OAI22_X1 port map( A1 => n13143, A2 => n13227, B1 => n13131, B2 => 
                           n11797, ZN => n6865);
   U3775 : OAI22_X1 port map( A1 => n13143, A2 => n13230, B1 => n13131, B2 => 
                           n11798, ZN => n6866);
   U3776 : OAI22_X1 port map( A1 => n13143, A2 => n13233, B1 => n13131, B2 => 
                           n11799, ZN => n6867);
   U3777 : OAI22_X1 port map( A1 => n13143, A2 => n13236, B1 => n13131, B2 => 
                           n11800, ZN => n6868);
   U3778 : OAI22_X1 port map( A1 => n13143, A2 => n13239, B1 => n13131, B2 => 
                           n11801, ZN => n6869);
   U3779 : OAI22_X1 port map( A1 => n13147, A2 => n13170, B1 => n1910, B2 => 
                           n11802, ZN => n6846);
   U3780 : OAI22_X1 port map( A1 => n12804, A2 => n13219, B1 => n12791, B2 => 
                           n11803, ZN => n5774);
   U3781 : OAI22_X1 port map( A1 => n12806, A2 => n13183, B1 => n12793, B2 => 
                           n11804, ZN => n5762);
   U3782 : OAI22_X1 port map( A1 => n12806, A2 => n13186, B1 => n12794, B2 => 
                           n11805, ZN => n5763);
   U3783 : OAI22_X1 port map( A1 => n12806, A2 => n13189, B1 => n12791, B2 => 
                           n11806, ZN => n5764);
   U3784 : OAI22_X1 port map( A1 => n12806, A2 => n13192, B1 => n12793, B2 => 
                           n11807, ZN => n5765);
   U3785 : OAI22_X1 port map( A1 => n12805, A2 => n13198, B1 => n12794, B2 => 
                           n11808, ZN => n5767);
   U3786 : OAI22_X1 port map( A1 => n12805, A2 => n13201, B1 => n12790, B2 => 
                           n11809, ZN => n5768);
   U3787 : OAI22_X1 port map( A1 => n12805, A2 => n13204, B1 => n1936, B2 => 
                           n11810, ZN => n5769);
   U3788 : OAI22_X1 port map( A1 => n12726, A2 => n13183, B1 => n12712, B2 => 
                           n11811, ZN => n5506);
   U3789 : OAI22_X1 port map( A1 => n12726, A2 => n13186, B1 => n12714, B2 => 
                           n11812, ZN => n5507);
   U3790 : OAI22_X1 port map( A1 => n12726, A2 => n13189, B1 => n12711, B2 => 
                           n11813, ZN => n5508);
   U3791 : OAI22_X1 port map( A1 => n12726, A2 => n13192, B1 => n12712, B2 => 
                           n11814, ZN => n5509);
   U3792 : OAI22_X1 port map( A1 => n12726, A2 => n13195, B1 => n12714, B2 => 
                           n11815, ZN => n5510);
   U3793 : OAI22_X1 port map( A1 => n12725, A2 => n13198, B1 => n12710, B2 => 
                           n11816, ZN => n5511);
   U3794 : OAI22_X1 port map( A1 => n12725, A2 => n13201, B1 => n1940, B2 => 
                           n11817, ZN => n5512);
   U3795 : OAI22_X1 port map( A1 => n12725, A2 => n13204, B1 => n1940, B2 => 
                           n11818, ZN => n5513);
   U3796 : OAI22_X1 port map( A1 => n12725, A2 => n13207, B1 => n12711, B2 => 
                           n11819, ZN => n5514);
   U3797 : OAI22_X1 port map( A1 => n12725, A2 => n13210, B1 => n12711, B2 => 
                           n11820, ZN => n5515);
   U3798 : OAI22_X1 port map( A1 => n12806, A2 => n13195, B1 => n1936, B2 => 
                           n11821, ZN => n5766);
   U3799 : OAI22_X1 port map( A1 => n12805, A2 => n13207, B1 => n12791, B2 => 
                           n11822, ZN => n5770);
   U3800 : OAI22_X1 port map( A1 => n12805, A2 => n13210, B1 => n12791, B2 => 
                           n11823, ZN => n5771);
   U3801 : OAI22_X1 port map( A1 => n12804, A2 => n13213, B1 => n12791, B2 => 
                           n11824, ZN => n5772);
   U3802 : OAI22_X1 port map( A1 => n12804, A2 => n13216, B1 => n12791, B2 => 
                           n11825, ZN => n5773);
   U3803 : OAI22_X1 port map( A1 => n12804, A2 => n13222, B1 => n12791, B2 => 
                           n11826, ZN => n5775);
   U3804 : OAI22_X1 port map( A1 => n12804, A2 => n13225, B1 => n12791, B2 => 
                           n11827, ZN => n5776);
   U3805 : OAI22_X1 port map( A1 => n12803, A2 => n13228, B1 => n12791, B2 => 
                           n11828, ZN => n5777);
   U3806 : OAI22_X1 port map( A1 => n12803, A2 => n13231, B1 => n12791, B2 => 
                           n11829, ZN => n5778);
   U3807 : OAI22_X1 port map( A1 => n12803, A2 => n13234, B1 => n12791, B2 => 
                           n11830, ZN => n5779);
   U3808 : OAI22_X1 port map( A1 => n12803, A2 => n13237, B1 => n12791, B2 => 
                           n11831, ZN => n5780);
   U3809 : OAI22_X1 port map( A1 => n12803, A2 => n13240, B1 => n12791, B2 => 
                           n11832, ZN => n5781);
   U3810 : OAI22_X1 port map( A1 => n12724, A2 => n13213, B1 => n12711, B2 => 
                           n11833, ZN => n5516);
   U3811 : OAI22_X1 port map( A1 => n12724, A2 => n13216, B1 => n12711, B2 => 
                           n11834, ZN => n5517);
   U3812 : OAI22_X1 port map( A1 => n12724, A2 => n13219, B1 => n12711, B2 => 
                           n11835, ZN => n5518);
   U3813 : OAI22_X1 port map( A1 => n12724, A2 => n13222, B1 => n12711, B2 => 
                           n11836, ZN => n5519);
   U3814 : OAI22_X1 port map( A1 => n12724, A2 => n13225, B1 => n12711, B2 => 
                           n11837, ZN => n5520);
   U3815 : OAI22_X1 port map( A1 => n12723, A2 => n13228, B1 => n12711, B2 => 
                           n11838, ZN => n5521);
   U3816 : OAI22_X1 port map( A1 => n12723, A2 => n13231, B1 => n12711, B2 => 
                           n11839, ZN => n5522);
   U3817 : OAI22_X1 port map( A1 => n12723, A2 => n13234, B1 => n12711, B2 => 
                           n11840, ZN => n5523);
   U3818 : OAI22_X1 port map( A1 => n12723, A2 => n13237, B1 => n12711, B2 => 
                           n11841, ZN => n5524);
   U3819 : OAI22_X1 port map( A1 => n12723, A2 => n13240, B1 => n12711, B2 => 
                           n11842, ZN => n5525);
   U3820 : OAI22_X1 port map( A1 => n12727, A2 => n13171, B1 => n1940, B2 => 
                           n11843, ZN => n5502);
   U3821 : OAI22_X1 port map( A1 => n12727, A2 => n13174, B1 => n1940, B2 => 
                           n11844, ZN => n5503);
   U3822 : OAI22_X1 port map( A1 => n12727, A2 => n13177, B1 => n1940, B2 => 
                           n11845, ZN => n5504);
   U3823 : OAI22_X1 port map( A1 => n12727, A2 => n13180, B1 => n1940, B2 => 
                           n11846, ZN => n5505);
   U3824 : OAI22_X1 port map( A1 => n12747, A2 => n13171, B1 => n12731, B2 => 
                           n11998, ZN => n5566);
   U3825 : OAI22_X1 port map( A1 => n12747, A2 => n13174, B1 => n12731, B2 => 
                           n11999, ZN => n5567);
   U3826 : OAI22_X1 port map( A1 => n12747, A2 => n13177, B1 => n12731, B2 => 
                           n12000, ZN => n5568);
   U3827 : OAI22_X1 port map( A1 => n12747, A2 => n13180, B1 => n12731, B2 => 
                           n12001, ZN => n5569);
   U3828 : OAI22_X1 port map( A1 => n12746, A2 => n13183, B1 => n12731, B2 => 
                           n12002, ZN => n5570);
   U3829 : OAI22_X1 port map( A1 => n12746, A2 => n13186, B1 => n12731, B2 => 
                           n12003, ZN => n5571);
   U3830 : OAI22_X1 port map( A1 => n12746, A2 => n13189, B1 => n12731, B2 => 
                           n12004, ZN => n5572);
   U3831 : OAI22_X1 port map( A1 => n12746, A2 => n13192, B1 => n12731, B2 => 
                           n12005, ZN => n5573);
   U3832 : OAI22_X1 port map( A1 => n12746, A2 => n13195, B1 => n12731, B2 => 
                           n12006, ZN => n5574);
   U3833 : OAI22_X1 port map( A1 => n12745, A2 => n13198, B1 => n12731, B2 => 
                           n12007, ZN => n5575);
   U3834 : OAI22_X1 port map( A1 => n12745, A2 => n13201, B1 => n12731, B2 => 
                           n12008, ZN => n5576);
   U3835 : OAI22_X1 port map( A1 => n12745, A2 => n13204, B1 => n12731, B2 => 
                           n12009, ZN => n5577);
   U3836 : OAI22_X1 port map( A1 => n12745, A2 => n13207, B1 => n12733, B2 => 
                           n12010, ZN => n5578);
   U3837 : OAI22_X1 port map( A1 => n12745, A2 => n13210, B1 => n12734, B2 => 
                           n12011, ZN => n5579);
   U3838 : OAI22_X1 port map( A1 => n12744, A2 => n13213, B1 => n12731, B2 => 
                           n12012, ZN => n5580);
   U3839 : OAI22_X1 port map( A1 => n12744, A2 => n13216, B1 => n12733, B2 => 
                           n12013, ZN => n5581);
   U3840 : OAI22_X1 port map( A1 => n12744, A2 => n13219, B1 => n12734, B2 => 
                           n12014, ZN => n5582);
   U3841 : OAI22_X1 port map( A1 => n12744, A2 => n13222, B1 => n12730, B2 => 
                           n12015, ZN => n5583);
   U3842 : OAI22_X1 port map( A1 => n12744, A2 => n13225, B1 => n1939, B2 => 
                           n12016, ZN => n5584);
   U3843 : OAI22_X1 port map( A1 => n12743, A2 => n13228, B1 => n1939, B2 => 
                           n12017, ZN => n5585);
   U3844 : OAI22_X1 port map( A1 => n12743, A2 => n13231, B1 => n1939, B2 => 
                           n12018, ZN => n5586);
   U3845 : OAI22_X1 port map( A1 => n12743, A2 => n13234, B1 => n1939, B2 => 
                           n12019, ZN => n5587);
   U3846 : OAI22_X1 port map( A1 => n12743, A2 => n13237, B1 => n1939, B2 => 
                           n12020, ZN => n5588);
   U3847 : OAI22_X1 port map( A1 => n12743, A2 => n13240, B1 => n1939, B2 => 
                           n12021, ZN => n5589);
   U3848 : OAI22_X1 port map( A1 => n12807, A2 => n13171, B1 => n1936, B2 => 
                           n11847, ZN => n5758);
   U3849 : OAI22_X1 port map( A1 => n12807, A2 => n13174, B1 => n1936, B2 => 
                           n11848, ZN => n5759);
   U3850 : OAI22_X1 port map( A1 => n12807, A2 => n13177, B1 => n1936, B2 => 
                           n11849, ZN => n5760);
   U3851 : OAI22_X1 port map( A1 => n12807, A2 => n13180, B1 => n1936, B2 => 
                           n11850, ZN => n5761);
   U3852 : OAI22_X1 port map( A1 => n12827, A2 => n13171, B1 => n12811, B2 => 
                           n12022, ZN => n5822);
   U3853 : OAI22_X1 port map( A1 => n12827, A2 => n13174, B1 => n12811, B2 => 
                           n12023, ZN => n5823);
   U3854 : OAI22_X1 port map( A1 => n12827, A2 => n13177, B1 => n12811, B2 => 
                           n12024, ZN => n5824);
   U3855 : OAI22_X1 port map( A1 => n12827, A2 => n13180, B1 => n12811, B2 => 
                           n12025, ZN => n5825);
   U3856 : OAI22_X1 port map( A1 => n12826, A2 => n13183, B1 => n12811, B2 => 
                           n12026, ZN => n5826);
   U3857 : OAI22_X1 port map( A1 => n12826, A2 => n13186, B1 => n12811, B2 => 
                           n12027, ZN => n5827);
   U3858 : OAI22_X1 port map( A1 => n12826, A2 => n13189, B1 => n12811, B2 => 
                           n12028, ZN => n5828);
   U3859 : OAI22_X1 port map( A1 => n12826, A2 => n13192, B1 => n12811, B2 => 
                           n12029, ZN => n5829);
   U3860 : OAI22_X1 port map( A1 => n12826, A2 => n13195, B1 => n12811, B2 => 
                           n12030, ZN => n5830);
   U3861 : OAI22_X1 port map( A1 => n12825, A2 => n13198, B1 => n12811, B2 => 
                           n12031, ZN => n5831);
   U3862 : OAI22_X1 port map( A1 => n12825, A2 => n13201, B1 => n12811, B2 => 
                           n12032, ZN => n5832);
   U3863 : OAI22_X1 port map( A1 => n12825, A2 => n13204, B1 => n12811, B2 => 
                           n12033, ZN => n5833);
   U3864 : OAI22_X1 port map( A1 => n12825, A2 => n13207, B1 => n12813, B2 => 
                           n12034, ZN => n5834);
   U3865 : OAI22_X1 port map( A1 => n12825, A2 => n13210, B1 => n12814, B2 => 
                           n12035, ZN => n5835);
   U3866 : OAI22_X1 port map( A1 => n12824, A2 => n13213, B1 => n12811, B2 => 
                           n12036, ZN => n5836);
   U3867 : OAI22_X1 port map( A1 => n12824, A2 => n13216, B1 => n12813, B2 => 
                           n12037, ZN => n5837);
   U3868 : OAI22_X1 port map( A1 => n12824, A2 => n13219, B1 => n12814, B2 => 
                           n12038, ZN => n5838);
   U3869 : OAI22_X1 port map( A1 => n12824, A2 => n13222, B1 => n12810, B2 => 
                           n12039, ZN => n5839);
   U3870 : OAI22_X1 port map( A1 => n12824, A2 => n13225, B1 => n1935, B2 => 
                           n12040, ZN => n5840);
   U3871 : OAI22_X1 port map( A1 => n12823, A2 => n13228, B1 => n1935, B2 => 
                           n12041, ZN => n5841);
   U3872 : OAI22_X1 port map( A1 => n12823, A2 => n13231, B1 => n1935, B2 => 
                           n12042, ZN => n5842);
   U3873 : OAI22_X1 port map( A1 => n12823, A2 => n13234, B1 => n1935, B2 => 
                           n12043, ZN => n5843);
   U3874 : OAI22_X1 port map( A1 => n12823, A2 => n13237, B1 => n1935, B2 => 
                           n12044, ZN => n5844);
   U3875 : OAI22_X1 port map( A1 => n12823, A2 => n13240, B1 => n1935, B2 => 
                           n12045, ZN => n5845);
   U3876 : OAI22_X1 port map( A1 => n13125, A2 => n13209, B1 => n13111, B2 => 
                           n12046, ZN => n6795);
   U3877 : OAI22_X1 port map( A1 => n13124, A2 => n13212, B1 => n13111, B2 => 
                           n12047, ZN => n6796);
   U3878 : OAI22_X1 port map( A1 => n13124, A2 => n13215, B1 => n13111, B2 => 
                           n12048, ZN => n6797);
   U3879 : OAI22_X1 port map( A1 => n13124, A2 => n13218, B1 => n13111, B2 => 
                           n12049, ZN => n6798);
   U3880 : OAI22_X1 port map( A1 => n13124, A2 => n13221, B1 => n13111, B2 => 
                           n12050, ZN => n6799);
   U3881 : OAI22_X1 port map( A1 => n13124, A2 => n13224, B1 => n13111, B2 => 
                           n12051, ZN => n6800);
   U3882 : OAI22_X1 port map( A1 => n13123, A2 => n13227, B1 => n13111, B2 => 
                           n12052, ZN => n6801);
   U3883 : OAI22_X1 port map( A1 => n13123, A2 => n13230, B1 => n13111, B2 => 
                           n12053, ZN => n6802);
   U3884 : OAI22_X1 port map( A1 => n13123, A2 => n13233, B1 => n13111, B2 => 
                           n12054, ZN => n6803);
   U3885 : OAI22_X1 port map( A1 => n13123, A2 => n13236, B1 => n13111, B2 => 
                           n12055, ZN => n6804);
   U3886 : OAI22_X1 port map( A1 => n13123, A2 => n13239, B1 => n13111, B2 => 
                           n12056, ZN => n6805);
   U3887 : OAI22_X1 port map( A1 => n13142, A2 => n13242, B1 => n13132, B2 => 
                           n11851, ZN => n6870);
   U3888 : OAI22_X1 port map( A1 => n13142, A2 => n13245, B1 => n13132, B2 => 
                           n11852, ZN => n6871);
   U3889 : OAI22_X1 port map( A1 => n13142, A2 => n13248, B1 => n13132, B2 => 
                           n11853, ZN => n6872);
   U3890 : OAI22_X1 port map( A1 => n13142, A2 => n13251, B1 => n13132, B2 => 
                           n11854, ZN => n6873);
   U3891 : OAI22_X1 port map( A1 => n13142, A2 => n13254, B1 => n13132, B2 => 
                           n11855, ZN => n6874);
   U3892 : OAI22_X1 port map( A1 => n13141, A2 => n13257, B1 => n13132, B2 => 
                           n11856, ZN => n6875);
   U3893 : OAI22_X1 port map( A1 => n13141, A2 => n13260, B1 => n13132, B2 => 
                           n11857, ZN => n6876);
   U3894 : OAI22_X1 port map( A1 => n13141, A2 => n13263, B1 => n13132, B2 => 
                           n11858, ZN => n6877);
   U3895 : OAI22_X1 port map( A1 => n13141, A2 => n13266, B1 => n13132, B2 => 
                           n11859, ZN => n6878);
   U3896 : OAI22_X1 port map( A1 => n13141, A2 => n13269, B1 => n13132, B2 => 
                           n11860, ZN => n6879);
   U3897 : OAI22_X1 port map( A1 => n13140, A2 => n13272, B1 => n13132, B2 => 
                           n11861, ZN => n6880);
   U3898 : OAI22_X1 port map( A1 => n13140, A2 => n13275, B1 => n13132, B2 => 
                           n11862, ZN => n6881);
   U3899 : OAI22_X1 port map( A1 => n13140, A2 => n13278, B1 => n13133, B2 => 
                           n11863, ZN => n6882);
   U3900 : OAI22_X1 port map( A1 => n13140, A2 => n13281, B1 => n13133, B2 => 
                           n11864, ZN => n6883);
   U3901 : OAI22_X1 port map( A1 => n13140, A2 => n13284, B1 => n13133, B2 => 
                           n11865, ZN => n6884);
   U3902 : OAI22_X1 port map( A1 => n13139, A2 => n13287, B1 => n13133, B2 => 
                           n11866, ZN => n6885);
   U3903 : OAI22_X1 port map( A1 => n13139, A2 => n13290, B1 => n13133, B2 => 
                           n11867, ZN => n6886);
   U3904 : OAI22_X1 port map( A1 => n13139, A2 => n13293, B1 => n13133, B2 => 
                           n11868, ZN => n6887);
   U3905 : OAI22_X1 port map( A1 => n13139, A2 => n13296, B1 => n13133, B2 => 
                           n11869, ZN => n6888);
   U3906 : OAI22_X1 port map( A1 => n13139, A2 => n13299, B1 => n13133, B2 => 
                           n11870, ZN => n6889);
   U3907 : OAI22_X1 port map( A1 => n13138, A2 => n13302, B1 => n13133, B2 => 
                           n11871, ZN => n6890);
   U3908 : OAI22_X1 port map( A1 => n13138, A2 => n13305, B1 => n13133, B2 => 
                           n11872, ZN => n6891);
   U3909 : OAI22_X1 port map( A1 => n13138, A2 => n13308, B1 => n13133, B2 => 
                           n11873, ZN => n6892);
   U3910 : OAI22_X1 port map( A1 => n13138, A2 => n13311, B1 => n13133, B2 => 
                           n11874, ZN => n6893);
   U3911 : OAI22_X1 port map( A1 => n13138, A2 => n13314, B1 => n13134, B2 => 
                           n11875, ZN => n6894);
   U3912 : OAI22_X1 port map( A1 => n13137, A2 => n13317, B1 => n13134, B2 => 
                           n11876, ZN => n6895);
   U3913 : OAI22_X1 port map( A1 => n13137, A2 => n13320, B1 => n13134, B2 => 
                           n11877, ZN => n6896);
   U3914 : OAI22_X1 port map( A1 => n13137, A2 => n13323, B1 => n13134, B2 => 
                           n11878, ZN => n6897);
   U3915 : OAI22_X1 port map( A1 => n13137, A2 => n13326, B1 => n13134, B2 => 
                           n11879, ZN => n6898);
   U3916 : OAI22_X1 port map( A1 => n13137, A2 => n13329, B1 => n13134, B2 => 
                           n11880, ZN => n6899);
   U3917 : OAI22_X1 port map( A1 => n13136, A2 => n13332, B1 => n13134, B2 => 
                           n11881, ZN => n6900);
   U3918 : OAI22_X1 port map( A1 => n13136, A2 => n13335, B1 => n13134, B2 => 
                           n11882, ZN => n6901);
   U3919 : OAI22_X1 port map( A1 => n13136, A2 => n13338, B1 => n13134, B2 => 
                           n11883, ZN => n6902);
   U3920 : OAI22_X1 port map( A1 => n13136, A2 => n13341, B1 => n13134, B2 => 
                           n11884, ZN => n6903);
   U3921 : OAI22_X1 port map( A1 => n13136, A2 => n13344, B1 => n13134, B2 => 
                           n11885, ZN => n6904);
   U3922 : OAI22_X1 port map( A1 => n13135, A2 => n13347, B1 => n13134, B2 => 
                           n11886, ZN => n6905);
   U3923 : OAI22_X1 port map( A1 => n12802, A2 => n13243, B1 => n12792, B2 => 
                           n11887, ZN => n5782);
   U3924 : OAI22_X1 port map( A1 => n12802, A2 => n13246, B1 => n12792, B2 => 
                           n11888, ZN => n5783);
   U3925 : OAI22_X1 port map( A1 => n12802, A2 => n13249, B1 => n12792, B2 => 
                           n11889, ZN => n5784);
   U3926 : OAI22_X1 port map( A1 => n12802, A2 => n13252, B1 => n12792, B2 => 
                           n11890, ZN => n5785);
   U3927 : OAI22_X1 port map( A1 => n12802, A2 => n13255, B1 => n12792, B2 => 
                           n11891, ZN => n5786);
   U3928 : OAI22_X1 port map( A1 => n12801, A2 => n13258, B1 => n12792, B2 => 
                           n11892, ZN => n5787);
   U3929 : OAI22_X1 port map( A1 => n12801, A2 => n13261, B1 => n12792, B2 => 
                           n11893, ZN => n5788);
   U3930 : OAI22_X1 port map( A1 => n12801, A2 => n13264, B1 => n12792, B2 => 
                           n11894, ZN => n5789);
   U3931 : OAI22_X1 port map( A1 => n12801, A2 => n13267, B1 => n12792, B2 => 
                           n11895, ZN => n5790);
   U3932 : OAI22_X1 port map( A1 => n12801, A2 => n13270, B1 => n12792, B2 => 
                           n11896, ZN => n5791);
   U3933 : OAI22_X1 port map( A1 => n12800, A2 => n13273, B1 => n12792, B2 => 
                           n11897, ZN => n5792);
   U3934 : OAI22_X1 port map( A1 => n12800, A2 => n13276, B1 => n12792, B2 => 
                           n11898, ZN => n5793);
   U3935 : OAI22_X1 port map( A1 => n12800, A2 => n13279, B1 => n12793, B2 => 
                           n11899, ZN => n5794);
   U3936 : OAI22_X1 port map( A1 => n12800, A2 => n13282, B1 => n12793, B2 => 
                           n11900, ZN => n5795);
   U3937 : OAI22_X1 port map( A1 => n12800, A2 => n13285, B1 => n12793, B2 => 
                           n11901, ZN => n5796);
   U3938 : OAI22_X1 port map( A1 => n12799, A2 => n13288, B1 => n12793, B2 => 
                           n11902, ZN => n5797);
   U3939 : OAI22_X1 port map( A1 => n12799, A2 => n13291, B1 => n12793, B2 => 
                           n11903, ZN => n5798);
   U3940 : OAI22_X1 port map( A1 => n12799, A2 => n13294, B1 => n12793, B2 => 
                           n11904, ZN => n5799);
   U3941 : OAI22_X1 port map( A1 => n12799, A2 => n13297, B1 => n12793, B2 => 
                           n11905, ZN => n5800);
   U3942 : OAI22_X1 port map( A1 => n12799, A2 => n13300, B1 => n12793, B2 => 
                           n11906, ZN => n5801);
   U3943 : OAI22_X1 port map( A1 => n12798, A2 => n13303, B1 => n12793, B2 => 
                           n11907, ZN => n5802);
   U3944 : OAI22_X1 port map( A1 => n12798, A2 => n13306, B1 => n12793, B2 => 
                           n11908, ZN => n5803);
   U3945 : OAI22_X1 port map( A1 => n12798, A2 => n13309, B1 => n12793, B2 => 
                           n11909, ZN => n5804);
   U3946 : OAI22_X1 port map( A1 => n12722, A2 => n13249, B1 => n12712, B2 => 
                           n11910, ZN => n5528);
   U3947 : OAI22_X1 port map( A1 => n12722, A2 => n13252, B1 => n12712, B2 => 
                           n11911, ZN => n5529);
   U3948 : OAI22_X1 port map( A1 => n12722, A2 => n13255, B1 => n12712, B2 => 
                           n11912, ZN => n5530);
   U3949 : OAI22_X1 port map( A1 => n12721, A2 => n13258, B1 => n12712, B2 => 
                           n11913, ZN => n5531);
   U3950 : OAI22_X1 port map( A1 => n12721, A2 => n13261, B1 => n12712, B2 => 
                           n11914, ZN => n5532);
   U3951 : OAI22_X1 port map( A1 => n12721, A2 => n13264, B1 => n12712, B2 => 
                           n11915, ZN => n5533);
   U3952 : OAI22_X1 port map( A1 => n12721, A2 => n13267, B1 => n12712, B2 => 
                           n11916, ZN => n5534);
   U3953 : OAI22_X1 port map( A1 => n12721, A2 => n13270, B1 => n12712, B2 => 
                           n11917, ZN => n5535);
   U3954 : OAI22_X1 port map( A1 => n12720, A2 => n13273, B1 => n12712, B2 => 
                           n11918, ZN => n5536);
   U3955 : OAI22_X1 port map( A1 => n12720, A2 => n13276, B1 => n12712, B2 => 
                           n11919, ZN => n5537);
   U3956 : OAI22_X1 port map( A1 => n12720, A2 => n13279, B1 => n12713, B2 => 
                           n11920, ZN => n5538);
   U3957 : OAI22_X1 port map( A1 => n12720, A2 => n13282, B1 => n12713, B2 => 
                           n11921, ZN => n5539);
   U3958 : OAI22_X1 port map( A1 => n12720, A2 => n13285, B1 => n12713, B2 => 
                           n11922, ZN => n5540);
   U3959 : OAI22_X1 port map( A1 => n12719, A2 => n13288, B1 => n12713, B2 => 
                           n11923, ZN => n5541);
   U3960 : OAI22_X1 port map( A1 => n12719, A2 => n13291, B1 => n12713, B2 => 
                           n11924, ZN => n5542);
   U3961 : OAI22_X1 port map( A1 => n12719, A2 => n13294, B1 => n12713, B2 => 
                           n11925, ZN => n5543);
   U3962 : OAI22_X1 port map( A1 => n12719, A2 => n13297, B1 => n12713, B2 => 
                           n11926, ZN => n5544);
   U3963 : OAI22_X1 port map( A1 => n12719, A2 => n13300, B1 => n12713, B2 => 
                           n11927, ZN => n5545);
   U3964 : OAI22_X1 port map( A1 => n12718, A2 => n13303, B1 => n12713, B2 => 
                           n11928, ZN => n5546);
   U3965 : OAI22_X1 port map( A1 => n12718, A2 => n13306, B1 => n12713, B2 => 
                           n11929, ZN => n5547);
   U3966 : OAI22_X1 port map( A1 => n12718, A2 => n13309, B1 => n12713, B2 => 
                           n11930, ZN => n5548);
   U3967 : OAI22_X1 port map( A1 => n12718, A2 => n13312, B1 => n12713, B2 => 
                           n11931, ZN => n5549);
   U3968 : OAI22_X1 port map( A1 => n12718, A2 => n13315, B1 => n12714, B2 => 
                           n11932, ZN => n5550);
   U3969 : OAI22_X1 port map( A1 => n12717, A2 => n13318, B1 => n12714, B2 => 
                           n11933, ZN => n5551);
   U3970 : OAI22_X1 port map( A1 => n12722, A2 => n13243, B1 => n12712, B2 => 
                           n11934, ZN => n5526);
   U3971 : OAI22_X1 port map( A1 => n12722, A2 => n13246, B1 => n12712, B2 => 
                           n11935, ZN => n5527);
   U3972 : OAI22_X1 port map( A1 => n12717, A2 => n13321, B1 => n12714, B2 => 
                           n11936, ZN => n5552);
   U3973 : OAI22_X1 port map( A1 => n12717, A2 => n13324, B1 => n12714, B2 => 
                           n11937, ZN => n5553);
   U3974 : OAI22_X1 port map( A1 => n12717, A2 => n13327, B1 => n12714, B2 => 
                           n11938, ZN => n5554);
   U3975 : OAI22_X1 port map( A1 => n12717, A2 => n13330, B1 => n12714, B2 => 
                           n11939, ZN => n5555);
   U3976 : OAI22_X1 port map( A1 => n12716, A2 => n13333, B1 => n12714, B2 => 
                           n11940, ZN => n5556);
   U3977 : OAI22_X1 port map( A1 => n12716, A2 => n13336, B1 => n12714, B2 => 
                           n11941, ZN => n5557);
   U3978 : OAI22_X1 port map( A1 => n12716, A2 => n13339, B1 => n12714, B2 => 
                           n11942, ZN => n5558);
   U3979 : OAI22_X1 port map( A1 => n12716, A2 => n13342, B1 => n12714, B2 => 
                           n11943, ZN => n5559);
   U3980 : OAI22_X1 port map( A1 => n12716, A2 => n13345, B1 => n12714, B2 => 
                           n11944, ZN => n5560);
   U3981 : OAI22_X1 port map( A1 => n12715, A2 => n13348, B1 => n12714, B2 => 
                           n11945, ZN => n5561);
   U3982 : OAI22_X1 port map( A1 => n12742, A2 => n13243, B1 => n12732, B2 => 
                           n12057, ZN => n5590);
   U3983 : OAI22_X1 port map( A1 => n12742, A2 => n13246, B1 => n12732, B2 => 
                           n12058, ZN => n5591);
   U3984 : OAI22_X1 port map( A1 => n12742, A2 => n13249, B1 => n12732, B2 => 
                           n12059, ZN => n5592);
   U3985 : OAI22_X1 port map( A1 => n12742, A2 => n13252, B1 => n12732, B2 => 
                           n12060, ZN => n5593);
   U3986 : OAI22_X1 port map( A1 => n12742, A2 => n13255, B1 => n12732, B2 => 
                           n12061, ZN => n5594);
   U3987 : OAI22_X1 port map( A1 => n12741, A2 => n13258, B1 => n12732, B2 => 
                           n12062, ZN => n5595);
   U3988 : OAI22_X1 port map( A1 => n12741, A2 => n13261, B1 => n12732, B2 => 
                           n12063, ZN => n5596);
   U3989 : OAI22_X1 port map( A1 => n12741, A2 => n13264, B1 => n12732, B2 => 
                           n12064, ZN => n5597);
   U3990 : OAI22_X1 port map( A1 => n12741, A2 => n13267, B1 => n12732, B2 => 
                           n12065, ZN => n5598);
   U3991 : OAI22_X1 port map( A1 => n12741, A2 => n13270, B1 => n12732, B2 => 
                           n12066, ZN => n5599);
   U3992 : OAI22_X1 port map( A1 => n12740, A2 => n13273, B1 => n12732, B2 => 
                           n12067, ZN => n5600);
   U3993 : OAI22_X1 port map( A1 => n12740, A2 => n13276, B1 => n12732, B2 => 
                           n12068, ZN => n5601);
   U3994 : OAI22_X1 port map( A1 => n12740, A2 => n13279, B1 => n12733, B2 => 
                           n12069, ZN => n5602);
   U3995 : OAI22_X1 port map( A1 => n12740, A2 => n13282, B1 => n12733, B2 => 
                           n12070, ZN => n5603);
   U3996 : OAI22_X1 port map( A1 => n12740, A2 => n13285, B1 => n12733, B2 => 
                           n12071, ZN => n5604);
   U3997 : OAI22_X1 port map( A1 => n12739, A2 => n13288, B1 => n12733, B2 => 
                           n12072, ZN => n5605);
   U3998 : OAI22_X1 port map( A1 => n12739, A2 => n13291, B1 => n12733, B2 => 
                           n12073, ZN => n5606);
   U3999 : OAI22_X1 port map( A1 => n12739, A2 => n13294, B1 => n12733, B2 => 
                           n12074, ZN => n5607);
   U4000 : OAI22_X1 port map( A1 => n12739, A2 => n13297, B1 => n12733, B2 => 
                           n12075, ZN => n5608);
   U4001 : OAI22_X1 port map( A1 => n12739, A2 => n13300, B1 => n12733, B2 => 
                           n12076, ZN => n5609);
   U4002 : OAI22_X1 port map( A1 => n12738, A2 => n13303, B1 => n12733, B2 => 
                           n12077, ZN => n5610);
   U4003 : OAI22_X1 port map( A1 => n12738, A2 => n13306, B1 => n12733, B2 => 
                           n12078, ZN => n5611);
   U4004 : OAI22_X1 port map( A1 => n12738, A2 => n13309, B1 => n12733, B2 => 
                           n12079, ZN => n5612);
   U4005 : OAI22_X1 port map( A1 => n12738, A2 => n13312, B1 => n12733, B2 => 
                           n12080, ZN => n5613);
   U4006 : OAI22_X1 port map( A1 => n12738, A2 => n13315, B1 => n12734, B2 => 
                           n12081, ZN => n5614);
   U4007 : OAI22_X1 port map( A1 => n12737, A2 => n13318, B1 => n12734, B2 => 
                           n12082, ZN => n5615);
   U4008 : OAI22_X1 port map( A1 => n12737, A2 => n13321, B1 => n12734, B2 => 
                           n12083, ZN => n5616);
   U4009 : OAI22_X1 port map( A1 => n12737, A2 => n13324, B1 => n12734, B2 => 
                           n12084, ZN => n5617);
   U4010 : OAI22_X1 port map( A1 => n12737, A2 => n13327, B1 => n12734, B2 => 
                           n12085, ZN => n5618);
   U4011 : OAI22_X1 port map( A1 => n12737, A2 => n13330, B1 => n12734, B2 => 
                           n12086, ZN => n5619);
   U4012 : OAI22_X1 port map( A1 => n12736, A2 => n13333, B1 => n12734, B2 => 
                           n12087, ZN => n5620);
   U4013 : OAI22_X1 port map( A1 => n12736, A2 => n13336, B1 => n12734, B2 => 
                           n12088, ZN => n5621);
   U4014 : OAI22_X1 port map( A1 => n12736, A2 => n13339, B1 => n12734, B2 => 
                           n12089, ZN => n5622);
   U4015 : OAI22_X1 port map( A1 => n12736, A2 => n13342, B1 => n12734, B2 => 
                           n12090, ZN => n5623);
   U4016 : OAI22_X1 port map( A1 => n12736, A2 => n13345, B1 => n12734, B2 => 
                           n12091, ZN => n5624);
   U4017 : OAI22_X1 port map( A1 => n12735, A2 => n13348, B1 => n12734, B2 => 
                           n12092, ZN => n5625);
   U4018 : OAI22_X1 port map( A1 => n12798, A2 => n13312, B1 => n12793, B2 => 
                           n11946, ZN => n5805);
   U4019 : OAI22_X1 port map( A1 => n12798, A2 => n13315, B1 => n12794, B2 => 
                           n11947, ZN => n5806);
   U4020 : OAI22_X1 port map( A1 => n12797, A2 => n13318, B1 => n12794, B2 => 
                           n11948, ZN => n5807);
   U4021 : OAI22_X1 port map( A1 => n12797, A2 => n13321, B1 => n12794, B2 => 
                           n11949, ZN => n5808);
   U4022 : OAI22_X1 port map( A1 => n12797, A2 => n13324, B1 => n12794, B2 => 
                           n11950, ZN => n5809);
   U4023 : OAI22_X1 port map( A1 => n12797, A2 => n13327, B1 => n12794, B2 => 
                           n11951, ZN => n5810);
   U4024 : OAI22_X1 port map( A1 => n12797, A2 => n13330, B1 => n12794, B2 => 
                           n11952, ZN => n5811);
   U4025 : OAI22_X1 port map( A1 => n12796, A2 => n13333, B1 => n12794, B2 => 
                           n11953, ZN => n5812);
   U4026 : OAI22_X1 port map( A1 => n12796, A2 => n13336, B1 => n12794, B2 => 
                           n11954, ZN => n5813);
   U4027 : OAI22_X1 port map( A1 => n12796, A2 => n13339, B1 => n12794, B2 => 
                           n11955, ZN => n5814);
   U4028 : OAI22_X1 port map( A1 => n12796, A2 => n13342, B1 => n12794, B2 => 
                           n11956, ZN => n5815);
   U4029 : OAI22_X1 port map( A1 => n12796, A2 => n13345, B1 => n12794, B2 => 
                           n11957, ZN => n5816);
   U4030 : OAI22_X1 port map( A1 => n12795, A2 => n13348, B1 => n12794, B2 => 
                           n11958, ZN => n5817);
   U4031 : OAI22_X1 port map( A1 => n12822, A2 => n13243, B1 => n12812, B2 => 
                           n12093, ZN => n5846);
   U4032 : OAI22_X1 port map( A1 => n12822, A2 => n13246, B1 => n12812, B2 => 
                           n12094, ZN => n5847);
   U4033 : OAI22_X1 port map( A1 => n12822, A2 => n13249, B1 => n12812, B2 => 
                           n12095, ZN => n5848);
   U4034 : OAI22_X1 port map( A1 => n12822, A2 => n13252, B1 => n12812, B2 => 
                           n12096, ZN => n5849);
   U4035 : OAI22_X1 port map( A1 => n12822, A2 => n13255, B1 => n12812, B2 => 
                           n12097, ZN => n5850);
   U4036 : OAI22_X1 port map( A1 => n12821, A2 => n13258, B1 => n12812, B2 => 
                           n12098, ZN => n5851);
   U4037 : OAI22_X1 port map( A1 => n12821, A2 => n13261, B1 => n12812, B2 => 
                           n12099, ZN => n5852);
   U4038 : OAI22_X1 port map( A1 => n12821, A2 => n13264, B1 => n12812, B2 => 
                           n12100, ZN => n5853);
   U4039 : OAI22_X1 port map( A1 => n12821, A2 => n13267, B1 => n12812, B2 => 
                           n12101, ZN => n5854);
   U4040 : OAI22_X1 port map( A1 => n12821, A2 => n13270, B1 => n12812, B2 => 
                           n12102, ZN => n5855);
   U4041 : OAI22_X1 port map( A1 => n12820, A2 => n13273, B1 => n12812, B2 => 
                           n12103, ZN => n5856);
   U4042 : OAI22_X1 port map( A1 => n12820, A2 => n13276, B1 => n12812, B2 => 
                           n12104, ZN => n5857);
   U4043 : OAI22_X1 port map( A1 => n12820, A2 => n13279, B1 => n12813, B2 => 
                           n12105, ZN => n5858);
   U4044 : OAI22_X1 port map( A1 => n12820, A2 => n13282, B1 => n12813, B2 => 
                           n12106, ZN => n5859);
   U4045 : OAI22_X1 port map( A1 => n12820, A2 => n13285, B1 => n12813, B2 => 
                           n12107, ZN => n5860);
   U4046 : OAI22_X1 port map( A1 => n12819, A2 => n13288, B1 => n12813, B2 => 
                           n12108, ZN => n5861);
   U4047 : OAI22_X1 port map( A1 => n12819, A2 => n13291, B1 => n12813, B2 => 
                           n12109, ZN => n5862);
   U4048 : OAI22_X1 port map( A1 => n12819, A2 => n13294, B1 => n12813, B2 => 
                           n12110, ZN => n5863);
   U4049 : OAI22_X1 port map( A1 => n12819, A2 => n13297, B1 => n12813, B2 => 
                           n12111, ZN => n5864);
   U4050 : OAI22_X1 port map( A1 => n12819, A2 => n13300, B1 => n12813, B2 => 
                           n12112, ZN => n5865);
   U4051 : OAI22_X1 port map( A1 => n12818, A2 => n13303, B1 => n12813, B2 => 
                           n12113, ZN => n5866);
   U4052 : OAI22_X1 port map( A1 => n12818, A2 => n13306, B1 => n12813, B2 => 
                           n12114, ZN => n5867);
   U4053 : OAI22_X1 port map( A1 => n12818, A2 => n13309, B1 => n12813, B2 => 
                           n12115, ZN => n5868);
   U4054 : OAI22_X1 port map( A1 => n12818, A2 => n13312, B1 => n12813, B2 => 
                           n12116, ZN => n5869);
   U4055 : OAI22_X1 port map( A1 => n12818, A2 => n13315, B1 => n12814, B2 => 
                           n12117, ZN => n5870);
   U4056 : OAI22_X1 port map( A1 => n12817, A2 => n13318, B1 => n12814, B2 => 
                           n12118, ZN => n5871);
   U4057 : OAI22_X1 port map( A1 => n12817, A2 => n13321, B1 => n12814, B2 => 
                           n12119, ZN => n5872);
   U4058 : OAI22_X1 port map( A1 => n12817, A2 => n13324, B1 => n12814, B2 => 
                           n12120, ZN => n5873);
   U4059 : OAI22_X1 port map( A1 => n12817, A2 => n13327, B1 => n12814, B2 => 
                           n12121, ZN => n5874);
   U4060 : OAI22_X1 port map( A1 => n12817, A2 => n13330, B1 => n12814, B2 => 
                           n12122, ZN => n5875);
   U4061 : OAI22_X1 port map( A1 => n12816, A2 => n13333, B1 => n12814, B2 => 
                           n12123, ZN => n5876);
   U4062 : OAI22_X1 port map( A1 => n12816, A2 => n13336, B1 => n12814, B2 => 
                           n12124, ZN => n5877);
   U4063 : OAI22_X1 port map( A1 => n12816, A2 => n13339, B1 => n12814, B2 => 
                           n12125, ZN => n5878);
   U4064 : OAI22_X1 port map( A1 => n12816, A2 => n13342, B1 => n12814, B2 => 
                           n12126, ZN => n5879);
   U4065 : OAI22_X1 port map( A1 => n12816, A2 => n13345, B1 => n12814, B2 => 
                           n12127, ZN => n5880);
   U4066 : OAI22_X1 port map( A1 => n12815, A2 => n13348, B1 => n12814, B2 => 
                           n12128, ZN => n5881);
   U4067 : OAI22_X1 port map( A1 => n8515, A2 => n12551, B1 => n12571, B2 => 
                           n13184, ZN => n4994);
   U4068 : OAI22_X1 port map( A1 => n8498, A2 => n12551, B1 => n12571, B2 => 
                           n13187, ZN => n4995);
   U4069 : OAI22_X1 port map( A1 => n8481, A2 => n12551, B1 => n12571, B2 => 
                           n13190, ZN => n4996);
   U4070 : OAI22_X1 port map( A1 => n8464, A2 => n12551, B1 => n12571, B2 => 
                           n13193, ZN => n4997);
   U4071 : OAI22_X1 port map( A1 => n8447, A2 => n12551, B1 => n12570, B2 => 
                           n13196, ZN => n4998);
   U4072 : OAI22_X1 port map( A1 => n8430, A2 => n12551, B1 => n12570, B2 => 
                           n13199, ZN => n4999);
   U4073 : OAI22_X1 port map( A1 => n8413, A2 => n12551, B1 => n12570, B2 => 
                           n13202, ZN => n5000);
   U4074 : OAI22_X1 port map( A1 => n8396, A2 => n12551, B1 => n12570, B2 => 
                           n13205, ZN => n5001);
   U4075 : OAI22_X1 port map( A1 => n8379, A2 => n12552, B1 => n12569, B2 => 
                           n13208, ZN => n5002);
   U4076 : OAI22_X1 port map( A1 => n8362, A2 => n12552, B1 => n12569, B2 => 
                           n13211, ZN => n5003);
   U4077 : OAI22_X1 port map( A1 => n8345, A2 => n12552, B1 => n12569, B2 => 
                           n13214, ZN => n5004);
   U4078 : OAI22_X1 port map( A1 => n8328, A2 => n12552, B1 => n12569, B2 => 
                           n13217, ZN => n5005);
   U4079 : OAI22_X1 port map( A1 => n8311, A2 => n12552, B1 => n12568, B2 => 
                           n13220, ZN => n5006);
   U4080 : OAI22_X1 port map( A1 => n8294, A2 => n12552, B1 => n12568, B2 => 
                           n13223, ZN => n5007);
   U4081 : OAI22_X1 port map( A1 => n8277, A2 => n12552, B1 => n12568, B2 => 
                           n13226, ZN => n5008);
   U4082 : OAI22_X1 port map( A1 => n8260, A2 => n12552, B1 => n12568, B2 => 
                           n13229, ZN => n5009);
   U4083 : OAI22_X1 port map( A1 => n8243, A2 => n12552, B1 => n12567, B2 => 
                           n13232, ZN => n5010);
   U4084 : OAI22_X1 port map( A1 => n8226, A2 => n12552, B1 => n12567, B2 => 
                           n13235, ZN => n5011);
   U4085 : OAI22_X1 port map( A1 => n8209, A2 => n12552, B1 => n12567, B2 => 
                           n13238, ZN => n5012);
   U4086 : OAI22_X1 port map( A1 => n8192, A2 => n12552, B1 => n12567, B2 => 
                           n13241, ZN => n5013);
   U4087 : OAI22_X1 port map( A1 => n8175, A2 => n12553, B1 => n12566, B2 => 
                           n13244, ZN => n5014);
   U4088 : OAI22_X1 port map( A1 => n8158, A2 => n12553, B1 => n12566, B2 => 
                           n13247, ZN => n5015);
   U4089 : OAI22_X1 port map( A1 => n8141, A2 => n12553, B1 => n12566, B2 => 
                           n13250, ZN => n5016);
   U4090 : OAI22_X1 port map( A1 => n8124, A2 => n12553, B1 => n12566, B2 => 
                           n13253, ZN => n5017);
   U4091 : OAI22_X1 port map( A1 => n8107, A2 => n12553, B1 => n12565, B2 => 
                           n13256, ZN => n5018);
   U4092 : OAI22_X1 port map( A1 => n8090, A2 => n12553, B1 => n12565, B2 => 
                           n13259, ZN => n5019);
   U4093 : OAI22_X1 port map( A1 => n8073, A2 => n12553, B1 => n12565, B2 => 
                           n13262, ZN => n5020);
   U4094 : OAI22_X1 port map( A1 => n8056, A2 => n12553, B1 => n12565, B2 => 
                           n13265, ZN => n5021);
   U4095 : OAI22_X1 port map( A1 => n8039, A2 => n12553, B1 => n12564, B2 => 
                           n13268, ZN => n5022);
   U4096 : OAI22_X1 port map( A1 => n8022, A2 => n12553, B1 => n12564, B2 => 
                           n13271, ZN => n5023);
   U4097 : OAI22_X1 port map( A1 => n8005, A2 => n12553, B1 => n12564, B2 => 
                           n13274, ZN => n5024);
   U4098 : OAI22_X1 port map( A1 => n7988, A2 => n12553, B1 => n12564, B2 => 
                           n13277, ZN => n5025);
   U4099 : OAI22_X1 port map( A1 => n7971, A2 => n12554, B1 => n12563, B2 => 
                           n13280, ZN => n5026);
   U4100 : OAI22_X1 port map( A1 => n7954, A2 => n12554, B1 => n12563, B2 => 
                           n13283, ZN => n5027);
   U4101 : OAI22_X1 port map( A1 => n7937, A2 => n12554, B1 => n12563, B2 => 
                           n13286, ZN => n5028);
   U4102 : OAI22_X1 port map( A1 => n7920, A2 => n12554, B1 => n12563, B2 => 
                           n13289, ZN => n5029);
   U4103 : OAI22_X1 port map( A1 => n7903, A2 => n12554, B1 => n12562, B2 => 
                           n13292, ZN => n5030);
   U4104 : OAI22_X1 port map( A1 => n7886, A2 => n12554, B1 => n12562, B2 => 
                           n13295, ZN => n5031);
   U4105 : OAI22_X1 port map( A1 => n7869, A2 => n12554, B1 => n12562, B2 => 
                           n13298, ZN => n5032);
   U4106 : OAI22_X1 port map( A1 => n7852, A2 => n12554, B1 => n12562, B2 => 
                           n13301, ZN => n5033);
   U4107 : OAI22_X1 port map( A1 => n7835, A2 => n12554, B1 => n12561, B2 => 
                           n13304, ZN => n5034);
   U4108 : OAI22_X1 port map( A1 => n7818, A2 => n12554, B1 => n12561, B2 => 
                           n13307, ZN => n5035);
   U4109 : OAI22_X1 port map( A1 => n7801, A2 => n12554, B1 => n12561, B2 => 
                           n13310, ZN => n5036);
   U4110 : OAI22_X1 port map( A1 => n7784, A2 => n12554, B1 => n12561, B2 => 
                           n13313, ZN => n5037);
   U4111 : OAI22_X1 port map( A1 => n7767, A2 => n12555, B1 => n12560, B2 => 
                           n13316, ZN => n5038);
   U4112 : OAI22_X1 port map( A1 => n7750, A2 => n12555, B1 => n12560, B2 => 
                           n13319, ZN => n5039);
   U4113 : OAI22_X1 port map( A1 => n7648, A2 => n12555, B1 => n12560, B2 => 
                           n13322, ZN => n5040);
   U4114 : OAI22_X1 port map( A1 => n7631, A2 => n12555, B1 => n12560, B2 => 
                           n13325, ZN => n5041);
   U4115 : OAI22_X1 port map( A1 => n7527, A2 => n12555, B1 => n12559, B2 => 
                           n13328, ZN => n5042);
   U4116 : OAI22_X1 port map( A1 => n7510, A2 => n12555, B1 => n12559, B2 => 
                           n13331, ZN => n5043);
   U4117 : OAI22_X1 port map( A1 => n7493, A2 => n12555, B1 => n12559, B2 => 
                           n13334, ZN => n5044);
   U4118 : OAI22_X1 port map( A1 => n7391, A2 => n12555, B1 => n12559, B2 => 
                           n13337, ZN => n5045);
   U4119 : OAI22_X1 port map( A1 => n7374, A2 => n12555, B1 => n12558, B2 => 
                           n13340, ZN => n5046);
   U4120 : OAI22_X1 port map( A1 => n7275, A2 => n12555, B1 => n12558, B2 => 
                           n13343, ZN => n5047);
   U4121 : OAI22_X1 port map( A1 => n7258, A2 => n12555, B1 => n12558, B2 => 
                           n13346, ZN => n5048);
   U4122 : OAI22_X1 port map( A1 => n7241, A2 => n12555, B1 => n12558, B2 => 
                           n13349, ZN => n5049);
   U4123 : OAI22_X1 port map( A1 => n7144, A2 => n12556, B1 => n12557, B2 => 
                           n13352, ZN => n5050);
   U4124 : OAI22_X1 port map( A1 => n7127, A2 => n12556, B1 => n12557, B2 => 
                           n13355, ZN => n5051);
   U4125 : OAI22_X1 port map( A1 => n7110, A2 => n12556, B1 => n12557, B2 => 
                           n13358, ZN => n5052);
   U4126 : OAI22_X1 port map( A1 => n4849, A2 => n12556, B1 => n12557, B2 => 
                           n13381, ZN => n5053);
   U4127 : OAI22_X1 port map( A1 => n8583, A2 => n12551, B1 => n12572, B2 => 
                           n13172, ZN => n4990);
   U4128 : OAI22_X1 port map( A1 => n8566, A2 => n12551, B1 => n12572, B2 => 
                           n13175, ZN => n4991);
   U4129 : OAI22_X1 port map( A1 => n8549, A2 => n12551, B1 => n12572, B2 => 
                           n13178, ZN => n4992);
   U4130 : OAI22_X1 port map( A1 => n8532, A2 => n12551, B1 => n12572, B2 => 
                           n13181, ZN => n4993);
   U4131 : OAI22_X1 port map( A1 => n12927, A2 => n13171, B1 => n8575, B2 => 
                           n12911, ZN => n6142);
   U4132 : OAI22_X1 port map( A1 => n12927, A2 => n13174, B1 => n8558, B2 => 
                           n12911, ZN => n6143);
   U4133 : OAI22_X1 port map( A1 => n12927, A2 => n13177, B1 => n8541, B2 => 
                           n12911, ZN => n6144);
   U4134 : OAI22_X1 port map( A1 => n12927, A2 => n13180, B1 => n8524, B2 => 
                           n12911, ZN => n6145);
   U4135 : OAI22_X1 port map( A1 => n12926, A2 => n13183, B1 => n8507, B2 => 
                           n12911, ZN => n6146);
   U4136 : OAI22_X1 port map( A1 => n12926, A2 => n13186, B1 => n8490, B2 => 
                           n12911, ZN => n6147);
   U4137 : OAI22_X1 port map( A1 => n12926, A2 => n13189, B1 => n8473, B2 => 
                           n12911, ZN => n6148);
   U4138 : OAI22_X1 port map( A1 => n12926, A2 => n13192, B1 => n8456, B2 => 
                           n12911, ZN => n6149);
   U4139 : OAI22_X1 port map( A1 => n12926, A2 => n13195, B1 => n8439, B2 => 
                           n12911, ZN => n6150);
   U4140 : OAI22_X1 port map( A1 => n12925, A2 => n13198, B1 => n8422, B2 => 
                           n12911, ZN => n6151);
   U4141 : OAI22_X1 port map( A1 => n12925, A2 => n13201, B1 => n8405, B2 => 
                           n12911, ZN => n6152);
   U4142 : OAI22_X1 port map( A1 => n12925, A2 => n13204, B1 => n8388, B2 => 
                           n12911, ZN => n6153);
   U4143 : OAI22_X1 port map( A1 => n12925, A2 => n13207, B1 => n8371, B2 => 
                           n12913, ZN => n6154);
   U4144 : OAI22_X1 port map( A1 => n12925, A2 => n13210, B1 => n8354, B2 => 
                           n12914, ZN => n6155);
   U4145 : OAI22_X1 port map( A1 => n12924, A2 => n13213, B1 => n8337, B2 => 
                           n12911, ZN => n6156);
   U4146 : OAI22_X1 port map( A1 => n12924, A2 => n13216, B1 => n8320, B2 => 
                           n12913, ZN => n6157);
   U4147 : OAI22_X1 port map( A1 => n12924, A2 => n13219, B1 => n8303, B2 => 
                           n12914, ZN => n6158);
   U4148 : OAI22_X1 port map( A1 => n12924, A2 => n13222, B1 => n8286, B2 => 
                           n12910, ZN => n6159);
   U4149 : OAI22_X1 port map( A1 => n12924, A2 => n13225, B1 => n8269, B2 => 
                           n1929, ZN => n6160);
   U4150 : OAI22_X1 port map( A1 => n12923, A2 => n13228, B1 => n8252, B2 => 
                           n1929, ZN => n6161);
   U4151 : OAI22_X1 port map( A1 => n12923, A2 => n13231, B1 => n8235, B2 => 
                           n1929, ZN => n6162);
   U4152 : OAI22_X1 port map( A1 => n12923, A2 => n13234, B1 => n8218, B2 => 
                           n1929, ZN => n6163);
   U4153 : OAI22_X1 port map( A1 => n12923, A2 => n13237, B1 => n8201, B2 => 
                           n1929, ZN => n6164);
   U4154 : OAI22_X1 port map( A1 => n12923, A2 => n13240, B1 => n8184, B2 => 
                           n1929, ZN => n6165);
   U4155 : OAI22_X1 port map( A1 => n12593, A2 => n13172, B1 => n8584, B2 => 
                           n12578, ZN => n5054);
   U4156 : OAI22_X1 port map( A1 => n12593, A2 => n13175, B1 => n8567, B2 => 
                           n12577, ZN => n5055);
   U4157 : OAI22_X1 port map( A1 => n12593, A2 => n13178, B1 => n8550, B2 => 
                           n12577, ZN => n5056);
   U4158 : OAI22_X1 port map( A1 => n12592, A2 => n13184, B1 => n8516, B2 => 
                           n1948, ZN => n5058);
   U4159 : OAI22_X1 port map( A1 => n12593, A2 => n13181, B1 => n8533, B2 => 
                           n1948, ZN => n5057);
   U4160 : OAI22_X1 port map( A1 => n12592, A2 => n13187, B1 => n8499, B2 => 
                           n1948, ZN => n5059);
   U4161 : OAI22_X1 port map( A1 => n12592, A2 => n13190, B1 => n8482, B2 => 
                           n1948, ZN => n5060);
   U4162 : OAI22_X1 port map( A1 => n12592, A2 => n13193, B1 => n8465, B2 => 
                           n1948, ZN => n5061);
   U4163 : OAI22_X1 port map( A1 => n12592, A2 => n13196, B1 => n8448, B2 => 
                           n12577, ZN => n5062);
   U4164 : OAI22_X1 port map( A1 => n12591, A2 => n13199, B1 => n8431, B2 => 
                           n12577, ZN => n5063);
   U4165 : OAI22_X1 port map( A1 => n12591, A2 => n13202, B1 => n8414, B2 => 
                           n12577, ZN => n5064);
   U4166 : OAI22_X1 port map( A1 => n12591, A2 => n13205, B1 => n8397, B2 => 
                           n12577, ZN => n5065);
   U4167 : OAI22_X1 port map( A1 => n12591, A2 => n13208, B1 => n8380, B2 => 
                           n12579, ZN => n5066);
   U4168 : OAI22_X1 port map( A1 => n12591, A2 => n13211, B1 => n8363, B2 => 
                           n12580, ZN => n5067);
   U4169 : OAI22_X1 port map( A1 => n12590, A2 => n13214, B1 => n8346, B2 => 
                           n12578, ZN => n5068);
   U4170 : OAI22_X1 port map( A1 => n12590, A2 => n13217, B1 => n8329, B2 => 
                           n12579, ZN => n5069);
   U4171 : OAI22_X1 port map( A1 => n12590, A2 => n13220, B1 => n8312, B2 => 
                           n12580, ZN => n5070);
   U4172 : OAI22_X1 port map( A1 => n12590, A2 => n13223, B1 => n8295, B2 => 
                           n12577, ZN => n5071);
   U4173 : OAI22_X1 port map( A1 => n12590, A2 => n13226, B1 => n8278, B2 => 
                           n1948, ZN => n5072);
   U4174 : OAI22_X1 port map( A1 => n12589, A2 => n13229, B1 => n8261, B2 => 
                           n1948, ZN => n5073);
   U4175 : OAI22_X1 port map( A1 => n12589, A2 => n13232, B1 => n8244, B2 => 
                           n1948, ZN => n5074);
   U4176 : OAI22_X1 port map( A1 => n12589, A2 => n13235, B1 => n8227, B2 => 
                           n1948, ZN => n5075);
   U4177 : OAI22_X1 port map( A1 => n12589, A2 => n13238, B1 => n8210, B2 => 
                           n1948, ZN => n5076);
   U4178 : OAI22_X1 port map( A1 => n12589, A2 => n13241, B1 => n8193, B2 => 
                           n1948, ZN => n5077);
   U4179 : OAI22_X1 port map( A1 => n13007, A2 => n13170, B1 => n8573, B2 => 
                           n12991, ZN => n6398);
   U4180 : OAI22_X1 port map( A1 => n13007, A2 => n13173, B1 => n8556, B2 => 
                           n12991, ZN => n6399);
   U4181 : OAI22_X1 port map( A1 => n13007, A2 => n13176, B1 => n8539, B2 => 
                           n12991, ZN => n6400);
   U4182 : OAI22_X1 port map( A1 => n13007, A2 => n13179, B1 => n8522, B2 => 
                           n12991, ZN => n6401);
   U4183 : OAI22_X1 port map( A1 => n13006, A2 => n13182, B1 => n8505, B2 => 
                           n12991, ZN => n6402);
   U4184 : OAI22_X1 port map( A1 => n13006, A2 => n13185, B1 => n8488, B2 => 
                           n12991, ZN => n6403);
   U4185 : OAI22_X1 port map( A1 => n13006, A2 => n13188, B1 => n8471, B2 => 
                           n12991, ZN => n6404);
   U4186 : OAI22_X1 port map( A1 => n13006, A2 => n13191, B1 => n8454, B2 => 
                           n12991, ZN => n6405);
   U4187 : OAI22_X1 port map( A1 => n13006, A2 => n13194, B1 => n8437, B2 => 
                           n12991, ZN => n6406);
   U4188 : OAI22_X1 port map( A1 => n13005, A2 => n13197, B1 => n8420, B2 => 
                           n12991, ZN => n6407);
   U4189 : OAI22_X1 port map( A1 => n13005, A2 => n13200, B1 => n8403, B2 => 
                           n12991, ZN => n6408);
   U4190 : OAI22_X1 port map( A1 => n13005, A2 => n13203, B1 => n8386, B2 => 
                           n12991, ZN => n6409);
   U4191 : OAI22_X1 port map( A1 => n13005, A2 => n13206, B1 => n8369, B2 => 
                           n12993, ZN => n6410);
   U4192 : OAI22_X1 port map( A1 => n13005, A2 => n13209, B1 => n8352, B2 => 
                           n12994, ZN => n6411);
   U4193 : OAI22_X1 port map( A1 => n13004, A2 => n13212, B1 => n8335, B2 => 
                           n12991, ZN => n6412);
   U4194 : OAI22_X1 port map( A1 => n13004, A2 => n13215, B1 => n8318, B2 => 
                           n12993, ZN => n6413);
   U4195 : OAI22_X1 port map( A1 => n13004, A2 => n13218, B1 => n8301, B2 => 
                           n12994, ZN => n6414);
   U4196 : OAI22_X1 port map( A1 => n13004, A2 => n13221, B1 => n8284, B2 => 
                           n12990, ZN => n6415);
   U4197 : OAI22_X1 port map( A1 => n13004, A2 => n13224, B1 => n8267, B2 => 
                           n1925, ZN => n6416);
   U4198 : OAI22_X1 port map( A1 => n13003, A2 => n13227, B1 => n8250, B2 => 
                           n1925, ZN => n6417);
   U4199 : OAI22_X1 port map( A1 => n13003, A2 => n13230, B1 => n8233, B2 => 
                           n1925, ZN => n6418);
   U4200 : OAI22_X1 port map( A1 => n13003, A2 => n13233, B1 => n8216, B2 => 
                           n1925, ZN => n6419);
   U4201 : OAI22_X1 port map( A1 => n13003, A2 => n13236, B1 => n8199, B2 => 
                           n1925, ZN => n6420);
   U4202 : OAI22_X1 port map( A1 => n13003, A2 => n13239, B1 => n8182, B2 => 
                           n1925, ZN => n6421);
   U4203 : OAI22_X1 port map( A1 => n12847, A2 => n13171, B1 => n8577, B2 => 
                           n12831, ZN => n5886);
   U4204 : OAI22_X1 port map( A1 => n12847, A2 => n13174, B1 => n8560, B2 => 
                           n12831, ZN => n5887);
   U4205 : OAI22_X1 port map( A1 => n12847, A2 => n13177, B1 => n8543, B2 => 
                           n12831, ZN => n5888);
   U4206 : OAI22_X1 port map( A1 => n12847, A2 => n13180, B1 => n8526, B2 => 
                           n12831, ZN => n5889);
   U4207 : OAI22_X1 port map( A1 => n12846, A2 => n13183, B1 => n8509, B2 => 
                           n12831, ZN => n5890);
   U4208 : OAI22_X1 port map( A1 => n12846, A2 => n13186, B1 => n8492, B2 => 
                           n12831, ZN => n5891);
   U4209 : OAI22_X1 port map( A1 => n12846, A2 => n13189, B1 => n8475, B2 => 
                           n12831, ZN => n5892);
   U4210 : OAI22_X1 port map( A1 => n12846, A2 => n13192, B1 => n8458, B2 => 
                           n12831, ZN => n5893);
   U4211 : OAI22_X1 port map( A1 => n12846, A2 => n13195, B1 => n8441, B2 => 
                           n12831, ZN => n5894);
   U4212 : OAI22_X1 port map( A1 => n12845, A2 => n13198, B1 => n8424, B2 => 
                           n12831, ZN => n5895);
   U4213 : OAI22_X1 port map( A1 => n12845, A2 => n13201, B1 => n8407, B2 => 
                           n12831, ZN => n5896);
   U4214 : OAI22_X1 port map( A1 => n12845, A2 => n13204, B1 => n8390, B2 => 
                           n12831, ZN => n5897);
   U4215 : OAI22_X1 port map( A1 => n12845, A2 => n13207, B1 => n8373, B2 => 
                           n12833, ZN => n5898);
   U4216 : OAI22_X1 port map( A1 => n12845, A2 => n13210, B1 => n8356, B2 => 
                           n12834, ZN => n5899);
   U4217 : OAI22_X1 port map( A1 => n12844, A2 => n13213, B1 => n8339, B2 => 
                           n12831, ZN => n5900);
   U4218 : OAI22_X1 port map( A1 => n12844, A2 => n13216, B1 => n8322, B2 => 
                           n12833, ZN => n5901);
   U4219 : OAI22_X1 port map( A1 => n12844, A2 => n13219, B1 => n8305, B2 => 
                           n12834, ZN => n5902);
   U4220 : OAI22_X1 port map( A1 => n12844, A2 => n13222, B1 => n8288, B2 => 
                           n12830, ZN => n5903);
   U4221 : OAI22_X1 port map( A1 => n12844, A2 => n13225, B1 => n8271, B2 => 
                           n1934, ZN => n5904);
   U4222 : OAI22_X1 port map( A1 => n12843, A2 => n13228, B1 => n8254, B2 => 
                           n1934, ZN => n5905);
   U4223 : OAI22_X1 port map( A1 => n12843, A2 => n13231, B1 => n8237, B2 => 
                           n1934, ZN => n5906);
   U4224 : OAI22_X1 port map( A1 => n12843, A2 => n13234, B1 => n8220, B2 => 
                           n1934, ZN => n5907);
   U4225 : OAI22_X1 port map( A1 => n12843, A2 => n13237, B1 => n8203, B2 => 
                           n1934, ZN => n5908);
   U4226 : OAI22_X1 port map( A1 => n12843, A2 => n13240, B1 => n8186, B2 => 
                           n1934, ZN => n5909);
   U4227 : OAI22_X1 port map( A1 => n12787, A2 => n13171, B1 => n8580, B2 => 
                           n12771, ZN => n5694);
   U4228 : OAI22_X1 port map( A1 => n12787, A2 => n13174, B1 => n8563, B2 => 
                           n12771, ZN => n5695);
   U4229 : OAI22_X1 port map( A1 => n12787, A2 => n13177, B1 => n8546, B2 => 
                           n12771, ZN => n5696);
   U4230 : OAI22_X1 port map( A1 => n12787, A2 => n13180, B1 => n8529, B2 => 
                           n12771, ZN => n5697);
   U4231 : OAI22_X1 port map( A1 => n12786, A2 => n13183, B1 => n8512, B2 => 
                           n12771, ZN => n5698);
   U4232 : OAI22_X1 port map( A1 => n12786, A2 => n13186, B1 => n8495, B2 => 
                           n12771, ZN => n5699);
   U4233 : OAI22_X1 port map( A1 => n12786, A2 => n13189, B1 => n8478, B2 => 
                           n12771, ZN => n5700);
   U4234 : OAI22_X1 port map( A1 => n12786, A2 => n13192, B1 => n8461, B2 => 
                           n12771, ZN => n5701);
   U4235 : OAI22_X1 port map( A1 => n12786, A2 => n13195, B1 => n8444, B2 => 
                           n12771, ZN => n5702);
   U4236 : OAI22_X1 port map( A1 => n12785, A2 => n13198, B1 => n8427, B2 => 
                           n12771, ZN => n5703);
   U4237 : OAI22_X1 port map( A1 => n12785, A2 => n13201, B1 => n8410, B2 => 
                           n12771, ZN => n5704);
   U4238 : OAI22_X1 port map( A1 => n12785, A2 => n13204, B1 => n8393, B2 => 
                           n12771, ZN => n5705);
   U4239 : OAI22_X1 port map( A1 => n12785, A2 => n13207, B1 => n8376, B2 => 
                           n12773, ZN => n5706);
   U4240 : OAI22_X1 port map( A1 => n12785, A2 => n13210, B1 => n8359, B2 => 
                           n12774, ZN => n5707);
   U4241 : OAI22_X1 port map( A1 => n12784, A2 => n13213, B1 => n8342, B2 => 
                           n12771, ZN => n5708);
   U4242 : OAI22_X1 port map( A1 => n12784, A2 => n13216, B1 => n8325, B2 => 
                           n12773, ZN => n5709);
   U4243 : OAI22_X1 port map( A1 => n12784, A2 => n13219, B1 => n8308, B2 => 
                           n12774, ZN => n5710);
   U4244 : OAI22_X1 port map( A1 => n12784, A2 => n13222, B1 => n8291, B2 => 
                           n12770, ZN => n5711);
   U4245 : OAI22_X1 port map( A1 => n12784, A2 => n13225, B1 => n8274, B2 => 
                           n1937, ZN => n5712);
   U4246 : OAI22_X1 port map( A1 => n12783, A2 => n13228, B1 => n8257, B2 => 
                           n1937, ZN => n5713);
   U4247 : OAI22_X1 port map( A1 => n12783, A2 => n13231, B1 => n8240, B2 => 
                           n1937, ZN => n5714);
   U4248 : OAI22_X1 port map( A1 => n12783, A2 => n13234, B1 => n8223, B2 => 
                           n1937, ZN => n5715);
   U4249 : OAI22_X1 port map( A1 => n12783, A2 => n13237, B1 => n8206, B2 => 
                           n1937, ZN => n5716);
   U4250 : OAI22_X1 port map( A1 => n12783, A2 => n13240, B1 => n8189, B2 => 
                           n1937, ZN => n5717);
   U4251 : OAI22_X1 port map( A1 => n12767, A2 => n13171, B1 => n8579, B2 => 
                           n12751, ZN => n5630);
   U4252 : OAI22_X1 port map( A1 => n12767, A2 => n13174, B1 => n8562, B2 => 
                           n12751, ZN => n5631);
   U4253 : OAI22_X1 port map( A1 => n12767, A2 => n13177, B1 => n8545, B2 => 
                           n12751, ZN => n5632);
   U4254 : OAI22_X1 port map( A1 => n12767, A2 => n13180, B1 => n8528, B2 => 
                           n12751, ZN => n5633);
   U4255 : OAI22_X1 port map( A1 => n12766, A2 => n13183, B1 => n8511, B2 => 
                           n12751, ZN => n5634);
   U4256 : OAI22_X1 port map( A1 => n12766, A2 => n13186, B1 => n8494, B2 => 
                           n12751, ZN => n5635);
   U4257 : OAI22_X1 port map( A1 => n12766, A2 => n13189, B1 => n8477, B2 => 
                           n12751, ZN => n5636);
   U4258 : OAI22_X1 port map( A1 => n12766, A2 => n13192, B1 => n8460, B2 => 
                           n12751, ZN => n5637);
   U4259 : OAI22_X1 port map( A1 => n12766, A2 => n13195, B1 => n8443, B2 => 
                           n12751, ZN => n5638);
   U4260 : OAI22_X1 port map( A1 => n12765, A2 => n13198, B1 => n8426, B2 => 
                           n12751, ZN => n5639);
   U4261 : OAI22_X1 port map( A1 => n12765, A2 => n13201, B1 => n8409, B2 => 
                           n12751, ZN => n5640);
   U4262 : OAI22_X1 port map( A1 => n12765, A2 => n13204, B1 => n8392, B2 => 
                           n12751, ZN => n5641);
   U4263 : OAI22_X1 port map( A1 => n12765, A2 => n13207, B1 => n8375, B2 => 
                           n12753, ZN => n5642);
   U4264 : OAI22_X1 port map( A1 => n12765, A2 => n13210, B1 => n8358, B2 => 
                           n12754, ZN => n5643);
   U4265 : OAI22_X1 port map( A1 => n12764, A2 => n13213, B1 => n8341, B2 => 
                           n12751, ZN => n5644);
   U4266 : OAI22_X1 port map( A1 => n12764, A2 => n13216, B1 => n8324, B2 => 
                           n12753, ZN => n5645);
   U4267 : OAI22_X1 port map( A1 => n12764, A2 => n13219, B1 => n8307, B2 => 
                           n12754, ZN => n5646);
   U4268 : OAI22_X1 port map( A1 => n12764, A2 => n13222, B1 => n8290, B2 => 
                           n12750, ZN => n5647);
   U4269 : OAI22_X1 port map( A1 => n12764, A2 => n13225, B1 => n8273, B2 => 
                           n1938, ZN => n5648);
   U4270 : OAI22_X1 port map( A1 => n12763, A2 => n13228, B1 => n8256, B2 => 
                           n1938, ZN => n5649);
   U4271 : OAI22_X1 port map( A1 => n12763, A2 => n13231, B1 => n8239, B2 => 
                           n1938, ZN => n5650);
   U4272 : OAI22_X1 port map( A1 => n12763, A2 => n13234, B1 => n8222, B2 => 
                           n1938, ZN => n5651);
   U4273 : OAI22_X1 port map( A1 => n12763, A2 => n13237, B1 => n8205, B2 => 
                           n1938, ZN => n5652);
   U4274 : OAI22_X1 port map( A1 => n12763, A2 => n13240, B1 => n8188, B2 => 
                           n1938, ZN => n5653);
   U4275 : OAI22_X1 port map( A1 => n12650, A2 => n13172, B1 => n8581, B2 => 
                           n12635, ZN => n5246);
   U4276 : OAI22_X1 port map( A1 => n12669, A2 => n13172, B1 => n8582, B2 => 
                           n12654, ZN => n5310);
   U4277 : OAI22_X1 port map( A1 => n12650, A2 => n13175, B1 => n8564, B2 => 
                           n12634, ZN => n5247);
   U4278 : OAI22_X1 port map( A1 => n12650, A2 => n13178, B1 => n8547, B2 => 
                           n12634, ZN => n5248);
   U4279 : OAI22_X1 port map( A1 => n12649, A2 => n13184, B1 => n8513, B2 => 
                           n1945, ZN => n5250);
   U4280 : OAI22_X1 port map( A1 => n12650, A2 => n13181, B1 => n8530, B2 => 
                           n1945, ZN => n5249);
   U4281 : OAI22_X1 port map( A1 => n12649, A2 => n13187, B1 => n8496, B2 => 
                           n1945, ZN => n5251);
   U4282 : OAI22_X1 port map( A1 => n12649, A2 => n13190, B1 => n8479, B2 => 
                           n1945, ZN => n5252);
   U4283 : OAI22_X1 port map( A1 => n12649, A2 => n13193, B1 => n8462, B2 => 
                           n1945, ZN => n5253);
   U4284 : OAI22_X1 port map( A1 => n12649, A2 => n13196, B1 => n8445, B2 => 
                           n12634, ZN => n5254);
   U4285 : OAI22_X1 port map( A1 => n12648, A2 => n13199, B1 => n8428, B2 => 
                           n12634, ZN => n5255);
   U4286 : OAI22_X1 port map( A1 => n12648, A2 => n13202, B1 => n8411, B2 => 
                           n12634, ZN => n5256);
   U4287 : OAI22_X1 port map( A1 => n12648, A2 => n13205, B1 => n8394, B2 => 
                           n12634, ZN => n5257);
   U4288 : OAI22_X1 port map( A1 => n12648, A2 => n13208, B1 => n8377, B2 => 
                           n12636, ZN => n5258);
   U4289 : OAI22_X1 port map( A1 => n12648, A2 => n13211, B1 => n8360, B2 => 
                           n12637, ZN => n5259);
   U4290 : OAI22_X1 port map( A1 => n12647, A2 => n13214, B1 => n8343, B2 => 
                           n12635, ZN => n5260);
   U4291 : OAI22_X1 port map( A1 => n12647, A2 => n13217, B1 => n8326, B2 => 
                           n12636, ZN => n5261);
   U4292 : OAI22_X1 port map( A1 => n12647, A2 => n13220, B1 => n8309, B2 => 
                           n12637, ZN => n5262);
   U4293 : OAI22_X1 port map( A1 => n12647, A2 => n13223, B1 => n8292, B2 => 
                           n12634, ZN => n5263);
   U4294 : OAI22_X1 port map( A1 => n12647, A2 => n13226, B1 => n8275, B2 => 
                           n1945, ZN => n5264);
   U4295 : OAI22_X1 port map( A1 => n12646, A2 => n13229, B1 => n8258, B2 => 
                           n1945, ZN => n5265);
   U4296 : OAI22_X1 port map( A1 => n12646, A2 => n13232, B1 => n8241, B2 => 
                           n1945, ZN => n5266);
   U4297 : OAI22_X1 port map( A1 => n12646, A2 => n13235, B1 => n8224, B2 => 
                           n1945, ZN => n5267);
   U4298 : OAI22_X1 port map( A1 => n12646, A2 => n13238, B1 => n8207, B2 => 
                           n1945, ZN => n5268);
   U4299 : OAI22_X1 port map( A1 => n12646, A2 => n13241, B1 => n8190, B2 => 
                           n1945, ZN => n5269);
   U4300 : OAI22_X1 port map( A1 => n12669, A2 => n13175, B1 => n8565, B2 => 
                           n12653, ZN => n5311);
   U4301 : OAI22_X1 port map( A1 => n12669, A2 => n13178, B1 => n8548, B2 => 
                           n12653, ZN => n5312);
   U4302 : OAI22_X1 port map( A1 => n12668, A2 => n13184, B1 => n8514, B2 => 
                           n1944, ZN => n5314);
   U4303 : OAI22_X1 port map( A1 => n12669, A2 => n13181, B1 => n8531, B2 => 
                           n1944, ZN => n5313);
   U4304 : OAI22_X1 port map( A1 => n12668, A2 => n13187, B1 => n8497, B2 => 
                           n1944, ZN => n5315);
   U4305 : OAI22_X1 port map( A1 => n12668, A2 => n13190, B1 => n8480, B2 => 
                           n1944, ZN => n5316);
   U4306 : OAI22_X1 port map( A1 => n12668, A2 => n13193, B1 => n8463, B2 => 
                           n1944, ZN => n5317);
   U4307 : OAI22_X1 port map( A1 => n12668, A2 => n13196, B1 => n8446, B2 => 
                           n12653, ZN => n5318);
   U4308 : OAI22_X1 port map( A1 => n12667, A2 => n13199, B1 => n8429, B2 => 
                           n12653, ZN => n5319);
   U4309 : OAI22_X1 port map( A1 => n12667, A2 => n13202, B1 => n8412, B2 => 
                           n12653, ZN => n5320);
   U4310 : OAI22_X1 port map( A1 => n12667, A2 => n13205, B1 => n8395, B2 => 
                           n12653, ZN => n5321);
   U4311 : OAI22_X1 port map( A1 => n12667, A2 => n13208, B1 => n8378, B2 => 
                           n12655, ZN => n5322);
   U4312 : OAI22_X1 port map( A1 => n12667, A2 => n13211, B1 => n8361, B2 => 
                           n12656, ZN => n5323);
   U4313 : OAI22_X1 port map( A1 => n12666, A2 => n13214, B1 => n8344, B2 => 
                           n12654, ZN => n5324);
   U4314 : OAI22_X1 port map( A1 => n12666, A2 => n13217, B1 => n8327, B2 => 
                           n12655, ZN => n5325);
   U4315 : OAI22_X1 port map( A1 => n12666, A2 => n13220, B1 => n8310, B2 => 
                           n12656, ZN => n5326);
   U4316 : OAI22_X1 port map( A1 => n12666, A2 => n13223, B1 => n8293, B2 => 
                           n12653, ZN => n5327);
   U4317 : OAI22_X1 port map( A1 => n12666, A2 => n13226, B1 => n8276, B2 => 
                           n1944, ZN => n5328);
   U4318 : OAI22_X1 port map( A1 => n12665, A2 => n13229, B1 => n8259, B2 => 
                           n1944, ZN => n5329);
   U4319 : OAI22_X1 port map( A1 => n12665, A2 => n13232, B1 => n8242, B2 => 
                           n1944, ZN => n5330);
   U4320 : OAI22_X1 port map( A1 => n12665, A2 => n13235, B1 => n8225, B2 => 
                           n1944, ZN => n5331);
   U4321 : OAI22_X1 port map( A1 => n12665, A2 => n13238, B1 => n8208, B2 => 
                           n1944, ZN => n5332);
   U4322 : OAI22_X1 port map( A1 => n12665, A2 => n13241, B1 => n8191, B2 => 
                           n1944, ZN => n5333);
   U4323 : OAI22_X1 port map( A1 => n13025, A2 => n13206, B1 => n8370, B2 => 
                           n13011, ZN => n6474);
   U4324 : OAI22_X1 port map( A1 => n13025, A2 => n13209, B1 => n8353, B2 => 
                           n13011, ZN => n6475);
   U4325 : OAI22_X1 port map( A1 => n13024, A2 => n13212, B1 => n8336, B2 => 
                           n13011, ZN => n6476);
   U4326 : OAI22_X1 port map( A1 => n13024, A2 => n13215, B1 => n8319, B2 => 
                           n13011, ZN => n6477);
   U4327 : OAI22_X1 port map( A1 => n13024, A2 => n13218, B1 => n8302, B2 => 
                           n13011, ZN => n6478);
   U4328 : OAI22_X1 port map( A1 => n13024, A2 => n13221, B1 => n8285, B2 => 
                           n13011, ZN => n6479);
   U4329 : OAI22_X1 port map( A1 => n13024, A2 => n13224, B1 => n8268, B2 => 
                           n13011, ZN => n6480);
   U4330 : OAI22_X1 port map( A1 => n13023, A2 => n13227, B1 => n8251, B2 => 
                           n13011, ZN => n6481);
   U4331 : OAI22_X1 port map( A1 => n13023, A2 => n13230, B1 => n8234, B2 => 
                           n13011, ZN => n6482);
   U4332 : OAI22_X1 port map( A1 => n13023, A2 => n13233, B1 => n8217, B2 => 
                           n13011, ZN => n6483);
   U4333 : OAI22_X1 port map( A1 => n13023, A2 => n13236, B1 => n8200, B2 => 
                           n13011, ZN => n6484);
   U4334 : OAI22_X1 port map( A1 => n13023, A2 => n13239, B1 => n8183, B2 => 
                           n13011, ZN => n6485);
   U4335 : OAI22_X1 port map( A1 => n13065, A2 => n13206, B1 => n8367, B2 => 
                           n13051, ZN => n6602);
   U4336 : OAI22_X1 port map( A1 => n13065, A2 => n13209, B1 => n8350, B2 => 
                           n13051, ZN => n6603);
   U4337 : OAI22_X1 port map( A1 => n13064, A2 => n13212, B1 => n8333, B2 => 
                           n13051, ZN => n6604);
   U4338 : OAI22_X1 port map( A1 => n13064, A2 => n13215, B1 => n8316, B2 => 
                           n13051, ZN => n6605);
   U4339 : OAI22_X1 port map( A1 => n13064, A2 => n13218, B1 => n8299, B2 => 
                           n13051, ZN => n6606);
   U4340 : OAI22_X1 port map( A1 => n13064, A2 => n13221, B1 => n8282, B2 => 
                           n13051, ZN => n6607);
   U4341 : OAI22_X1 port map( A1 => n13064, A2 => n13224, B1 => n8265, B2 => 
                           n13051, ZN => n6608);
   U4342 : OAI22_X1 port map( A1 => n13063, A2 => n13227, B1 => n8248, B2 => 
                           n13051, ZN => n6609);
   U4343 : OAI22_X1 port map( A1 => n13063, A2 => n13230, B1 => n8231, B2 => 
                           n13051, ZN => n6610);
   U4344 : OAI22_X1 port map( A1 => n13063, A2 => n13233, B1 => n8214, B2 => 
                           n13051, ZN => n6611);
   U4345 : OAI22_X1 port map( A1 => n13063, A2 => n13236, B1 => n8197, B2 => 
                           n13051, ZN => n6612);
   U4346 : OAI22_X1 port map( A1 => n13063, A2 => n13239, B1 => n8180, B2 => 
                           n13051, ZN => n6613);
   U4347 : OAI22_X1 port map( A1 => n13045, A2 => n13206, B1 => n8368, B2 => 
                           n13031, ZN => n6538);
   U4348 : OAI22_X1 port map( A1 => n13045, A2 => n13209, B1 => n8351, B2 => 
                           n13031, ZN => n6539);
   U4349 : OAI22_X1 port map( A1 => n13044, A2 => n13212, B1 => n8334, B2 => 
                           n13031, ZN => n6540);
   U4350 : OAI22_X1 port map( A1 => n13044, A2 => n13215, B1 => n8317, B2 => 
                           n13031, ZN => n6541);
   U4351 : OAI22_X1 port map( A1 => n13044, A2 => n13218, B1 => n8300, B2 => 
                           n13031, ZN => n6542);
   U4352 : OAI22_X1 port map( A1 => n13044, A2 => n13221, B1 => n8283, B2 => 
                           n13031, ZN => n6543);
   U4353 : OAI22_X1 port map( A1 => n13044, A2 => n13224, B1 => n8266, B2 => 
                           n13031, ZN => n6544);
   U4354 : OAI22_X1 port map( A1 => n13043, A2 => n13227, B1 => n8249, B2 => 
                           n13031, ZN => n6545);
   U4355 : OAI22_X1 port map( A1 => n13043, A2 => n13230, B1 => n8232, B2 => 
                           n13031, ZN => n6546);
   U4356 : OAI22_X1 port map( A1 => n13043, A2 => n13233, B1 => n8215, B2 => 
                           n13031, ZN => n6547);
   U4357 : OAI22_X1 port map( A1 => n13043, A2 => n13236, B1 => n8198, B2 => 
                           n13031, ZN => n6548);
   U4358 : OAI22_X1 port map( A1 => n13043, A2 => n13239, B1 => n8181, B2 => 
                           n13031, ZN => n6549);
   U4359 : OAI22_X1 port map( A1 => n12922, A2 => n13243, B1 => n8167, B2 => 
                           n12912, ZN => n6166);
   U4360 : OAI22_X1 port map( A1 => n12922, A2 => n13246, B1 => n8150, B2 => 
                           n12912, ZN => n6167);
   U4361 : OAI22_X1 port map( A1 => n12922, A2 => n13249, B1 => n8133, B2 => 
                           n12912, ZN => n6168);
   U4362 : OAI22_X1 port map( A1 => n12922, A2 => n13252, B1 => n8116, B2 => 
                           n12912, ZN => n6169);
   U4363 : OAI22_X1 port map( A1 => n12922, A2 => n13255, B1 => n8099, B2 => 
                           n12912, ZN => n6170);
   U4364 : OAI22_X1 port map( A1 => n12921, A2 => n13258, B1 => n8082, B2 => 
                           n12912, ZN => n6171);
   U4365 : OAI22_X1 port map( A1 => n12921, A2 => n13261, B1 => n8065, B2 => 
                           n12912, ZN => n6172);
   U4366 : OAI22_X1 port map( A1 => n12921, A2 => n13264, B1 => n8048, B2 => 
                           n12912, ZN => n6173);
   U4367 : OAI22_X1 port map( A1 => n12921, A2 => n13267, B1 => n8031, B2 => 
                           n12912, ZN => n6174);
   U4368 : OAI22_X1 port map( A1 => n12921, A2 => n13270, B1 => n8014, B2 => 
                           n12912, ZN => n6175);
   U4369 : OAI22_X1 port map( A1 => n12920, A2 => n13273, B1 => n7997, B2 => 
                           n12912, ZN => n6176);
   U4370 : OAI22_X1 port map( A1 => n12920, A2 => n13276, B1 => n7980, B2 => 
                           n12912, ZN => n6177);
   U4371 : OAI22_X1 port map( A1 => n12920, A2 => n13279, B1 => n7963, B2 => 
                           n12913, ZN => n6178);
   U4372 : OAI22_X1 port map( A1 => n12920, A2 => n13282, B1 => n7946, B2 => 
                           n12913, ZN => n6179);
   U4373 : OAI22_X1 port map( A1 => n12920, A2 => n13285, B1 => n7929, B2 => 
                           n12913, ZN => n6180);
   U4374 : OAI22_X1 port map( A1 => n12919, A2 => n13288, B1 => n7912, B2 => 
                           n12913, ZN => n6181);
   U4375 : OAI22_X1 port map( A1 => n12919, A2 => n13291, B1 => n7895, B2 => 
                           n12913, ZN => n6182);
   U4376 : OAI22_X1 port map( A1 => n12919, A2 => n13294, B1 => n7878, B2 => 
                           n12913, ZN => n6183);
   U4377 : OAI22_X1 port map( A1 => n12919, A2 => n13297, B1 => n7861, B2 => 
                           n12913, ZN => n6184);
   U4378 : OAI22_X1 port map( A1 => n12919, A2 => n13300, B1 => n7844, B2 => 
                           n12913, ZN => n6185);
   U4379 : OAI22_X1 port map( A1 => n12918, A2 => n13303, B1 => n7827, B2 => 
                           n12913, ZN => n6186);
   U4380 : OAI22_X1 port map( A1 => n12918, A2 => n13306, B1 => n7810, B2 => 
                           n12913, ZN => n6187);
   U4381 : OAI22_X1 port map( A1 => n12918, A2 => n13309, B1 => n7793, B2 => 
                           n12913, ZN => n6188);
   U4382 : OAI22_X1 port map( A1 => n12918, A2 => n13312, B1 => n7776, B2 => 
                           n12913, ZN => n6189);
   U4383 : OAI22_X1 port map( A1 => n12918, A2 => n13315, B1 => n7759, B2 => 
                           n12914, ZN => n6190);
   U4384 : OAI22_X1 port map( A1 => n12917, A2 => n13318, B1 => n7742, B2 => 
                           n12914, ZN => n6191);
   U4385 : OAI22_X1 port map( A1 => n12917, A2 => n13321, B1 => n7640, B2 => 
                           n12914, ZN => n6192);
   U4386 : OAI22_X1 port map( A1 => n12917, A2 => n13324, B1 => n7623, B2 => 
                           n12914, ZN => n6193);
   U4387 : OAI22_X1 port map( A1 => n12917, A2 => n13327, B1 => n7519, B2 => 
                           n12914, ZN => n6194);
   U4388 : OAI22_X1 port map( A1 => n12917, A2 => n13330, B1 => n7502, B2 => 
                           n12914, ZN => n6195);
   U4389 : OAI22_X1 port map( A1 => n12916, A2 => n13333, B1 => n7400, B2 => 
                           n12914, ZN => n6196);
   U4390 : OAI22_X1 port map( A1 => n12916, A2 => n13336, B1 => n7383, B2 => 
                           n12914, ZN => n6197);
   U4391 : OAI22_X1 port map( A1 => n12916, A2 => n13339, B1 => n7366, B2 => 
                           n12914, ZN => n6198);
   U4392 : OAI22_X1 port map( A1 => n12916, A2 => n13342, B1 => n7267, B2 => 
                           n12914, ZN => n6199);
   U4393 : OAI22_X1 port map( A1 => n12916, A2 => n13345, B1 => n7250, B2 => 
                           n12914, ZN => n6200);
   U4394 : OAI22_X1 port map( A1 => n12915, A2 => n13348, B1 => n7153, B2 => 
                           n12914, ZN => n6201);
   U4395 : OAI22_X1 port map( A1 => n12942, A2 => n13243, B1 => n8168, B2 => 
                           n12932, ZN => n6230);
   U4396 : OAI22_X1 port map( A1 => n12942, A2 => n13246, B1 => n8151, B2 => 
                           n12932, ZN => n6231);
   U4397 : OAI22_X1 port map( A1 => n12942, A2 => n13249, B1 => n8134, B2 => 
                           n12932, ZN => n6232);
   U4398 : OAI22_X1 port map( A1 => n12942, A2 => n13252, B1 => n8117, B2 => 
                           n12932, ZN => n6233);
   U4399 : OAI22_X1 port map( A1 => n12942, A2 => n13255, B1 => n8100, B2 => 
                           n12932, ZN => n6234);
   U4400 : OAI22_X1 port map( A1 => n12941, A2 => n13258, B1 => n8083, B2 => 
                           n12932, ZN => n6235);
   U4401 : OAI22_X1 port map( A1 => n12941, A2 => n13261, B1 => n8066, B2 => 
                           n12932, ZN => n6236);
   U4402 : OAI22_X1 port map( A1 => n12941, A2 => n13264, B1 => n8049, B2 => 
                           n12932, ZN => n6237);
   U4403 : OAI22_X1 port map( A1 => n12941, A2 => n13267, B1 => n8032, B2 => 
                           n12932, ZN => n6238);
   U4404 : OAI22_X1 port map( A1 => n12941, A2 => n13270, B1 => n8015, B2 => 
                           n12932, ZN => n6239);
   U4405 : OAI22_X1 port map( A1 => n12940, A2 => n13273, B1 => n7998, B2 => 
                           n12932, ZN => n6240);
   U4406 : OAI22_X1 port map( A1 => n12940, A2 => n13276, B1 => n7981, B2 => 
                           n12932, ZN => n6241);
   U4407 : OAI22_X1 port map( A1 => n12940, A2 => n13279, B1 => n7964, B2 => 
                           n12933, ZN => n6242);
   U4408 : OAI22_X1 port map( A1 => n12940, A2 => n13282, B1 => n7947, B2 => 
                           n12933, ZN => n6243);
   U4409 : OAI22_X1 port map( A1 => n12940, A2 => n13285, B1 => n7930, B2 => 
                           n12933, ZN => n6244);
   U4410 : OAI22_X1 port map( A1 => n12939, A2 => n13288, B1 => n7913, B2 => 
                           n12933, ZN => n6245);
   U4411 : OAI22_X1 port map( A1 => n12939, A2 => n13291, B1 => n7896, B2 => 
                           n12933, ZN => n6246);
   U4412 : OAI22_X1 port map( A1 => n12939, A2 => n13294, B1 => n7879, B2 => 
                           n12933, ZN => n6247);
   U4413 : OAI22_X1 port map( A1 => n12939, A2 => n13297, B1 => n7862, B2 => 
                           n12933, ZN => n6248);
   U4414 : OAI22_X1 port map( A1 => n12939, A2 => n13300, B1 => n7845, B2 => 
                           n12933, ZN => n6249);
   U4415 : OAI22_X1 port map( A1 => n12938, A2 => n13303, B1 => n7828, B2 => 
                           n12933, ZN => n6250);
   U4416 : OAI22_X1 port map( A1 => n12938, A2 => n13306, B1 => n7811, B2 => 
                           n12933, ZN => n6251);
   U4417 : OAI22_X1 port map( A1 => n12938, A2 => n13309, B1 => n7794, B2 => 
                           n12933, ZN => n6252);
   U4418 : OAI22_X1 port map( A1 => n12938, A2 => n13312, B1 => n7777, B2 => 
                           n12933, ZN => n6253);
   U4419 : OAI22_X1 port map( A1 => n12938, A2 => n13315, B1 => n7760, B2 => 
                           n12934, ZN => n6254);
   U4420 : OAI22_X1 port map( A1 => n12937, A2 => n13318, B1 => n7743, B2 => 
                           n12934, ZN => n6255);
   U4421 : OAI22_X1 port map( A1 => n12937, A2 => n13321, B1 => n7641, B2 => 
                           n12934, ZN => n6256);
   U4422 : OAI22_X1 port map( A1 => n12937, A2 => n13324, B1 => n7624, B2 => 
                           n12934, ZN => n6257);
   U4423 : OAI22_X1 port map( A1 => n12937, A2 => n13327, B1 => n7520, B2 => 
                           n12934, ZN => n6258);
   U4424 : OAI22_X1 port map( A1 => n12937, A2 => n13330, B1 => n7503, B2 => 
                           n12934, ZN => n6259);
   U4425 : OAI22_X1 port map( A1 => n12936, A2 => n13333, B1 => n7401, B2 => 
                           n12934, ZN => n6260);
   U4426 : OAI22_X1 port map( A1 => n12936, A2 => n13336, B1 => n7384, B2 => 
                           n12934, ZN => n6261);
   U4427 : OAI22_X1 port map( A1 => n12936, A2 => n13339, B1 => n7367, B2 => 
                           n12934, ZN => n6262);
   U4428 : OAI22_X1 port map( A1 => n12936, A2 => n13342, B1 => n7268, B2 => 
                           n12934, ZN => n6263);
   U4429 : OAI22_X1 port map( A1 => n12936, A2 => n13345, B1 => n7251, B2 => 
                           n12934, ZN => n6264);
   U4430 : OAI22_X1 port map( A1 => n12935, A2 => n13348, B1 => n7234, B2 => 
                           n12934, ZN => n6265);
   U4431 : OAI22_X1 port map( A1 => n13022, A2 => n13242, B1 => n8166, B2 => 
                           n13012, ZN => n6486);
   U4432 : OAI22_X1 port map( A1 => n13022, A2 => n13245, B1 => n8149, B2 => 
                           n13012, ZN => n6487);
   U4433 : OAI22_X1 port map( A1 => n13022, A2 => n13248, B1 => n8132, B2 => 
                           n13012, ZN => n6488);
   U4434 : OAI22_X1 port map( A1 => n13022, A2 => n13251, B1 => n8115, B2 => 
                           n13012, ZN => n6489);
   U4435 : OAI22_X1 port map( A1 => n13022, A2 => n13254, B1 => n8098, B2 => 
                           n13012, ZN => n6490);
   U4436 : OAI22_X1 port map( A1 => n13021, A2 => n13257, B1 => n8081, B2 => 
                           n13012, ZN => n6491);
   U4437 : OAI22_X1 port map( A1 => n13021, A2 => n13260, B1 => n8064, B2 => 
                           n13012, ZN => n6492);
   U4438 : OAI22_X1 port map( A1 => n13021, A2 => n13263, B1 => n8047, B2 => 
                           n13012, ZN => n6493);
   U4439 : OAI22_X1 port map( A1 => n13021, A2 => n13266, B1 => n8030, B2 => 
                           n13012, ZN => n6494);
   U4440 : OAI22_X1 port map( A1 => n13021, A2 => n13269, B1 => n8013, B2 => 
                           n13012, ZN => n6495);
   U4441 : OAI22_X1 port map( A1 => n13020, A2 => n13272, B1 => n7996, B2 => 
                           n13012, ZN => n6496);
   U4442 : OAI22_X1 port map( A1 => n13020, A2 => n13275, B1 => n7979, B2 => 
                           n13012, ZN => n6497);
   U4443 : OAI22_X1 port map( A1 => n13020, A2 => n13278, B1 => n7962, B2 => 
                           n13013, ZN => n6498);
   U4444 : OAI22_X1 port map( A1 => n13020, A2 => n13281, B1 => n7945, B2 => 
                           n13013, ZN => n6499);
   U4445 : OAI22_X1 port map( A1 => n13020, A2 => n13284, B1 => n7928, B2 => 
                           n13013, ZN => n6500);
   U4446 : OAI22_X1 port map( A1 => n13019, A2 => n13287, B1 => n7911, B2 => 
                           n13013, ZN => n6501);
   U4447 : OAI22_X1 port map( A1 => n13019, A2 => n13290, B1 => n7894, B2 => 
                           n13013, ZN => n6502);
   U4448 : OAI22_X1 port map( A1 => n13019, A2 => n13293, B1 => n7877, B2 => 
                           n13013, ZN => n6503);
   U4449 : OAI22_X1 port map( A1 => n13019, A2 => n13296, B1 => n7860, B2 => 
                           n13013, ZN => n6504);
   U4450 : OAI22_X1 port map( A1 => n13019, A2 => n13299, B1 => n7843, B2 => 
                           n13013, ZN => n6505);
   U4451 : OAI22_X1 port map( A1 => n13018, A2 => n13302, B1 => n7826, B2 => 
                           n13013, ZN => n6506);
   U4452 : OAI22_X1 port map( A1 => n13018, A2 => n13305, B1 => n7809, B2 => 
                           n13013, ZN => n6507);
   U4453 : OAI22_X1 port map( A1 => n13018, A2 => n13308, B1 => n7792, B2 => 
                           n13013, ZN => n6508);
   U4454 : OAI22_X1 port map( A1 => n13018, A2 => n13311, B1 => n7775, B2 => 
                           n13013, ZN => n6509);
   U4455 : OAI22_X1 port map( A1 => n13018, A2 => n13314, B1 => n7758, B2 => 
                           n13014, ZN => n6510);
   U4456 : OAI22_X1 port map( A1 => n13017, A2 => n13317, B1 => n7656, B2 => 
                           n13014, ZN => n6511);
   U4457 : OAI22_X1 port map( A1 => n13017, A2 => n13320, B1 => n7639, B2 => 
                           n13014, ZN => n6512);
   U4458 : OAI22_X1 port map( A1 => n13017, A2 => n13323, B1 => n7622, B2 => 
                           n13014, ZN => n6513);
   U4459 : OAI22_X1 port map( A1 => n13017, A2 => n13326, B1 => n7518, B2 => 
                           n13014, ZN => n6514);
   U4460 : OAI22_X1 port map( A1 => n13017, A2 => n13329, B1 => n7501, B2 => 
                           n13014, ZN => n6515);
   U4461 : OAI22_X1 port map( A1 => n13016, A2 => n13332, B1 => n7399, B2 => 
                           n13014, ZN => n6516);
   U4462 : OAI22_X1 port map( A1 => n13016, A2 => n13335, B1 => n7382, B2 => 
                           n13014, ZN => n6517);
   U4463 : OAI22_X1 port map( A1 => n13016, A2 => n13338, B1 => n7365, B2 => 
                           n13014, ZN => n6518);
   U4464 : OAI22_X1 port map( A1 => n13016, A2 => n13341, B1 => n7266, B2 => 
                           n13014, ZN => n6519);
   U4465 : OAI22_X1 port map( A1 => n13016, A2 => n13344, B1 => n7249, B2 => 
                           n13014, ZN => n6520);
   U4466 : OAI22_X1 port map( A1 => n13015, A2 => n13347, B1 => n7152, B2 => 
                           n13014, ZN => n6521);
   U4467 : OAI22_X1 port map( A1 => n13002, A2 => n13242, B1 => n8165, B2 => 
                           n12992, ZN => n6422);
   U4468 : OAI22_X1 port map( A1 => n13002, A2 => n13245, B1 => n8148, B2 => 
                           n12992, ZN => n6423);
   U4469 : OAI22_X1 port map( A1 => n13002, A2 => n13248, B1 => n8131, B2 => 
                           n12992, ZN => n6424);
   U4470 : OAI22_X1 port map( A1 => n13002, A2 => n13251, B1 => n8114, B2 => 
                           n12992, ZN => n6425);
   U4471 : OAI22_X1 port map( A1 => n13002, A2 => n13254, B1 => n8097, B2 => 
                           n12992, ZN => n6426);
   U4472 : OAI22_X1 port map( A1 => n13001, A2 => n13257, B1 => n8080, B2 => 
                           n12992, ZN => n6427);
   U4473 : OAI22_X1 port map( A1 => n13001, A2 => n13260, B1 => n8063, B2 => 
                           n12992, ZN => n6428);
   U4474 : OAI22_X1 port map( A1 => n13001, A2 => n13263, B1 => n8046, B2 => 
                           n12992, ZN => n6429);
   U4475 : OAI22_X1 port map( A1 => n13001, A2 => n13266, B1 => n8029, B2 => 
                           n12992, ZN => n6430);
   U4476 : OAI22_X1 port map( A1 => n13001, A2 => n13269, B1 => n8012, B2 => 
                           n12992, ZN => n6431);
   U4477 : OAI22_X1 port map( A1 => n13000, A2 => n13272, B1 => n7995, B2 => 
                           n12992, ZN => n6432);
   U4478 : OAI22_X1 port map( A1 => n13000, A2 => n13275, B1 => n7978, B2 => 
                           n12992, ZN => n6433);
   U4479 : OAI22_X1 port map( A1 => n13000, A2 => n13278, B1 => n7961, B2 => 
                           n12993, ZN => n6434);
   U4480 : OAI22_X1 port map( A1 => n13000, A2 => n13281, B1 => n7944, B2 => 
                           n12993, ZN => n6435);
   U4481 : OAI22_X1 port map( A1 => n13000, A2 => n13284, B1 => n7927, B2 => 
                           n12993, ZN => n6436);
   U4482 : OAI22_X1 port map( A1 => n12999, A2 => n13287, B1 => n7910, B2 => 
                           n12993, ZN => n6437);
   U4483 : OAI22_X1 port map( A1 => n12999, A2 => n13290, B1 => n7893, B2 => 
                           n12993, ZN => n6438);
   U4484 : OAI22_X1 port map( A1 => n12999, A2 => n13293, B1 => n7876, B2 => 
                           n12993, ZN => n6439);
   U4485 : OAI22_X1 port map( A1 => n12999, A2 => n13296, B1 => n7859, B2 => 
                           n12993, ZN => n6440);
   U4486 : OAI22_X1 port map( A1 => n12999, A2 => n13299, B1 => n7842, B2 => 
                           n12993, ZN => n6441);
   U4487 : OAI22_X1 port map( A1 => n12998, A2 => n13302, B1 => n7825, B2 => 
                           n12993, ZN => n6442);
   U4488 : OAI22_X1 port map( A1 => n12998, A2 => n13305, B1 => n7808, B2 => 
                           n12993, ZN => n6443);
   U4489 : OAI22_X1 port map( A1 => n12998, A2 => n13308, B1 => n7791, B2 => 
                           n12993, ZN => n6444);
   U4490 : OAI22_X1 port map( A1 => n12998, A2 => n13311, B1 => n7774, B2 => 
                           n12993, ZN => n6445);
   U4491 : OAI22_X1 port map( A1 => n12998, A2 => n13314, B1 => n7757, B2 => 
                           n12994, ZN => n6446);
   U4492 : OAI22_X1 port map( A1 => n12997, A2 => n13317, B1 => n7655, B2 => 
                           n12994, ZN => n6447);
   U4493 : OAI22_X1 port map( A1 => n12997, A2 => n13320, B1 => n7638, B2 => 
                           n12994, ZN => n6448);
   U4494 : OAI22_X1 port map( A1 => n12997, A2 => n13323, B1 => n7621, B2 => 
                           n12994, ZN => n6449);
   U4495 : OAI22_X1 port map( A1 => n12997, A2 => n13326, B1 => n7517, B2 => 
                           n12994, ZN => n6450);
   U4496 : OAI22_X1 port map( A1 => n12997, A2 => n13329, B1 => n7500, B2 => 
                           n12994, ZN => n6451);
   U4497 : OAI22_X1 port map( A1 => n12996, A2 => n13332, B1 => n7398, B2 => 
                           n12994, ZN => n6452);
   U4498 : OAI22_X1 port map( A1 => n12996, A2 => n13335, B1 => n7381, B2 => 
                           n12994, ZN => n6453);
   U4499 : OAI22_X1 port map( A1 => n12996, A2 => n13338, B1 => n7364, B2 => 
                           n12994, ZN => n6454);
   U4500 : OAI22_X1 port map( A1 => n12996, A2 => n13341, B1 => n7265, B2 => 
                           n12994, ZN => n6455);
   U4501 : OAI22_X1 port map( A1 => n12996, A2 => n13344, B1 => n7248, B2 => 
                           n12994, ZN => n6456);
   U4502 : OAI22_X1 port map( A1 => n12995, A2 => n13347, B1 => n7151, B2 => 
                           n12994, ZN => n6457);
   U4503 : OAI22_X1 port map( A1 => n13062, A2 => n13242, B1 => n8163, B2 => 
                           n13052, ZN => n6614);
   U4504 : OAI22_X1 port map( A1 => n13062, A2 => n13245, B1 => n8146, B2 => 
                           n13052, ZN => n6615);
   U4505 : OAI22_X1 port map( A1 => n13062, A2 => n13248, B1 => n8129, B2 => 
                           n13052, ZN => n6616);
   U4506 : OAI22_X1 port map( A1 => n13062, A2 => n13251, B1 => n8112, B2 => 
                           n13052, ZN => n6617);
   U4507 : OAI22_X1 port map( A1 => n13062, A2 => n13254, B1 => n8095, B2 => 
                           n13052, ZN => n6618);
   U4508 : OAI22_X1 port map( A1 => n13061, A2 => n13257, B1 => n8078, B2 => 
                           n13052, ZN => n6619);
   U4509 : OAI22_X1 port map( A1 => n13061, A2 => n13260, B1 => n8061, B2 => 
                           n13052, ZN => n6620);
   U4510 : OAI22_X1 port map( A1 => n13061, A2 => n13263, B1 => n8044, B2 => 
                           n13052, ZN => n6621);
   U4511 : OAI22_X1 port map( A1 => n13061, A2 => n13266, B1 => n8027, B2 => 
                           n13052, ZN => n6622);
   U4512 : OAI22_X1 port map( A1 => n13061, A2 => n13269, B1 => n8010, B2 => 
                           n13052, ZN => n6623);
   U4513 : OAI22_X1 port map( A1 => n13060, A2 => n13272, B1 => n7993, B2 => 
                           n13052, ZN => n6624);
   U4514 : OAI22_X1 port map( A1 => n13060, A2 => n13275, B1 => n7976, B2 => 
                           n13052, ZN => n6625);
   U4515 : OAI22_X1 port map( A1 => n13060, A2 => n13278, B1 => n7959, B2 => 
                           n13053, ZN => n6626);
   U4516 : OAI22_X1 port map( A1 => n13060, A2 => n13281, B1 => n7942, B2 => 
                           n13053, ZN => n6627);
   U4517 : OAI22_X1 port map( A1 => n13060, A2 => n13284, B1 => n7925, B2 => 
                           n13053, ZN => n6628);
   U4518 : OAI22_X1 port map( A1 => n13059, A2 => n13287, B1 => n7908, B2 => 
                           n13053, ZN => n6629);
   U4519 : OAI22_X1 port map( A1 => n13059, A2 => n13290, B1 => n7891, B2 => 
                           n13053, ZN => n6630);
   U4520 : OAI22_X1 port map( A1 => n13059, A2 => n13293, B1 => n7874, B2 => 
                           n13053, ZN => n6631);
   U4521 : OAI22_X1 port map( A1 => n13059, A2 => n13296, B1 => n7857, B2 => 
                           n13053, ZN => n6632);
   U4522 : OAI22_X1 port map( A1 => n13059, A2 => n13299, B1 => n7840, B2 => 
                           n13053, ZN => n6633);
   U4523 : OAI22_X1 port map( A1 => n13058, A2 => n13302, B1 => n7823, B2 => 
                           n13053, ZN => n6634);
   U4524 : OAI22_X1 port map( A1 => n13058, A2 => n13305, B1 => n7806, B2 => 
                           n13053, ZN => n6635);
   U4525 : OAI22_X1 port map( A1 => n13058, A2 => n13308, B1 => n7789, B2 => 
                           n13053, ZN => n6636);
   U4526 : OAI22_X1 port map( A1 => n13058, A2 => n13311, B1 => n7772, B2 => 
                           n13053, ZN => n6637);
   U4527 : OAI22_X1 port map( A1 => n13058, A2 => n13314, B1 => n7755, B2 => 
                           n13054, ZN => n6638);
   U4528 : OAI22_X1 port map( A1 => n13057, A2 => n13317, B1 => n7653, B2 => 
                           n13054, ZN => n6639);
   U4529 : OAI22_X1 port map( A1 => n13057, A2 => n13320, B1 => n7636, B2 => 
                           n13054, ZN => n6640);
   U4530 : OAI22_X1 port map( A1 => n13057, A2 => n13323, B1 => n7619, B2 => 
                           n13054, ZN => n6641);
   U4531 : OAI22_X1 port map( A1 => n13057, A2 => n13326, B1 => n7515, B2 => 
                           n13054, ZN => n6642);
   U4532 : OAI22_X1 port map( A1 => n13057, A2 => n13329, B1 => n7498, B2 => 
                           n13054, ZN => n6643);
   U4533 : OAI22_X1 port map( A1 => n13056, A2 => n13332, B1 => n7396, B2 => 
                           n13054, ZN => n6644);
   U4534 : OAI22_X1 port map( A1 => n13056, A2 => n13335, B1 => n7379, B2 => 
                           n13054, ZN => n6645);
   U4535 : OAI22_X1 port map( A1 => n13056, A2 => n13338, B1 => n7362, B2 => 
                           n13054, ZN => n6646);
   U4536 : OAI22_X1 port map( A1 => n13056, A2 => n13341, B1 => n7263, B2 => 
                           n13054, ZN => n6647);
   U4537 : OAI22_X1 port map( A1 => n13056, A2 => n13344, B1 => n7246, B2 => 
                           n13054, ZN => n6648);
   U4538 : OAI22_X1 port map( A1 => n13055, A2 => n13347, B1 => n7149, B2 => 
                           n13054, ZN => n6649);
   U4539 : OAI22_X1 port map( A1 => n13042, A2 => n13242, B1 => n8164, B2 => 
                           n13032, ZN => n6550);
   U4540 : OAI22_X1 port map( A1 => n13042, A2 => n13245, B1 => n8147, B2 => 
                           n13032, ZN => n6551);
   U4541 : OAI22_X1 port map( A1 => n13042, A2 => n13248, B1 => n8130, B2 => 
                           n13032, ZN => n6552);
   U4542 : OAI22_X1 port map( A1 => n13042, A2 => n13251, B1 => n8113, B2 => 
                           n13032, ZN => n6553);
   U4543 : OAI22_X1 port map( A1 => n13042, A2 => n13254, B1 => n8096, B2 => 
                           n13032, ZN => n6554);
   U4544 : OAI22_X1 port map( A1 => n13041, A2 => n13257, B1 => n8079, B2 => 
                           n13032, ZN => n6555);
   U4545 : OAI22_X1 port map( A1 => n13041, A2 => n13260, B1 => n8062, B2 => 
                           n13032, ZN => n6556);
   U4546 : OAI22_X1 port map( A1 => n13041, A2 => n13263, B1 => n8045, B2 => 
                           n13032, ZN => n6557);
   U4547 : OAI22_X1 port map( A1 => n13041, A2 => n13266, B1 => n8028, B2 => 
                           n13032, ZN => n6558);
   U4548 : OAI22_X1 port map( A1 => n13041, A2 => n13269, B1 => n8011, B2 => 
                           n13032, ZN => n6559);
   U4549 : OAI22_X1 port map( A1 => n13040, A2 => n13272, B1 => n7994, B2 => 
                           n13032, ZN => n6560);
   U4550 : OAI22_X1 port map( A1 => n13040, A2 => n13275, B1 => n7977, B2 => 
                           n13032, ZN => n6561);
   U4551 : OAI22_X1 port map( A1 => n13040, A2 => n13278, B1 => n7960, B2 => 
                           n13033, ZN => n6562);
   U4552 : OAI22_X1 port map( A1 => n13040, A2 => n13281, B1 => n7943, B2 => 
                           n13033, ZN => n6563);
   U4553 : OAI22_X1 port map( A1 => n13040, A2 => n13284, B1 => n7926, B2 => 
                           n13033, ZN => n6564);
   U4554 : OAI22_X1 port map( A1 => n13039, A2 => n13287, B1 => n7909, B2 => 
                           n13033, ZN => n6565);
   U4555 : OAI22_X1 port map( A1 => n13039, A2 => n13290, B1 => n7892, B2 => 
                           n13033, ZN => n6566);
   U4556 : OAI22_X1 port map( A1 => n13039, A2 => n13293, B1 => n7875, B2 => 
                           n13033, ZN => n6567);
   U4557 : OAI22_X1 port map( A1 => n13039, A2 => n13296, B1 => n7858, B2 => 
                           n13033, ZN => n6568);
   U4558 : OAI22_X1 port map( A1 => n13039, A2 => n13299, B1 => n7841, B2 => 
                           n13033, ZN => n6569);
   U4559 : OAI22_X1 port map( A1 => n13038, A2 => n13302, B1 => n7824, B2 => 
                           n13033, ZN => n6570);
   U4560 : OAI22_X1 port map( A1 => n13038, A2 => n13305, B1 => n7807, B2 => 
                           n13033, ZN => n6571);
   U4561 : OAI22_X1 port map( A1 => n13038, A2 => n13308, B1 => n7790, B2 => 
                           n13033, ZN => n6572);
   U4562 : OAI22_X1 port map( A1 => n13038, A2 => n13311, B1 => n7773, B2 => 
                           n13033, ZN => n6573);
   U4563 : OAI22_X1 port map( A1 => n13038, A2 => n13314, B1 => n7756, B2 => 
                           n13034, ZN => n6574);
   U4564 : OAI22_X1 port map( A1 => n13037, A2 => n13317, B1 => n7654, B2 => 
                           n13034, ZN => n6575);
   U4565 : OAI22_X1 port map( A1 => n13037, A2 => n13320, B1 => n7637, B2 => 
                           n13034, ZN => n6576);
   U4566 : OAI22_X1 port map( A1 => n13037, A2 => n13323, B1 => n7620, B2 => 
                           n13034, ZN => n6577);
   U4567 : OAI22_X1 port map( A1 => n13037, A2 => n13326, B1 => n7516, B2 => 
                           n13034, ZN => n6578);
   U4568 : OAI22_X1 port map( A1 => n13037, A2 => n13329, B1 => n7499, B2 => 
                           n13034, ZN => n6579);
   U4569 : OAI22_X1 port map( A1 => n13036, A2 => n13332, B1 => n7397, B2 => 
                           n13034, ZN => n6580);
   U4570 : OAI22_X1 port map( A1 => n13036, A2 => n13335, B1 => n7380, B2 => 
                           n13034, ZN => n6581);
   U4571 : OAI22_X1 port map( A1 => n13036, A2 => n13338, B1 => n7363, B2 => 
                           n13034, ZN => n6582);
   U4572 : OAI22_X1 port map( A1 => n13036, A2 => n13341, B1 => n7264, B2 => 
                           n13034, ZN => n6583);
   U4573 : OAI22_X1 port map( A1 => n13036, A2 => n13344, B1 => n7247, B2 => 
                           n13034, ZN => n6584);
   U4574 : OAI22_X1 port map( A1 => n13035, A2 => n13347, B1 => n7150, B2 => 
                           n13034, ZN => n6585);
   U4575 : OAI22_X1 port map( A1 => n12865, A2 => n13207, B1 => n8374, B2 => 
                           n12851, ZN => n5962);
   U4576 : OAI22_X1 port map( A1 => n12865, A2 => n13210, B1 => n8357, B2 => 
                           n12851, ZN => n5963);
   U4577 : OAI22_X1 port map( A1 => n12864, A2 => n13213, B1 => n8340, B2 => 
                           n12851, ZN => n5964);
   U4578 : OAI22_X1 port map( A1 => n12864, A2 => n13216, B1 => n8323, B2 => 
                           n12851, ZN => n5965);
   U4579 : OAI22_X1 port map( A1 => n12864, A2 => n13219, B1 => n8306, B2 => 
                           n12851, ZN => n5966);
   U4580 : OAI22_X1 port map( A1 => n12864, A2 => n13222, B1 => n8289, B2 => 
                           n12851, ZN => n5967);
   U4581 : OAI22_X1 port map( A1 => n12864, A2 => n13225, B1 => n8272, B2 => 
                           n12851, ZN => n5968);
   U4582 : OAI22_X1 port map( A1 => n12863, A2 => n13228, B1 => n8255, B2 => 
                           n12851, ZN => n5969);
   U4583 : OAI22_X1 port map( A1 => n12863, A2 => n13231, B1 => n8238, B2 => 
                           n12851, ZN => n5970);
   U4584 : OAI22_X1 port map( A1 => n12863, A2 => n13234, B1 => n8221, B2 => 
                           n12851, ZN => n5971);
   U4585 : OAI22_X1 port map( A1 => n12863, A2 => n13237, B1 => n8204, B2 => 
                           n12851, ZN => n5972);
   U4586 : OAI22_X1 port map( A1 => n12863, A2 => n13240, B1 => n8187, B2 => 
                           n12851, ZN => n5973);
   U4587 : OAI22_X1 port map( A1 => n12862, A2 => n13243, B1 => n8170, B2 => 
                           n12852, ZN => n5974);
   U4588 : OAI22_X1 port map( A1 => n12862, A2 => n13246, B1 => n8153, B2 => 
                           n12852, ZN => n5975);
   U4589 : OAI22_X1 port map( A1 => n12862, A2 => n13249, B1 => n8136, B2 => 
                           n12852, ZN => n5976);
   U4590 : OAI22_X1 port map( A1 => n12862, A2 => n13252, B1 => n8119, B2 => 
                           n12852, ZN => n5977);
   U4591 : OAI22_X1 port map( A1 => n12862, A2 => n13255, B1 => n8102, B2 => 
                           n12852, ZN => n5978);
   U4592 : OAI22_X1 port map( A1 => n12861, A2 => n13258, B1 => n8085, B2 => 
                           n12852, ZN => n5979);
   U4593 : OAI22_X1 port map( A1 => n12861, A2 => n13261, B1 => n8068, B2 => 
                           n12852, ZN => n5980);
   U4594 : OAI22_X1 port map( A1 => n12861, A2 => n13264, B1 => n8051, B2 => 
                           n12852, ZN => n5981);
   U4595 : OAI22_X1 port map( A1 => n12861, A2 => n13267, B1 => n8034, B2 => 
                           n12852, ZN => n5982);
   U4596 : OAI22_X1 port map( A1 => n12861, A2 => n13270, B1 => n8017, B2 => 
                           n12852, ZN => n5983);
   U4597 : OAI22_X1 port map( A1 => n12860, A2 => n13273, B1 => n8000, B2 => 
                           n12852, ZN => n5984);
   U4598 : OAI22_X1 port map( A1 => n12860, A2 => n13276, B1 => n7983, B2 => 
                           n12852, ZN => n5985);
   U4599 : OAI22_X1 port map( A1 => n12860, A2 => n13279, B1 => n7966, B2 => 
                           n12853, ZN => n5986);
   U4600 : OAI22_X1 port map( A1 => n12860, A2 => n13282, B1 => n7949, B2 => 
                           n12853, ZN => n5987);
   U4601 : OAI22_X1 port map( A1 => n12860, A2 => n13285, B1 => n7932, B2 => 
                           n12853, ZN => n5988);
   U4602 : OAI22_X1 port map( A1 => n12859, A2 => n13288, B1 => n7915, B2 => 
                           n12853, ZN => n5989);
   U4603 : OAI22_X1 port map( A1 => n12859, A2 => n13291, B1 => n7898, B2 => 
                           n12853, ZN => n5990);
   U4604 : OAI22_X1 port map( A1 => n12859, A2 => n13294, B1 => n7881, B2 => 
                           n12853, ZN => n5991);
   U4605 : OAI22_X1 port map( A1 => n12859, A2 => n13297, B1 => n7864, B2 => 
                           n12853, ZN => n5992);
   U4606 : OAI22_X1 port map( A1 => n12859, A2 => n13300, B1 => n7847, B2 => 
                           n12853, ZN => n5993);
   U4607 : OAI22_X1 port map( A1 => n12858, A2 => n13303, B1 => n7830, B2 => 
                           n12853, ZN => n5994);
   U4608 : OAI22_X1 port map( A1 => n12858, A2 => n13306, B1 => n7813, B2 => 
                           n12853, ZN => n5995);
   U4609 : OAI22_X1 port map( A1 => n12858, A2 => n13309, B1 => n7796, B2 => 
                           n12853, ZN => n5996);
   U4610 : OAI22_X1 port map( A1 => n12858, A2 => n13312, B1 => n7779, B2 => 
                           n12853, ZN => n5997);
   U4611 : OAI22_X1 port map( A1 => n12858, A2 => n13315, B1 => n7762, B2 => 
                           n12854, ZN => n5998);
   U4612 : OAI22_X1 port map( A1 => n12857, A2 => n13318, B1 => n7745, B2 => 
                           n12854, ZN => n5999);
   U4613 : OAI22_X1 port map( A1 => n12857, A2 => n13321, B1 => n7643, B2 => 
                           n12854, ZN => n6000);
   U4614 : OAI22_X1 port map( A1 => n12857, A2 => n13324, B1 => n7626, B2 => 
                           n12854, ZN => n6001);
   U4615 : OAI22_X1 port map( A1 => n12857, A2 => n13327, B1 => n7522, B2 => 
                           n12854, ZN => n6002);
   U4616 : OAI22_X1 port map( A1 => n12857, A2 => n13330, B1 => n7505, B2 => 
                           n12854, ZN => n6003);
   U4617 : OAI22_X1 port map( A1 => n12856, A2 => n13333, B1 => n7403, B2 => 
                           n12854, ZN => n6004);
   U4618 : OAI22_X1 port map( A1 => n12856, A2 => n13336, B1 => n7386, B2 => 
                           n12854, ZN => n6005);
   U4619 : OAI22_X1 port map( A1 => n12856, A2 => n13339, B1 => n7369, B2 => 
                           n12854, ZN => n6006);
   U4620 : OAI22_X1 port map( A1 => n12856, A2 => n13342, B1 => n7270, B2 => 
                           n12854, ZN => n6007);
   U4621 : OAI22_X1 port map( A1 => n12856, A2 => n13345, B1 => n7253, B2 => 
                           n12854, ZN => n6008);
   U4622 : OAI22_X1 port map( A1 => n12855, A2 => n13348, B1 => n7236, B2 => 
                           n12854, ZN => n6009);
   U4623 : OAI22_X1 port map( A1 => n12842, A2 => n13243, B1 => n8169, B2 => 
                           n12832, ZN => n5910);
   U4624 : OAI22_X1 port map( A1 => n12842, A2 => n13246, B1 => n8152, B2 => 
                           n12832, ZN => n5911);
   U4625 : OAI22_X1 port map( A1 => n12842, A2 => n13249, B1 => n8135, B2 => 
                           n12832, ZN => n5912);
   U4626 : OAI22_X1 port map( A1 => n12842, A2 => n13252, B1 => n8118, B2 => 
                           n12832, ZN => n5913);
   U4627 : OAI22_X1 port map( A1 => n12842, A2 => n13255, B1 => n8101, B2 => 
                           n12832, ZN => n5914);
   U4628 : OAI22_X1 port map( A1 => n12841, A2 => n13258, B1 => n8084, B2 => 
                           n12832, ZN => n5915);
   U4629 : OAI22_X1 port map( A1 => n12841, A2 => n13261, B1 => n8067, B2 => 
                           n12832, ZN => n5916);
   U4630 : OAI22_X1 port map( A1 => n12841, A2 => n13264, B1 => n8050, B2 => 
                           n12832, ZN => n5917);
   U4631 : OAI22_X1 port map( A1 => n12841, A2 => n13267, B1 => n8033, B2 => 
                           n12832, ZN => n5918);
   U4632 : OAI22_X1 port map( A1 => n12841, A2 => n13270, B1 => n8016, B2 => 
                           n12832, ZN => n5919);
   U4633 : OAI22_X1 port map( A1 => n12840, A2 => n13273, B1 => n7999, B2 => 
                           n12832, ZN => n5920);
   U4634 : OAI22_X1 port map( A1 => n12840, A2 => n13276, B1 => n7982, B2 => 
                           n12832, ZN => n5921);
   U4635 : OAI22_X1 port map( A1 => n12840, A2 => n13279, B1 => n7965, B2 => 
                           n12833, ZN => n5922);
   U4636 : OAI22_X1 port map( A1 => n12840, A2 => n13282, B1 => n7948, B2 => 
                           n12833, ZN => n5923);
   U4637 : OAI22_X1 port map( A1 => n12840, A2 => n13285, B1 => n7931, B2 => 
                           n12833, ZN => n5924);
   U4638 : OAI22_X1 port map( A1 => n12839, A2 => n13288, B1 => n7914, B2 => 
                           n12833, ZN => n5925);
   U4639 : OAI22_X1 port map( A1 => n12839, A2 => n13291, B1 => n7897, B2 => 
                           n12833, ZN => n5926);
   U4640 : OAI22_X1 port map( A1 => n12839, A2 => n13294, B1 => n7880, B2 => 
                           n12833, ZN => n5927);
   U4641 : OAI22_X1 port map( A1 => n12839, A2 => n13297, B1 => n7863, B2 => 
                           n12833, ZN => n5928);
   U4642 : OAI22_X1 port map( A1 => n12839, A2 => n13300, B1 => n7846, B2 => 
                           n12833, ZN => n5929);
   U4643 : OAI22_X1 port map( A1 => n12838, A2 => n13303, B1 => n7829, B2 => 
                           n12833, ZN => n5930);
   U4644 : OAI22_X1 port map( A1 => n12838, A2 => n13306, B1 => n7812, B2 => 
                           n12833, ZN => n5931);
   U4645 : OAI22_X1 port map( A1 => n12838, A2 => n13309, B1 => n7795, B2 => 
                           n12833, ZN => n5932);
   U4646 : OAI22_X1 port map( A1 => n12838, A2 => n13312, B1 => n7778, B2 => 
                           n12833, ZN => n5933);
   U4647 : OAI22_X1 port map( A1 => n12838, A2 => n13315, B1 => n7761, B2 => 
                           n12834, ZN => n5934);
   U4648 : OAI22_X1 port map( A1 => n12837, A2 => n13318, B1 => n7744, B2 => 
                           n12834, ZN => n5935);
   U4649 : OAI22_X1 port map( A1 => n12837, A2 => n13321, B1 => n7642, B2 => 
                           n12834, ZN => n5936);
   U4650 : OAI22_X1 port map( A1 => n12837, A2 => n13324, B1 => n7625, B2 => 
                           n12834, ZN => n5937);
   U4651 : OAI22_X1 port map( A1 => n12837, A2 => n13327, B1 => n7521, B2 => 
                           n12834, ZN => n5938);
   U4652 : OAI22_X1 port map( A1 => n12837, A2 => n13330, B1 => n7504, B2 => 
                           n12834, ZN => n5939);
   U4653 : OAI22_X1 port map( A1 => n12836, A2 => n13333, B1 => n7402, B2 => 
                           n12834, ZN => n5940);
   U4654 : OAI22_X1 port map( A1 => n12836, A2 => n13336, B1 => n7385, B2 => 
                           n12834, ZN => n5941);
   U4655 : OAI22_X1 port map( A1 => n12836, A2 => n13339, B1 => n7368, B2 => 
                           n12834, ZN => n5942);
   U4656 : OAI22_X1 port map( A1 => n12836, A2 => n13342, B1 => n7269, B2 => 
                           n12834, ZN => n5943);
   U4657 : OAI22_X1 port map( A1 => n12836, A2 => n13345, B1 => n7252, B2 => 
                           n12834, ZN => n5944);
   U4658 : OAI22_X1 port map( A1 => n12835, A2 => n13348, B1 => n7235, B2 => 
                           n12834, ZN => n5945);
   U4659 : OAI22_X1 port map( A1 => n12782, A2 => n13243, B1 => n8172, B2 => 
                           n12772, ZN => n5718);
   U4660 : OAI22_X1 port map( A1 => n12782, A2 => n13246, B1 => n8155, B2 => 
                           n12772, ZN => n5719);
   U4661 : OAI22_X1 port map( A1 => n12782, A2 => n13249, B1 => n8138, B2 => 
                           n12772, ZN => n5720);
   U4662 : OAI22_X1 port map( A1 => n12782, A2 => n13252, B1 => n8121, B2 => 
                           n12772, ZN => n5721);
   U4663 : OAI22_X1 port map( A1 => n12782, A2 => n13255, B1 => n8104, B2 => 
                           n12772, ZN => n5722);
   U4664 : OAI22_X1 port map( A1 => n12781, A2 => n13258, B1 => n8087, B2 => 
                           n12772, ZN => n5723);
   U4665 : OAI22_X1 port map( A1 => n12781, A2 => n13261, B1 => n8070, B2 => 
                           n12772, ZN => n5724);
   U4666 : OAI22_X1 port map( A1 => n12781, A2 => n13264, B1 => n8053, B2 => 
                           n12772, ZN => n5725);
   U4667 : OAI22_X1 port map( A1 => n12781, A2 => n13267, B1 => n8036, B2 => 
                           n12772, ZN => n5726);
   U4668 : OAI22_X1 port map( A1 => n12781, A2 => n13270, B1 => n8019, B2 => 
                           n12772, ZN => n5727);
   U4669 : OAI22_X1 port map( A1 => n12780, A2 => n13273, B1 => n8002, B2 => 
                           n12772, ZN => n5728);
   U4670 : OAI22_X1 port map( A1 => n12780, A2 => n13276, B1 => n7985, B2 => 
                           n12772, ZN => n5729);
   U4671 : OAI22_X1 port map( A1 => n12780, A2 => n13279, B1 => n7968, B2 => 
                           n12773, ZN => n5730);
   U4672 : OAI22_X1 port map( A1 => n12780, A2 => n13282, B1 => n7951, B2 => 
                           n12773, ZN => n5731);
   U4673 : OAI22_X1 port map( A1 => n12780, A2 => n13285, B1 => n7934, B2 => 
                           n12773, ZN => n5732);
   U4674 : OAI22_X1 port map( A1 => n12779, A2 => n13288, B1 => n7917, B2 => 
                           n12773, ZN => n5733);
   U4675 : OAI22_X1 port map( A1 => n12779, A2 => n13291, B1 => n7900, B2 => 
                           n12773, ZN => n5734);
   U4676 : OAI22_X1 port map( A1 => n12779, A2 => n13294, B1 => n7883, B2 => 
                           n12773, ZN => n5735);
   U4677 : OAI22_X1 port map( A1 => n12779, A2 => n13297, B1 => n7866, B2 => 
                           n12773, ZN => n5736);
   U4678 : OAI22_X1 port map( A1 => n12779, A2 => n13300, B1 => n7849, B2 => 
                           n12773, ZN => n5737);
   U4679 : OAI22_X1 port map( A1 => n12778, A2 => n13303, B1 => n7832, B2 => 
                           n12773, ZN => n5738);
   U4680 : OAI22_X1 port map( A1 => n12778, A2 => n13306, B1 => n7815, B2 => 
                           n12773, ZN => n5739);
   U4681 : OAI22_X1 port map( A1 => n12778, A2 => n13309, B1 => n7798, B2 => 
                           n12773, ZN => n5740);
   U4682 : OAI22_X1 port map( A1 => n12778, A2 => n13312, B1 => n7781, B2 => 
                           n12773, ZN => n5741);
   U4683 : OAI22_X1 port map( A1 => n12778, A2 => n13315, B1 => n7764, B2 => 
                           n12774, ZN => n5742);
   U4684 : OAI22_X1 port map( A1 => n12777, A2 => n13318, B1 => n7747, B2 => 
                           n12774, ZN => n5743);
   U4685 : OAI22_X1 port map( A1 => n12777, A2 => n13321, B1 => n7645, B2 => 
                           n12774, ZN => n5744);
   U4686 : OAI22_X1 port map( A1 => n12777, A2 => n13324, B1 => n7628, B2 => 
                           n12774, ZN => n5745);
   U4687 : OAI22_X1 port map( A1 => n12777, A2 => n13327, B1 => n7524, B2 => 
                           n12774, ZN => n5746);
   U4688 : OAI22_X1 port map( A1 => n12777, A2 => n13330, B1 => n7507, B2 => 
                           n12774, ZN => n5747);
   U4689 : OAI22_X1 port map( A1 => n12776, A2 => n13333, B1 => n7490, B2 => 
                           n12774, ZN => n5748);
   U4690 : OAI22_X1 port map( A1 => n12776, A2 => n13336, B1 => n7388, B2 => 
                           n12774, ZN => n5749);
   U4691 : OAI22_X1 port map( A1 => n12776, A2 => n13339, B1 => n7371, B2 => 
                           n12774, ZN => n5750);
   U4692 : OAI22_X1 port map( A1 => n12776, A2 => n13342, B1 => n7272, B2 => 
                           n12774, ZN => n5751);
   U4693 : OAI22_X1 port map( A1 => n12776, A2 => n13345, B1 => n7255, B2 => 
                           n12774, ZN => n5752);
   U4694 : OAI22_X1 port map( A1 => n12775, A2 => n13348, B1 => n7238, B2 => 
                           n12774, ZN => n5753);
   U4695 : OAI22_X1 port map( A1 => n12762, A2 => n13243, B1 => n8171, B2 => 
                           n12752, ZN => n5654);
   U4696 : OAI22_X1 port map( A1 => n12762, A2 => n13246, B1 => n8154, B2 => 
                           n12752, ZN => n5655);
   U4697 : OAI22_X1 port map( A1 => n12762, A2 => n13249, B1 => n8137, B2 => 
                           n12752, ZN => n5656);
   U4698 : OAI22_X1 port map( A1 => n12762, A2 => n13252, B1 => n8120, B2 => 
                           n12752, ZN => n5657);
   U4699 : OAI22_X1 port map( A1 => n12762, A2 => n13255, B1 => n8103, B2 => 
                           n12752, ZN => n5658);
   U4700 : OAI22_X1 port map( A1 => n12761, A2 => n13258, B1 => n8086, B2 => 
                           n12752, ZN => n5659);
   U4701 : OAI22_X1 port map( A1 => n12761, A2 => n13261, B1 => n8069, B2 => 
                           n12752, ZN => n5660);
   U4702 : OAI22_X1 port map( A1 => n12761, A2 => n13264, B1 => n8052, B2 => 
                           n12752, ZN => n5661);
   U4703 : OAI22_X1 port map( A1 => n12761, A2 => n13267, B1 => n8035, B2 => 
                           n12752, ZN => n5662);
   U4704 : OAI22_X1 port map( A1 => n12761, A2 => n13270, B1 => n8018, B2 => 
                           n12752, ZN => n5663);
   U4705 : OAI22_X1 port map( A1 => n12760, A2 => n13273, B1 => n8001, B2 => 
                           n12752, ZN => n5664);
   U4706 : OAI22_X1 port map( A1 => n12760, A2 => n13276, B1 => n7984, B2 => 
                           n12752, ZN => n5665);
   U4707 : OAI22_X1 port map( A1 => n12760, A2 => n13279, B1 => n7967, B2 => 
                           n12753, ZN => n5666);
   U4708 : OAI22_X1 port map( A1 => n12760, A2 => n13282, B1 => n7950, B2 => 
                           n12753, ZN => n5667);
   U4709 : OAI22_X1 port map( A1 => n12760, A2 => n13285, B1 => n7933, B2 => 
                           n12753, ZN => n5668);
   U4710 : OAI22_X1 port map( A1 => n12759, A2 => n13288, B1 => n7916, B2 => 
                           n12753, ZN => n5669);
   U4711 : OAI22_X1 port map( A1 => n12759, A2 => n13291, B1 => n7899, B2 => 
                           n12753, ZN => n5670);
   U4712 : OAI22_X1 port map( A1 => n12759, A2 => n13294, B1 => n7882, B2 => 
                           n12753, ZN => n5671);
   U4713 : OAI22_X1 port map( A1 => n12759, A2 => n13297, B1 => n7865, B2 => 
                           n12753, ZN => n5672);
   U4714 : OAI22_X1 port map( A1 => n12759, A2 => n13300, B1 => n7848, B2 => 
                           n12753, ZN => n5673);
   U4715 : OAI22_X1 port map( A1 => n12758, A2 => n13303, B1 => n7831, B2 => 
                           n12753, ZN => n5674);
   U4716 : OAI22_X1 port map( A1 => n12758, A2 => n13306, B1 => n7814, B2 => 
                           n12753, ZN => n5675);
   U4717 : OAI22_X1 port map( A1 => n12758, A2 => n13309, B1 => n7797, B2 => 
                           n12753, ZN => n5676);
   U4718 : OAI22_X1 port map( A1 => n12758, A2 => n13312, B1 => n7780, B2 => 
                           n12753, ZN => n5677);
   U4719 : OAI22_X1 port map( A1 => n12758, A2 => n13315, B1 => n7763, B2 => 
                           n12754, ZN => n5678);
   U4720 : OAI22_X1 port map( A1 => n12757, A2 => n13318, B1 => n7746, B2 => 
                           n12754, ZN => n5679);
   U4721 : OAI22_X1 port map( A1 => n12757, A2 => n13321, B1 => n7644, B2 => 
                           n12754, ZN => n5680);
   U4722 : OAI22_X1 port map( A1 => n12757, A2 => n13324, B1 => n7627, B2 => 
                           n12754, ZN => n5681);
   U4723 : OAI22_X1 port map( A1 => n12757, A2 => n13327, B1 => n7523, B2 => 
                           n12754, ZN => n5682);
   U4724 : OAI22_X1 port map( A1 => n12757, A2 => n13330, B1 => n7506, B2 => 
                           n12754, ZN => n5683);
   U4725 : OAI22_X1 port map( A1 => n12756, A2 => n13333, B1 => n7404, B2 => 
                           n12754, ZN => n5684);
   U4726 : OAI22_X1 port map( A1 => n12756, A2 => n13336, B1 => n7387, B2 => 
                           n12754, ZN => n5685);
   U4727 : OAI22_X1 port map( A1 => n12756, A2 => n13339, B1 => n7370, B2 => 
                           n12754, ZN => n5686);
   U4728 : OAI22_X1 port map( A1 => n12756, A2 => n13342, B1 => n7271, B2 => 
                           n12754, ZN => n5687);
   U4729 : OAI22_X1 port map( A1 => n12756, A2 => n13345, B1 => n7254, B2 => 
                           n12754, ZN => n5688);
   U4730 : OAI22_X1 port map( A1 => n12755, A2 => n13348, B1 => n7237, B2 => 
                           n12754, ZN => n5689);
   U4731 : OAI22_X1 port map( A1 => n12588, A2 => n13244, B1 => n8176, B2 => 
                           n12578, ZN => n5078);
   U4732 : OAI22_X1 port map( A1 => n12588, A2 => n13247, B1 => n8159, B2 => 
                           n12578, ZN => n5079);
   U4733 : OAI22_X1 port map( A1 => n12588, A2 => n13250, B1 => n8142, B2 => 
                           n12578, ZN => n5080);
   U4734 : OAI22_X1 port map( A1 => n12588, A2 => n13253, B1 => n8125, B2 => 
                           n12578, ZN => n5081);
   U4735 : OAI22_X1 port map( A1 => n12588, A2 => n13256, B1 => n8108, B2 => 
                           n12578, ZN => n5082);
   U4736 : OAI22_X1 port map( A1 => n12587, A2 => n13259, B1 => n8091, B2 => 
                           n12578, ZN => n5083);
   U4737 : OAI22_X1 port map( A1 => n12587, A2 => n13262, B1 => n8074, B2 => 
                           n12578, ZN => n5084);
   U4738 : OAI22_X1 port map( A1 => n12587, A2 => n13265, B1 => n8057, B2 => 
                           n12578, ZN => n5085);
   U4739 : OAI22_X1 port map( A1 => n12587, A2 => n13268, B1 => n8040, B2 => 
                           n12578, ZN => n5086);
   U4740 : OAI22_X1 port map( A1 => n12587, A2 => n13271, B1 => n8023, B2 => 
                           n12578, ZN => n5087);
   U4741 : OAI22_X1 port map( A1 => n12586, A2 => n13274, B1 => n8006, B2 => 
                           n12578, ZN => n5088);
   U4742 : OAI22_X1 port map( A1 => n12586, A2 => n13277, B1 => n7989, B2 => 
                           n12578, ZN => n5089);
   U4743 : OAI22_X1 port map( A1 => n12586, A2 => n13280, B1 => n7972, B2 => 
                           n12579, ZN => n5090);
   U4744 : OAI22_X1 port map( A1 => n12586, A2 => n13283, B1 => n7955, B2 => 
                           n12579, ZN => n5091);
   U4745 : OAI22_X1 port map( A1 => n12586, A2 => n13286, B1 => n7938, B2 => 
                           n12579, ZN => n5092);
   U4746 : OAI22_X1 port map( A1 => n12585, A2 => n13289, B1 => n7921, B2 => 
                           n12579, ZN => n5093);
   U4747 : OAI22_X1 port map( A1 => n12585, A2 => n13292, B1 => n7904, B2 => 
                           n12579, ZN => n5094);
   U4748 : OAI22_X1 port map( A1 => n12585, A2 => n13295, B1 => n7887, B2 => 
                           n12579, ZN => n5095);
   U4749 : OAI22_X1 port map( A1 => n12585, A2 => n13298, B1 => n7870, B2 => 
                           n12579, ZN => n5096);
   U4750 : OAI22_X1 port map( A1 => n12585, A2 => n13301, B1 => n7853, B2 => 
                           n12579, ZN => n5097);
   U4751 : OAI22_X1 port map( A1 => n12584, A2 => n13304, B1 => n7836, B2 => 
                           n12579, ZN => n5098);
   U4752 : OAI22_X1 port map( A1 => n12584, A2 => n13307, B1 => n7819, B2 => 
                           n12579, ZN => n5099);
   U4753 : OAI22_X1 port map( A1 => n12584, A2 => n13310, B1 => n7802, B2 => 
                           n12579, ZN => n5100);
   U4754 : OAI22_X1 port map( A1 => n12584, A2 => n13313, B1 => n7785, B2 => 
                           n12579, ZN => n5101);
   U4755 : OAI22_X1 port map( A1 => n12584, A2 => n13316, B1 => n7768, B2 => 
                           n12580, ZN => n5102);
   U4756 : OAI22_X1 port map( A1 => n12583, A2 => n13319, B1 => n7751, B2 => 
                           n12580, ZN => n5103);
   U4757 : OAI22_X1 port map( A1 => n12583, A2 => n13322, B1 => n7649, B2 => 
                           n12580, ZN => n5104);
   U4758 : OAI22_X1 port map( A1 => n12583, A2 => n13325, B1 => n7632, B2 => 
                           n12580, ZN => n5105);
   U4759 : OAI22_X1 port map( A1 => n12583, A2 => n13328, B1 => n7528, B2 => 
                           n12580, ZN => n5106);
   U4760 : OAI22_X1 port map( A1 => n12583, A2 => n13331, B1 => n7511, B2 => 
                           n12580, ZN => n5107);
   U4761 : OAI22_X1 port map( A1 => n12582, A2 => n13334, B1 => n7494, B2 => 
                           n12580, ZN => n5108);
   U4762 : OAI22_X1 port map( A1 => n12582, A2 => n13337, B1 => n7392, B2 => 
                           n12580, ZN => n5109);
   U4763 : OAI22_X1 port map( A1 => n12582, A2 => n13340, B1 => n7375, B2 => 
                           n12580, ZN => n5110);
   U4764 : OAI22_X1 port map( A1 => n12582, A2 => n13343, B1 => n7276, B2 => 
                           n12580, ZN => n5111);
   U4765 : OAI22_X1 port map( A1 => n12582, A2 => n13346, B1 => n7259, B2 => 
                           n12580, ZN => n5112);
   U4766 : OAI22_X1 port map( A1 => n12581, A2 => n13349, B1 => n7242, B2 => 
                           n12580, ZN => n5113);
   U4767 : OAI22_X1 port map( A1 => n12645, A2 => n13244, B1 => n8173, B2 => 
                           n12635, ZN => n5270);
   U4768 : OAI22_X1 port map( A1 => n12645, A2 => n13247, B1 => n8156, B2 => 
                           n12635, ZN => n5271);
   U4769 : OAI22_X1 port map( A1 => n12645, A2 => n13250, B1 => n8139, B2 => 
                           n12635, ZN => n5272);
   U4770 : OAI22_X1 port map( A1 => n12645, A2 => n13253, B1 => n8122, B2 => 
                           n12635, ZN => n5273);
   U4771 : OAI22_X1 port map( A1 => n12645, A2 => n13256, B1 => n8105, B2 => 
                           n12635, ZN => n5274);
   U4772 : OAI22_X1 port map( A1 => n12644, A2 => n13259, B1 => n8088, B2 => 
                           n12635, ZN => n5275);
   U4773 : OAI22_X1 port map( A1 => n12644, A2 => n13262, B1 => n8071, B2 => 
                           n12635, ZN => n5276);
   U4774 : OAI22_X1 port map( A1 => n12644, A2 => n13265, B1 => n8054, B2 => 
                           n12635, ZN => n5277);
   U4775 : OAI22_X1 port map( A1 => n12644, A2 => n13268, B1 => n8037, B2 => 
                           n12635, ZN => n5278);
   U4776 : OAI22_X1 port map( A1 => n12644, A2 => n13271, B1 => n8020, B2 => 
                           n12635, ZN => n5279);
   U4777 : OAI22_X1 port map( A1 => n12643, A2 => n13274, B1 => n8003, B2 => 
                           n12635, ZN => n5280);
   U4778 : OAI22_X1 port map( A1 => n12643, A2 => n13277, B1 => n7986, B2 => 
                           n12635, ZN => n5281);
   U4779 : OAI22_X1 port map( A1 => n12643, A2 => n13280, B1 => n7969, B2 => 
                           n12636, ZN => n5282);
   U4780 : OAI22_X1 port map( A1 => n12643, A2 => n13283, B1 => n7952, B2 => 
                           n12636, ZN => n5283);
   U4781 : OAI22_X1 port map( A1 => n12643, A2 => n13286, B1 => n7935, B2 => 
                           n12636, ZN => n5284);
   U4782 : OAI22_X1 port map( A1 => n12642, A2 => n13289, B1 => n7918, B2 => 
                           n12636, ZN => n5285);
   U4783 : OAI22_X1 port map( A1 => n12642, A2 => n13292, B1 => n7901, B2 => 
                           n12636, ZN => n5286);
   U4784 : OAI22_X1 port map( A1 => n12642, A2 => n13295, B1 => n7884, B2 => 
                           n12636, ZN => n5287);
   U4785 : OAI22_X1 port map( A1 => n12642, A2 => n13298, B1 => n7867, B2 => 
                           n12636, ZN => n5288);
   U4786 : OAI22_X1 port map( A1 => n12642, A2 => n13301, B1 => n7850, B2 => 
                           n12636, ZN => n5289);
   U4787 : OAI22_X1 port map( A1 => n12641, A2 => n13304, B1 => n7833, B2 => 
                           n12636, ZN => n5290);
   U4788 : OAI22_X1 port map( A1 => n12641, A2 => n13307, B1 => n7816, B2 => 
                           n12636, ZN => n5291);
   U4789 : OAI22_X1 port map( A1 => n12641, A2 => n13310, B1 => n7799, B2 => 
                           n12636, ZN => n5292);
   U4790 : OAI22_X1 port map( A1 => n12641, A2 => n13313, B1 => n7782, B2 => 
                           n12636, ZN => n5293);
   U4791 : OAI22_X1 port map( A1 => n12641, A2 => n13316, B1 => n7765, B2 => 
                           n12637, ZN => n5294);
   U4792 : OAI22_X1 port map( A1 => n12640, A2 => n13319, B1 => n7748, B2 => 
                           n12637, ZN => n5295);
   U4793 : OAI22_X1 port map( A1 => n12640, A2 => n13322, B1 => n7646, B2 => 
                           n12637, ZN => n5296);
   U4794 : OAI22_X1 port map( A1 => n12640, A2 => n13325, B1 => n7629, B2 => 
                           n12637, ZN => n5297);
   U4795 : OAI22_X1 port map( A1 => n12640, A2 => n13328, B1 => n7525, B2 => 
                           n12637, ZN => n5298);
   U4796 : OAI22_X1 port map( A1 => n12640, A2 => n13331, B1 => n7508, B2 => 
                           n12637, ZN => n5299);
   U4797 : OAI22_X1 port map( A1 => n12639, A2 => n13334, B1 => n7491, B2 => 
                           n12637, ZN => n5300);
   U4798 : OAI22_X1 port map( A1 => n12639, A2 => n13337, B1 => n7389, B2 => 
                           n12637, ZN => n5301);
   U4799 : OAI22_X1 port map( A1 => n12639, A2 => n13340, B1 => n7372, B2 => 
                           n12637, ZN => n5302);
   U4800 : OAI22_X1 port map( A1 => n12639, A2 => n13343, B1 => n7273, B2 => 
                           n12637, ZN => n5303);
   U4801 : OAI22_X1 port map( A1 => n12639, A2 => n13346, B1 => n7256, B2 => 
                           n12637, ZN => n5304);
   U4802 : OAI22_X1 port map( A1 => n12638, A2 => n13349, B1 => n7239, B2 => 
                           n12637, ZN => n5305);
   U4803 : OAI22_X1 port map( A1 => n12664, A2 => n13244, B1 => n8174, B2 => 
                           n12654, ZN => n5334);
   U4804 : OAI22_X1 port map( A1 => n12664, A2 => n13247, B1 => n8157, B2 => 
                           n12654, ZN => n5335);
   U4805 : OAI22_X1 port map( A1 => n12664, A2 => n13250, B1 => n8140, B2 => 
                           n12654, ZN => n5336);
   U4806 : OAI22_X1 port map( A1 => n12664, A2 => n13253, B1 => n8123, B2 => 
                           n12654, ZN => n5337);
   U4807 : OAI22_X1 port map( A1 => n12664, A2 => n13256, B1 => n8106, B2 => 
                           n12654, ZN => n5338);
   U4808 : OAI22_X1 port map( A1 => n12663, A2 => n13259, B1 => n8089, B2 => 
                           n12654, ZN => n5339);
   U4809 : OAI22_X1 port map( A1 => n12663, A2 => n13262, B1 => n8072, B2 => 
                           n12654, ZN => n5340);
   U4810 : OAI22_X1 port map( A1 => n12663, A2 => n13265, B1 => n8055, B2 => 
                           n12654, ZN => n5341);
   U4811 : OAI22_X1 port map( A1 => n12663, A2 => n13268, B1 => n8038, B2 => 
                           n12654, ZN => n5342);
   U4812 : OAI22_X1 port map( A1 => n12663, A2 => n13271, B1 => n8021, B2 => 
                           n12654, ZN => n5343);
   U4813 : OAI22_X1 port map( A1 => n12662, A2 => n13274, B1 => n8004, B2 => 
                           n12654, ZN => n5344);
   U4814 : OAI22_X1 port map( A1 => n12662, A2 => n13277, B1 => n7987, B2 => 
                           n12654, ZN => n5345);
   U4815 : OAI22_X1 port map( A1 => n12662, A2 => n13280, B1 => n7970, B2 => 
                           n12655, ZN => n5346);
   U4816 : OAI22_X1 port map( A1 => n12662, A2 => n13283, B1 => n7953, B2 => 
                           n12655, ZN => n5347);
   U4817 : OAI22_X1 port map( A1 => n12662, A2 => n13286, B1 => n7936, B2 => 
                           n12655, ZN => n5348);
   U4818 : OAI22_X1 port map( A1 => n12661, A2 => n13289, B1 => n7919, B2 => 
                           n12655, ZN => n5349);
   U4819 : OAI22_X1 port map( A1 => n12661, A2 => n13292, B1 => n7902, B2 => 
                           n12655, ZN => n5350);
   U4820 : OAI22_X1 port map( A1 => n12661, A2 => n13295, B1 => n7885, B2 => 
                           n12655, ZN => n5351);
   U4821 : OAI22_X1 port map( A1 => n12661, A2 => n13298, B1 => n7868, B2 => 
                           n12655, ZN => n5352);
   U4822 : OAI22_X1 port map( A1 => n12661, A2 => n13301, B1 => n7851, B2 => 
                           n12655, ZN => n5353);
   U4823 : OAI22_X1 port map( A1 => n12660, A2 => n13304, B1 => n7834, B2 => 
                           n12655, ZN => n5354);
   U4824 : OAI22_X1 port map( A1 => n12660, A2 => n13307, B1 => n7817, B2 => 
                           n12655, ZN => n5355);
   U4825 : OAI22_X1 port map( A1 => n12660, A2 => n13310, B1 => n7800, B2 => 
                           n12655, ZN => n5356);
   U4826 : OAI22_X1 port map( A1 => n12660, A2 => n13313, B1 => n7783, B2 => 
                           n12655, ZN => n5357);
   U4827 : OAI22_X1 port map( A1 => n12660, A2 => n13316, B1 => n7766, B2 => 
                           n12656, ZN => n5358);
   U4828 : OAI22_X1 port map( A1 => n12659, A2 => n13319, B1 => n7749, B2 => 
                           n12656, ZN => n5359);
   U4829 : OAI22_X1 port map( A1 => n12659, A2 => n13322, B1 => n7647, B2 => 
                           n12656, ZN => n5360);
   U4830 : OAI22_X1 port map( A1 => n12659, A2 => n13325, B1 => n7630, B2 => 
                           n12656, ZN => n5361);
   U4831 : OAI22_X1 port map( A1 => n12659, A2 => n13328, B1 => n7526, B2 => 
                           n12656, ZN => n5362);
   U4832 : OAI22_X1 port map( A1 => n12659, A2 => n13331, B1 => n7509, B2 => 
                           n12656, ZN => n5363);
   U4833 : OAI22_X1 port map( A1 => n12658, A2 => n13334, B1 => n7492, B2 => 
                           n12656, ZN => n5364);
   U4834 : OAI22_X1 port map( A1 => n12658, A2 => n13337, B1 => n7390, B2 => 
                           n12656, ZN => n5365);
   U4835 : OAI22_X1 port map( A1 => n12658, A2 => n13340, B1 => n7373, B2 => 
                           n12656, ZN => n5366);
   U4836 : OAI22_X1 port map( A1 => n12658, A2 => n13343, B1 => n7274, B2 => 
                           n12656, ZN => n5367);
   U4837 : OAI22_X1 port map( A1 => n12658, A2 => n13346, B1 => n7257, B2 => 
                           n12656, ZN => n5368);
   U4838 : OAI22_X1 port map( A1 => n12657, A2 => n13349, B1 => n7240, B2 => 
                           n12656, ZN => n5369);
   U4839 : OAI22_X1 port map( A1 => n12855, A2 => n13351, B1 => n7139, B2 => 
                           n12852, ZN => n6010);
   U4840 : OAI22_X1 port map( A1 => n12855, A2 => n13354, B1 => n7122, B2 => 
                           n12853, ZN => n6011);
   U4841 : OAI22_X1 port map( A1 => n12855, A2 => n13357, B1 => n4861, B2 => 
                           n12854, ZN => n6012);
   U4842 : OAI22_X1 port map( A1 => n12855, A2 => n13380, B1 => n4844, B2 => 
                           n12852, ZN => n6013);
   U4843 : OAI22_X1 port map( A1 => n12775, A2 => n13351, B1 => n7141, B2 => 
                           n12772, ZN => n5754);
   U4844 : OAI22_X1 port map( A1 => n12775, A2 => n13354, B1 => n7124, B2 => 
                           n12773, ZN => n5755);
   U4845 : OAI22_X1 port map( A1 => n12775, A2 => n13357, B1 => n7107, B2 => 
                           n12774, ZN => n5756);
   U4846 : OAI22_X1 port map( A1 => n12775, A2 => n13380, B1 => n4846, B2 => 
                           n12772, ZN => n5757);
   U4847 : OAI22_X1 port map( A1 => n12835, A2 => n13351, B1 => n7138, B2 => 
                           n12832, ZN => n5946);
   U4848 : OAI22_X1 port map( A1 => n12835, A2 => n13354, B1 => n7121, B2 => 
                           n12833, ZN => n5947);
   U4849 : OAI22_X1 port map( A1 => n12835, A2 => n13357, B1 => n4860, B2 => 
                           n12834, ZN => n5948);
   U4850 : OAI22_X1 port map( A1 => n12835, A2 => n13380, B1 => n4843, B2 => 
                           n12832, ZN => n5949);
   U4851 : OAI22_X1 port map( A1 => n12755, A2 => n13351, B1 => n7140, B2 => 
                           n12752, ZN => n5690);
   U4852 : OAI22_X1 port map( A1 => n12755, A2 => n13354, B1 => n7123, B2 => 
                           n12753, ZN => n5691);
   U4853 : OAI22_X1 port map( A1 => n12755, A2 => n13357, B1 => n7106, B2 => 
                           n12754, ZN => n5692);
   U4854 : OAI22_X1 port map( A1 => n12755, A2 => n13380, B1 => n4845, B2 => 
                           n12752, ZN => n5693);
   U4855 : OAI22_X1 port map( A1 => n13125, A2 => n13206, B1 => n8366, B2 => 
                           n13111, ZN => n6794);
   U4856 : OAI22_X1 port map( A1 => n12947, A2 => n13171, B1 => n8576, B2 => 
                           n12933, ZN => n6206);
   U4857 : OAI22_X1 port map( A1 => n12947, A2 => n13174, B1 => n8559, B2 => 
                           n12934, ZN => n6207);
   U4858 : OAI22_X1 port map( A1 => n12947, A2 => n13177, B1 => n8542, B2 => 
                           n12931, ZN => n6208);
   U4859 : OAI22_X1 port map( A1 => n12947, A2 => n13180, B1 => n8525, B2 => 
                           n12933, ZN => n6209);
   U4860 : OAI22_X1 port map( A1 => n12946, A2 => n13183, B1 => n8508, B2 => 
                           n12934, ZN => n6210);
   U4861 : OAI22_X1 port map( A1 => n12946, A2 => n13186, B1 => n8491, B2 => 
                           n12930, ZN => n6211);
   U4862 : OAI22_X1 port map( A1 => n12945, A2 => n13210, B1 => n8355, B2 => 
                           n12931, ZN => n6219);
   U4863 : OAI22_X1 port map( A1 => n12944, A2 => n13213, B1 => n8338, B2 => 
                           n12931, ZN => n6220);
   U4864 : OAI22_X1 port map( A1 => n12944, A2 => n13216, B1 => n8321, B2 => 
                           n12931, ZN => n6221);
   U4865 : OAI22_X1 port map( A1 => n12944, A2 => n13219, B1 => n8304, B2 => 
                           n12931, ZN => n6222);
   U4866 : OAI22_X1 port map( A1 => n12944, A2 => n13222, B1 => n8287, B2 => 
                           n12931, ZN => n6223);
   U4867 : OAI22_X1 port map( A1 => n12944, A2 => n13225, B1 => n8270, B2 => 
                           n12931, ZN => n6224);
   U4868 : OAI22_X1 port map( A1 => n12915, A2 => n13351, B1 => n7136, B2 => 
                           n12912, ZN => n6202);
   U4869 : OAI22_X1 port map( A1 => n12915, A2 => n13354, B1 => n7119, B2 => 
                           n12913, ZN => n6203);
   U4870 : OAI22_X1 port map( A1 => n12915, A2 => n13357, B1 => n4858, B2 => 
                           n12914, ZN => n6204);
   U4871 : OAI22_X1 port map( A1 => n12915, A2 => n13380, B1 => n4841, B2 => 
                           n12912, ZN => n6205);
   U4872 : OAI22_X1 port map( A1 => n12935, A2 => n13351, B1 => n7137, B2 => 
                           n12932, ZN => n6266);
   U4873 : OAI22_X1 port map( A1 => n12935, A2 => n13354, B1 => n7120, B2 => 
                           n12933, ZN => n6267);
   U4874 : OAI22_X1 port map( A1 => n12935, A2 => n13357, B1 => n4859, B2 => 
                           n12934, ZN => n6268);
   U4875 : OAI22_X1 port map( A1 => n12935, A2 => n13380, B1 => n4842, B2 => 
                           n12932, ZN => n6269);
   U4876 : OAI22_X1 port map( A1 => n13015, A2 => n13350, B1 => n7135, B2 => 
                           n13012, ZN => n6522);
   U4877 : OAI22_X1 port map( A1 => n13015, A2 => n13353, B1 => n7118, B2 => 
                           n13013, ZN => n6523);
   U4878 : OAI22_X1 port map( A1 => n13015, A2 => n13356, B1 => n4857, B2 => 
                           n13014, ZN => n6524);
   U4879 : OAI22_X1 port map( A1 => n13015, A2 => n13379, B1 => n4840, B2 => 
                           n13012, ZN => n6525);
   U4880 : OAI22_X1 port map( A1 => n12995, A2 => n13350, B1 => n7134, B2 => 
                           n12992, ZN => n6458);
   U4881 : OAI22_X1 port map( A1 => n12995, A2 => n13353, B1 => n7117, B2 => 
                           n12993, ZN => n6459);
   U4882 : OAI22_X1 port map( A1 => n12995, A2 => n13356, B1 => n4856, B2 => 
                           n12994, ZN => n6460);
   U4883 : OAI22_X1 port map( A1 => n12995, A2 => n13379, B1 => n4839, B2 => 
                           n12992, ZN => n6461);
   U4884 : OAI22_X1 port map( A1 => n13055, A2 => n13350, B1 => n7132, B2 => 
                           n13052, ZN => n6650);
   U4885 : OAI22_X1 port map( A1 => n13055, A2 => n13353, B1 => n7115, B2 => 
                           n13053, ZN => n6651);
   U4886 : OAI22_X1 port map( A1 => n13055, A2 => n13356, B1 => n4854, B2 => 
                           n13054, ZN => n6652);
   U4887 : OAI22_X1 port map( A1 => n13055, A2 => n13379, B1 => n4837, B2 => 
                           n13052, ZN => n6653);
   U4888 : OAI22_X1 port map( A1 => n13035, A2 => n13350, B1 => n7133, B2 => 
                           n13032, ZN => n6586);
   U4889 : OAI22_X1 port map( A1 => n13035, A2 => n13353, B1 => n7116, B2 => 
                           n13033, ZN => n6587);
   U4890 : OAI22_X1 port map( A1 => n13035, A2 => n13356, B1 => n4855, B2 => 
                           n13034, ZN => n6588);
   U4891 : OAI22_X1 port map( A1 => n13035, A2 => n13379, B1 => n4838, B2 => 
                           n13032, ZN => n6589);
   U4892 : OAI22_X1 port map( A1 => n12581, A2 => n13352, B1 => n7145, B2 => 
                           n12578, ZN => n5114);
   U4893 : OAI22_X1 port map( A1 => n12581, A2 => n13355, B1 => n7128, B2 => 
                           n12579, ZN => n5115);
   U4894 : OAI22_X1 port map( A1 => n12581, A2 => n13358, B1 => n7111, B2 => 
                           n12580, ZN => n5116);
   U4895 : OAI22_X1 port map( A1 => n12581, A2 => n13381, B1 => n4850, B2 => 
                           n12578, ZN => n5117);
   U4896 : OAI22_X1 port map( A1 => n12638, A2 => n13352, B1 => n7142, B2 => 
                           n12635, ZN => n5306);
   U4897 : OAI22_X1 port map( A1 => n12638, A2 => n13355, B1 => n7125, B2 => 
                           n12636, ZN => n5307);
   U4898 : OAI22_X1 port map( A1 => n12638, A2 => n13358, B1 => n7108, B2 => 
                           n12637, ZN => n5308);
   U4899 : OAI22_X1 port map( A1 => n12638, A2 => n13381, B1 => n4847, B2 => 
                           n12635, ZN => n5309);
   U4900 : OAI22_X1 port map( A1 => n12657, A2 => n13352, B1 => n7143, B2 => 
                           n12654, ZN => n5370);
   U4901 : OAI22_X1 port map( A1 => n12657, A2 => n13355, B1 => n7126, B2 => 
                           n12655, ZN => n5371);
   U4902 : OAI22_X1 port map( A1 => n12657, A2 => n13358, B1 => n7109, B2 => 
                           n12656, ZN => n5372);
   U4903 : OAI22_X1 port map( A1 => n12657, A2 => n13381, B1 => n4848, B2 => 
                           n12654, ZN => n5373);
   U4904 : OAI22_X1 port map( A1 => n13115, A2 => n13379, B1 => n13112, B2 => 
                           n13848, ZN => n6845);
   U4905 : OAI22_X1 port map( A1 => n13135, A2 => n13350, B1 => n13132, B2 => 
                           n13852, ZN => n6906);
   U4906 : OAI22_X1 port map( A1 => n13135, A2 => n13353, B1 => n13133, B2 => 
                           n13851, ZN => n6907);
   U4907 : OAI22_X1 port map( A1 => n13135, A2 => n13356, B1 => n13134, B2 => 
                           n13850, ZN => n6908);
   U4908 : OAI22_X1 port map( A1 => n13135, A2 => n13379, B1 => n13132, B2 => 
                           n13849, ZN => n6909);
   U4909 : OAI22_X1 port map( A1 => n12715, A2 => n13351, B1 => n12713, B2 => 
                           n13666, ZN => n5562);
   U4910 : OAI22_X1 port map( A1 => n12715, A2 => n13354, B1 => n12712, B2 => 
                           n13665, ZN => n5563);
   U4911 : OAI22_X1 port map( A1 => n12715, A2 => n13357, B1 => n12714, B2 => 
                           n13664, ZN => n5564);
   U4912 : OAI22_X1 port map( A1 => n12715, A2 => n13380, B1 => n12713, B2 => 
                           n13663, ZN => n5565);
   U4913 : OAI22_X1 port map( A1 => n12735, A2 => n13351, B1 => n12732, B2 => 
                           n13662, ZN => n5626);
   U4914 : OAI22_X1 port map( A1 => n12735, A2 => n13354, B1 => n12733, B2 => 
                           n13661, ZN => n5627);
   U4915 : OAI22_X1 port map( A1 => n12735, A2 => n13357, B1 => n12734, B2 => 
                           n13660, ZN => n5628);
   U4916 : OAI22_X1 port map( A1 => n12735, A2 => n13380, B1 => n12732, B2 => 
                           n13659, ZN => n5629);
   U4917 : OAI22_X1 port map( A1 => n12795, A2 => n13351, B1 => n12792, B2 => 
                           n13658, ZN => n5818);
   U4918 : OAI22_X1 port map( A1 => n12795, A2 => n13354, B1 => n12793, B2 => 
                           n13657, ZN => n5819);
   U4919 : OAI22_X1 port map( A1 => n12795, A2 => n13357, B1 => n12794, B2 => 
                           n13656, ZN => n5820);
   U4920 : OAI22_X1 port map( A1 => n12795, A2 => n13380, B1 => n12792, B2 => 
                           n13655, ZN => n5821);
   U4921 : OAI22_X1 port map( A1 => n12815, A2 => n13351, B1 => n12812, B2 => 
                           n13654, ZN => n5882);
   U4922 : OAI22_X1 port map( A1 => n12815, A2 => n13354, B1 => n12813, B2 => 
                           n13653, ZN => n5883);
   U4923 : OAI22_X1 port map( A1 => n12815, A2 => n13357, B1 => n12814, B2 => 
                           n13652, ZN => n5884);
   U4924 : OAI22_X1 port map( A1 => n12815, A2 => n13380, B1 => n12812, B2 => 
                           n13651, ZN => n5885);
   U4925 : OAI21_X1 port map( B1 => n4833, B2 => n12544, A => n3180, ZN => 
                           n4926);
   U4926 : OAI21_X1 port map( B1 => n3181, B2 => n3182, A => n12549, ZN => 
                           n3180);
   U4927 : NAND4_X1 port map( A1 => n3183, A2 => n3184, A3 => n3185, A4 => 
                           n3186, ZN => n3182);
   U4928 : NAND4_X1 port map( A1 => n3199, A2 => n3200, A3 => n3201, A4 => 
                           n3202, ZN => n3181);
   U4929 : OAI21_X1 port map( B1 => n4832, B2 => n12543, A => n3161, ZN => 
                           n4927);
   U4930 : OAI21_X1 port map( B1 => n3162, B2 => n3163, A => n12549, ZN => 
                           n3161);
   U4931 : NAND4_X1 port map( A1 => n3164, A2 => n3165, A3 => n3166, A4 => 
                           n3167, ZN => n3163);
   U4932 : NAND4_X1 port map( A1 => n3172, A2 => n3173, A3 => n3174, A4 => 
                           n3175, ZN => n3162);
   U4933 : OAI21_X1 port map( B1 => n4831, B2 => n12544, A => n3142, ZN => 
                           n4928);
   U4934 : OAI21_X1 port map( B1 => n3143, B2 => n3144, A => n12549, ZN => 
                           n3142);
   U4935 : NAND4_X1 port map( A1 => n3145, A2 => n3146, A3 => n3147, A4 => 
                           n3148, ZN => n3144);
   U4936 : NAND4_X1 port map( A1 => n3153, A2 => n3154, A3 => n3155, A4 => 
                           n3156, ZN => n3143);
   U4937 : OAI21_X1 port map( B1 => n4830, B2 => n12543, A => n3123, ZN => 
                           n4929);
   U4938 : OAI21_X1 port map( B1 => n3124, B2 => n3125, A => n12548, ZN => 
                           n3123);
   U4939 : NAND4_X1 port map( A1 => n3126, A2 => n3127, A3 => n3128, A4 => 
                           n3129, ZN => n3125);
   U4940 : NAND4_X1 port map( A1 => n3134, A2 => n3135, A3 => n3136, A4 => 
                           n3137, ZN => n3124);
   U4941 : OAI21_X1 port map( B1 => n4829, B2 => n12543, A => n3104, ZN => 
                           n4930);
   U4942 : OAI21_X1 port map( B1 => n3105, B2 => n3106, A => n12548, ZN => 
                           n3104);
   U4943 : NAND4_X1 port map( A1 => n3107, A2 => n3108, A3 => n3109, A4 => 
                           n3110, ZN => n3106);
   U4944 : NAND4_X1 port map( A1 => n3115, A2 => n3116, A3 => n3117, A4 => 
                           n3118, ZN => n3105);
   U4945 : OAI21_X1 port map( B1 => n4828, B2 => n12544, A => n3085, ZN => 
                           n4931);
   U4946 : OAI21_X1 port map( B1 => n3086, B2 => n3087, A => n12548, ZN => 
                           n3085);
   U4947 : NAND4_X1 port map( A1 => n3088, A2 => n3089, A3 => n3090, A4 => 
                           n3091, ZN => n3087);
   U4948 : NAND4_X1 port map( A1 => n3096, A2 => n3097, A3 => n3098, A4 => 
                           n3099, ZN => n3086);
   U4949 : OAI21_X1 port map( B1 => n4827, B2 => n12544, A => n3066, ZN => 
                           n4932);
   U4950 : OAI21_X1 port map( B1 => n3067, B2 => n3068, A => n12548, ZN => 
                           n3066);
   U4951 : NAND4_X1 port map( A1 => n3069, A2 => n3070, A3 => n3071, A4 => 
                           n3072, ZN => n3068);
   U4952 : NAND4_X1 port map( A1 => n3077, A2 => n3078, A3 => n3079, A4 => 
                           n3080, ZN => n3067);
   U4953 : OAI21_X1 port map( B1 => n4826, B2 => n12543, A => n3047, ZN => 
                           n4933);
   U4954 : OAI21_X1 port map( B1 => n3048, B2 => n3049, A => n12548, ZN => 
                           n3047);
   U4955 : NAND4_X1 port map( A1 => n3050, A2 => n3051, A3 => n3052, A4 => 
                           n3053, ZN => n3049);
   U4956 : NAND4_X1 port map( A1 => n3058, A2 => n3059, A3 => n3060, A4 => 
                           n3061, ZN => n3048);
   U4957 : OAI21_X1 port map( B1 => n4825, B2 => n12543, A => n3028, ZN => 
                           n4934);
   U4958 : OAI21_X1 port map( B1 => n3029, B2 => n3030, A => n12547, ZN => 
                           n3028);
   U4959 : NAND4_X1 port map( A1 => n3031, A2 => n3032, A3 => n3033, A4 => 
                           n3034, ZN => n3030);
   U4960 : NAND4_X1 port map( A1 => n3039, A2 => n3040, A3 => n3041, A4 => 
                           n3042, ZN => n3029);
   U4961 : OAI21_X1 port map( B1 => n4824, B2 => n12543, A => n3009, ZN => 
                           n4935);
   U4962 : OAI21_X1 port map( B1 => n3010, B2 => n3011, A => n12547, ZN => 
                           n3009);
   U4963 : NAND4_X1 port map( A1 => n3012, A2 => n3013, A3 => n3014, A4 => 
                           n3015, ZN => n3011);
   U4964 : NAND4_X1 port map( A1 => n3020, A2 => n3021, A3 => n3022, A4 => 
                           n3023, ZN => n3010);
   U4965 : OAI21_X1 port map( B1 => n4823, B2 => n12542, A => n2990, ZN => 
                           n4936);
   U4966 : OAI21_X1 port map( B1 => n2991, B2 => n2992, A => n12546, ZN => 
                           n2990);
   U4967 : NAND4_X1 port map( A1 => n2993, A2 => n2994, A3 => n2995, A4 => 
                           n2996, ZN => n2992);
   U4968 : NAND4_X1 port map( A1 => n3001, A2 => n3002, A3 => n3003, A4 => 
                           n3004, ZN => n2991);
   U4969 : OAI21_X1 port map( B1 => n4822, B2 => n12543, A => n2971, ZN => 
                           n4937);
   U4970 : OAI21_X1 port map( B1 => n2972, B2 => n2973, A => n12546, ZN => 
                           n2971);
   U4971 : NAND4_X1 port map( A1 => n2974, A2 => n2975, A3 => n2976, A4 => 
                           n2977, ZN => n2973);
   U4972 : NAND4_X1 port map( A1 => n2982, A2 => n2983, A3 => n2984, A4 => 
                           n2985, ZN => n2972);
   U4973 : OAI21_X1 port map( B1 => n4821, B2 => n12543, A => n2952, ZN => 
                           n4938);
   U4974 : OAI21_X1 port map( B1 => n2953, B2 => n2954, A => n12546, ZN => 
                           n2952);
   U4975 : NAND4_X1 port map( A1 => n2955, A2 => n2956, A3 => n2957, A4 => 
                           n2958, ZN => n2954);
   U4976 : NAND4_X1 port map( A1 => n2963, A2 => n2964, A3 => n2965, A4 => 
                           n2966, ZN => n2953);
   U4977 : OAI21_X1 port map( B1 => n4820, B2 => n12543, A => n2933, ZN => 
                           n4939);
   U4978 : OAI21_X1 port map( B1 => n2934, B2 => n2935, A => n12545, ZN => 
                           n2933);
   U4979 : NAND4_X1 port map( A1 => n2936, A2 => n2937, A3 => n2938, A4 => 
                           n2939, ZN => n2935);
   U4980 : NAND4_X1 port map( A1 => n2944, A2 => n2945, A3 => n2946, A4 => 
                           n2947, ZN => n2934);
   U4981 : OAI21_X1 port map( B1 => n4819, B2 => n12543, A => n2914, ZN => 
                           n4940);
   U4982 : OAI21_X1 port map( B1 => n2915, B2 => n2916, A => n12547, ZN => 
                           n2914);
   U4983 : NAND4_X1 port map( A1 => n2917, A2 => n2918, A3 => n2919, A4 => 
                           n2920, ZN => n2916);
   U4984 : NAND4_X1 port map( A1 => n2925, A2 => n2926, A3 => n2927, A4 => 
                           n2928, ZN => n2915);
   U4985 : OAI21_X1 port map( B1 => n4818, B2 => n12543, A => n2895, ZN => 
                           n4941);
   U4986 : OAI21_X1 port map( B1 => n2896, B2 => n2897, A => n12546, ZN => 
                           n2895);
   U4987 : NAND4_X1 port map( A1 => n2898, A2 => n2899, A3 => n2900, A4 => 
                           n2901, ZN => n2897);
   U4988 : NAND4_X1 port map( A1 => n2906, A2 => n2907, A3 => n2908, A4 => 
                           n2909, ZN => n2896);
   U4989 : OAI21_X1 port map( B1 => n4817, B2 => n12542, A => n2876, ZN => 
                           n4942);
   U4990 : OAI21_X1 port map( B1 => n2877, B2 => n2878, A => n12544, ZN => 
                           n2876);
   U4991 : NAND4_X1 port map( A1 => n2879, A2 => n2880, A3 => n2881, A4 => 
                           n2882, ZN => n2878);
   U4992 : NAND4_X1 port map( A1 => n2887, A2 => n2888, A3 => n2889, A4 => 
                           n2890, ZN => n2877);
   U4993 : OAI21_X1 port map( B1 => n4816, B2 => n12542, A => n2857, ZN => 
                           n4943);
   U4994 : OAI21_X1 port map( B1 => n2858, B2 => n2859, A => n12546, ZN => 
                           n2857);
   U4995 : NAND4_X1 port map( A1 => n2860, A2 => n2861, A3 => n2862, A4 => 
                           n2863, ZN => n2859);
   U4996 : NAND4_X1 port map( A1 => n2868, A2 => n2869, A3 => n2870, A4 => 
                           n2871, ZN => n2858);
   U4997 : OAI21_X1 port map( B1 => n4815, B2 => n12543, A => n2838, ZN => 
                           n4944);
   U4998 : OAI21_X1 port map( B1 => n2839, B2 => n2840, A => n12545, ZN => 
                           n2838);
   U4999 : NAND4_X1 port map( A1 => n2841, A2 => n2842, A3 => n2843, A4 => 
                           n2844, ZN => n2840);
   U5000 : NAND4_X1 port map( A1 => n2849, A2 => n2850, A3 => n2851, A4 => 
                           n2852, ZN => n2839);
   U5001 : OAI21_X1 port map( B1 => n4814, B2 => n12542, A => n2819, ZN => 
                           n4945);
   U5002 : OAI21_X1 port map( B1 => n2820, B2 => n2821, A => n12546, ZN => 
                           n2819);
   U5003 : NAND4_X1 port map( A1 => n2822, A2 => n2823, A3 => n2824, A4 => 
                           n2825, ZN => n2821);
   U5004 : NAND4_X1 port map( A1 => n2830, A2 => n2831, A3 => n2832, A4 => 
                           n2833, ZN => n2820);
   U5005 : OAI21_X1 port map( B1 => n4813, B2 => n12542, A => n2800, ZN => 
                           n4946);
   U5006 : OAI21_X1 port map( B1 => n2801, B2 => n2802, A => n12544, ZN => 
                           n2800);
   U5007 : NAND4_X1 port map( A1 => n2803, A2 => n2804, A3 => n2805, A4 => 
                           n2806, ZN => n2802);
   U5008 : NAND4_X1 port map( A1 => n2811, A2 => n2812, A3 => n2813, A4 => 
                           n2814, ZN => n2801);
   U5009 : OAI21_X1 port map( B1 => n4812, B2 => n12542, A => n2781, ZN => 
                           n4947);
   U5010 : OAI21_X1 port map( B1 => n2782, B2 => n2783, A => n12545, ZN => 
                           n2781);
   U5011 : NAND4_X1 port map( A1 => n2784, A2 => n2785, A3 => n2786, A4 => 
                           n2787, ZN => n2783);
   U5012 : NAND4_X1 port map( A1 => n2792, A2 => n2793, A3 => n2794, A4 => 
                           n2795, ZN => n2782);
   U5013 : OAI21_X1 port map( B1 => n4811, B2 => n12542, A => n2762, ZN => 
                           n4948);
   U5014 : OAI21_X1 port map( B1 => n2763, B2 => n2764, A => n12544, ZN => 
                           n2762);
   U5015 : NAND4_X1 port map( A1 => n2765, A2 => n2766, A3 => n2767, A4 => 
                           n2768, ZN => n2764);
   U5016 : NAND4_X1 port map( A1 => n2773, A2 => n2774, A3 => n2775, A4 => 
                           n2776, ZN => n2763);
   U5017 : OAI21_X1 port map( B1 => n4810, B2 => n12542, A => n2743, ZN => 
                           n4949);
   U5018 : OAI21_X1 port map( B1 => n2744, B2 => n2745, A => n12545, ZN => 
                           n2743);
   U5019 : NAND4_X1 port map( A1 => n2746, A2 => n2747, A3 => n2748, A4 => 
                           n2749, ZN => n2745);
   U5020 : NAND4_X1 port map( A1 => n2754, A2 => n2755, A3 => n2756, A4 => 
                           n2757, ZN => n2744);
   U5021 : OAI21_X1 port map( B1 => n4809, B2 => n12542, A => n2724, ZN => 
                           n4950);
   U5022 : OAI21_X1 port map( B1 => n2725, B2 => n2726, A => n12544, ZN => 
                           n2724);
   U5023 : NAND4_X1 port map( A1 => n2727, A2 => n2728, A3 => n2729, A4 => 
                           n2730, ZN => n2726);
   U5024 : NAND4_X1 port map( A1 => n2735, A2 => n2736, A3 => n2737, A4 => 
                           n2738, ZN => n2725);
   U5025 : OAI21_X1 port map( B1 => n4808, B2 => n12542, A => n2705, ZN => 
                           n4951);
   U5026 : OAI21_X1 port map( B1 => n2706, B2 => n2707, A => n12545, ZN => 
                           n2705);
   U5027 : NAND4_X1 port map( A1 => n2708, A2 => n2709, A3 => n2710, A4 => 
                           n2711, ZN => n2707);
   U5028 : NAND4_X1 port map( A1 => n2716, A2 => n2717, A3 => n2718, A4 => 
                           n2719, ZN => n2706);
   U5029 : OAI21_X1 port map( B1 => n4807, B2 => n12542, A => n2686, ZN => 
                           n4952);
   U5030 : OAI21_X1 port map( B1 => n2687, B2 => n2688, A => n12545, ZN => 
                           n2686);
   U5031 : NAND4_X1 port map( A1 => n2689, A2 => n2690, A3 => n2691, A4 => 
                           n2692, ZN => n2688);
   U5032 : NAND4_X1 port map( A1 => n2697, A2 => n2698, A3 => n2699, A4 => 
                           n2700, ZN => n2687);
   U5033 : OAI21_X1 port map( B1 => n4806, B2 => n12541, A => n2667, ZN => 
                           n4953);
   U5034 : OAI21_X1 port map( B1 => n2668, B2 => n2669, A => n12544, ZN => 
                           n2667);
   U5035 : NAND4_X1 port map( A1 => n2670, A2 => n2671, A3 => n2672, A4 => 
                           n2673, ZN => n2669);
   U5036 : NAND4_X1 port map( A1 => n2678, A2 => n2679, A3 => n2680, A4 => 
                           n2681, ZN => n2668);
   U5037 : OAI21_X1 port map( B1 => n4805, B2 => n12541, A => n2648, ZN => 
                           n4954);
   U5038 : OAI21_X1 port map( B1 => n2649, B2 => n2650, A => n12544, ZN => 
                           n2648);
   U5039 : NAND4_X1 port map( A1 => n2651, A2 => n2652, A3 => n2653, A4 => 
                           n2654, ZN => n2650);
   U5040 : NAND4_X1 port map( A1 => n2659, A2 => n2660, A3 => n2661, A4 => 
                           n2662, ZN => n2649);
   U5041 : OAI21_X1 port map( B1 => n4804, B2 => n12541, A => n2629, ZN => 
                           n4955);
   U5042 : OAI21_X1 port map( B1 => n2630, B2 => n2631, A => n12545, ZN => 
                           n2629);
   U5043 : NAND4_X1 port map( A1 => n2632, A2 => n2633, A3 => n2634, A4 => 
                           n2635, ZN => n2631);
   U5044 : NAND4_X1 port map( A1 => n2640, A2 => n2641, A3 => n2642, A4 => 
                           n2643, ZN => n2630);
   U5045 : OAI21_X1 port map( B1 => n4803, B2 => n12541, A => n2610, ZN => 
                           n4956);
   U5046 : OAI21_X1 port map( B1 => n2611, B2 => n2612, A => n12544, ZN => 
                           n2610);
   U5047 : NAND4_X1 port map( A1 => n2613, A2 => n2614, A3 => n2615, A4 => 
                           n2616, ZN => n2612);
   U5048 : NAND4_X1 port map( A1 => n2621, A2 => n2622, A3 => n2623, A4 => 
                           n2624, ZN => n2611);
   U5049 : OAI21_X1 port map( B1 => n4797, B2 => n12542, A => n2591, ZN => 
                           n4957);
   U5050 : OAI21_X1 port map( B1 => n2592, B2 => n2593, A => n12544, ZN => 
                           n2591);
   U5051 : NAND4_X1 port map( A1 => n2594, A2 => n2595, A3 => n2596, A4 => 
                           n2597, ZN => n2593);
   U5052 : NAND4_X1 port map( A1 => n2602, A2 => n2603, A3 => n2604, A4 => 
                           n2605, ZN => n2592);
   U5053 : OAI21_X1 port map( B1 => n4796, B2 => n12541, A => n2572, ZN => 
                           n4958);
   U5054 : OAI21_X1 port map( B1 => n2573, B2 => n2574, A => n12545, ZN => 
                           n2572);
   U5055 : NAND4_X1 port map( A1 => n2575, A2 => n2576, A3 => n2577, A4 => 
                           n2578, ZN => n2574);
   U5056 : NAND4_X1 port map( A1 => n2583, A2 => n2584, A3 => n2585, A4 => 
                           n2586, ZN => n2573);
   U5057 : OAI21_X1 port map( B1 => n4795, B2 => n12541, A => n2553, ZN => 
                           n4959);
   U5058 : OAI21_X1 port map( B1 => n2554, B2 => n2555, A => n12545, ZN => 
                           n2553);
   U5059 : NAND4_X1 port map( A1 => n2556, A2 => n2557, A3 => n2558, A4 => 
                           n2559, ZN => n2555);
   U5060 : NAND4_X1 port map( A1 => n2564, A2 => n2565, A3 => n2566, A4 => 
                           n2567, ZN => n2554);
   U5061 : OAI21_X1 port map( B1 => n4794, B2 => n12541, A => n2534, ZN => 
                           n4960);
   U5062 : OAI21_X1 port map( B1 => n2535, B2 => n2536, A => n12545, ZN => 
                           n2534);
   U5063 : NAND4_X1 port map( A1 => n2537, A2 => n2538, A3 => n2539, A4 => 
                           n2540, ZN => n2536);
   U5064 : NAND4_X1 port map( A1 => n2545, A2 => n2546, A3 => n2547, A4 => 
                           n2548, ZN => n2535);
   U5065 : OAI21_X1 port map( B1 => n4793, B2 => n12541, A => n2515, ZN => 
                           n4961);
   U5066 : OAI21_X1 port map( B1 => n2516, B2 => n2517, A => n12546, ZN => 
                           n2515);
   U5067 : NAND4_X1 port map( A1 => n2518, A2 => n2519, A3 => n2520, A4 => 
                           n2521, ZN => n2517);
   U5068 : NAND4_X1 port map( A1 => n2526, A2 => n2527, A3 => n2528, A4 => 
                           n2529, ZN => n2516);
   U5069 : OAI21_X1 port map( B1 => n4792, B2 => n12541, A => n2496, ZN => 
                           n4962);
   U5070 : OAI21_X1 port map( B1 => n2497, B2 => n2498, A => n12545, ZN => 
                           n2496);
   U5071 : NAND4_X1 port map( A1 => n2499, A2 => n2500, A3 => n2501, A4 => 
                           n2502, ZN => n2498);
   U5072 : NAND4_X1 port map( A1 => n2507, A2 => n2508, A3 => n2509, A4 => 
                           n2510, ZN => n2497);
   U5073 : OAI21_X1 port map( B1 => n4791, B2 => n12541, A => n2477, ZN => 
                           n4963);
   U5074 : OAI21_X1 port map( B1 => n2478, B2 => n2479, A => n12545, ZN => 
                           n2477);
   U5075 : NAND4_X1 port map( A1 => n2480, A2 => n2481, A3 => n2482, A4 => 
                           n2483, ZN => n2479);
   U5076 : NAND4_X1 port map( A1 => n2488, A2 => n2489, A3 => n2490, A4 => 
                           n2491, ZN => n2478);
   U5077 : OAI21_X1 port map( B1 => n4790, B2 => n12541, A => n2458, ZN => 
                           n4964);
   U5078 : OAI21_X1 port map( B1 => n2459, B2 => n2460, A => n12547, ZN => 
                           n2458);
   U5079 : NAND4_X1 port map( A1 => n2461, A2 => n2462, A3 => n2463, A4 => 
                           n2464, ZN => n2460);
   U5080 : NAND4_X1 port map( A1 => n2469, A2 => n2470, A3 => n2471, A4 => 
                           n2472, ZN => n2459);
   U5081 : OAI21_X1 port map( B1 => n4789, B2 => n12540, A => n2439, ZN => 
                           n4965);
   U5082 : OAI21_X1 port map( B1 => n2440, B2 => n2441, A => n12547, ZN => 
                           n2439);
   U5083 : NAND4_X1 port map( A1 => n2442, A2 => n2443, A3 => n2444, A4 => 
                           n2445, ZN => n2441);
   U5084 : NAND4_X1 port map( A1 => n2450, A2 => n2451, A3 => n2452, A4 => 
                           n2453, ZN => n2440);
   U5085 : OAI21_X1 port map( B1 => n4788, B2 => n12540, A => n2420, ZN => 
                           n4966);
   U5086 : OAI21_X1 port map( B1 => n2421, B2 => n2422, A => n12546, ZN => 
                           n2420);
   U5087 : NAND4_X1 port map( A1 => n2423, A2 => n2424, A3 => n2425, A4 => 
                           n2426, ZN => n2422);
   U5088 : NAND4_X1 port map( A1 => n2431, A2 => n2432, A3 => n2433, A4 => 
                           n2434, ZN => n2421);
   U5089 : OAI21_X1 port map( B1 => n4787, B2 => n12540, A => n2401, ZN => 
                           n4967);
   U5090 : OAI21_X1 port map( B1 => n2402, B2 => n2403, A => n12546, ZN => 
                           n2401);
   U5091 : NAND4_X1 port map( A1 => n2404, A2 => n2405, A3 => n2406, A4 => 
                           n2407, ZN => n2403);
   U5092 : NAND4_X1 port map( A1 => n2412, A2 => n2413, A3 => n2414, A4 => 
                           n2415, ZN => n2402);
   U5093 : OAI21_X1 port map( B1 => n4786, B2 => n12540, A => n2382, ZN => 
                           n4968);
   U5094 : OAI21_X1 port map( B1 => n2383, B2 => n2384, A => n12546, ZN => 
                           n2382);
   U5095 : NAND4_X1 port map( A1 => n2385, A2 => n2386, A3 => n2387, A4 => 
                           n2388, ZN => n2384);
   U5096 : NAND4_X1 port map( A1 => n2393, A2 => n2394, A3 => n2395, A4 => 
                           n2396, ZN => n2383);
   U5097 : OAI21_X1 port map( B1 => n4785, B2 => n12540, A => n2363, ZN => 
                           n4969);
   U5098 : OAI21_X1 port map( B1 => n2364, B2 => n2365, A => n12546, ZN => 
                           n2363);
   U5099 : NAND4_X1 port map( A1 => n2366, A2 => n2367, A3 => n2368, A4 => 
                           n2369, ZN => n2365);
   U5100 : NAND4_X1 port map( A1 => n2374, A2 => n2375, A3 => n2376, A4 => 
                           n2377, ZN => n2364);
   U5101 : OAI21_X1 port map( B1 => n4784, B2 => n12540, A => n2344, ZN => 
                           n4970);
   U5102 : OAI21_X1 port map( B1 => n2345, B2 => n2346, A => n12547, ZN => 
                           n2344);
   U5103 : NAND4_X1 port map( A1 => n2347, A2 => n2348, A3 => n2349, A4 => 
                           n2350, ZN => n2346);
   U5104 : NAND4_X1 port map( A1 => n2355, A2 => n2356, A3 => n2357, A4 => 
                           n2358, ZN => n2345);
   U5105 : OAI21_X1 port map( B1 => n4783, B2 => n12540, A => n2325, ZN => 
                           n4971);
   U5106 : OAI21_X1 port map( B1 => n2326, B2 => n2327, A => n12546, ZN => 
                           n2325);
   U5107 : NAND4_X1 port map( A1 => n2328, A2 => n2329, A3 => n2330, A4 => 
                           n2331, ZN => n2327);
   U5108 : NAND4_X1 port map( A1 => n2336, A2 => n2337, A3 => n2338, A4 => 
                           n2339, ZN => n2326);
   U5109 : OAI21_X1 port map( B1 => n4782, B2 => n12540, A => n2306, ZN => 
                           n4972);
   U5110 : OAI21_X1 port map( B1 => n2307, B2 => n2308, A => n12547, ZN => 
                           n2306);
   U5111 : NAND4_X1 port map( A1 => n2309, A2 => n2310, A3 => n2311, A4 => 
                           n2312, ZN => n2308);
   U5112 : NAND4_X1 port map( A1 => n2317, A2 => n2318, A3 => n2319, A4 => 
                           n2320, ZN => n2307);
   U5113 : OAI21_X1 port map( B1 => n4781, B2 => n12540, A => n2287, ZN => 
                           n4973);
   U5114 : OAI21_X1 port map( B1 => n2288, B2 => n2289, A => n12547, ZN => 
                           n2287);
   U5115 : NAND4_X1 port map( A1 => n2290, A2 => n2291, A3 => n2292, A4 => 
                           n2293, ZN => n2289);
   U5116 : NAND4_X1 port map( A1 => n2298, A2 => n2299, A3 => n2300, A4 => 
                           n2301, ZN => n2288);
   U5117 : OAI21_X1 port map( B1 => n4780, B2 => n12540, A => n2268, ZN => 
                           n4974);
   U5118 : OAI21_X1 port map( B1 => n2269, B2 => n2270, A => n12547, ZN => 
                           n2268);
   U5119 : NAND4_X1 port map( A1 => n2271, A2 => n2272, A3 => n2273, A4 => 
                           n2274, ZN => n2270);
   U5120 : NAND4_X1 port map( A1 => n2279, A2 => n2280, A3 => n2281, A4 => 
                           n2282, ZN => n2269);
   U5121 : OAI21_X1 port map( B1 => n4779, B2 => n12540, A => n2249, ZN => 
                           n4975);
   U5122 : OAI21_X1 port map( B1 => n2250, B2 => n2251, A => n12547, ZN => 
                           n2249);
   U5123 : NAND4_X1 port map( A1 => n2252, A2 => n2253, A3 => n2254, A4 => 
                           n2255, ZN => n2251);
   U5124 : NAND4_X1 port map( A1 => n2260, A2 => n2261, A3 => n2262, A4 => 
                           n2263, ZN => n2250);
   U5125 : OAI21_X1 port map( B1 => n4778, B2 => n12540, A => n2230, ZN => 
                           n4976);
   U5126 : OAI21_X1 port map( B1 => n2231, B2 => n2232, A => n12548, ZN => 
                           n2230);
   U5127 : NAND4_X1 port map( A1 => n2233, A2 => n2234, A3 => n2235, A4 => 
                           n2236, ZN => n2232);
   U5128 : NAND4_X1 port map( A1 => n2241, A2 => n2242, A3 => n2243, A4 => 
                           n2244, ZN => n2231);
   U5129 : OAI21_X1 port map( B1 => n4777, B2 => n12539, A => n2211, ZN => 
                           n4977);
   U5130 : OAI21_X1 port map( B1 => n2212, B2 => n2213, A => n12547, ZN => 
                           n2211);
   U5131 : NAND4_X1 port map( A1 => n2214, A2 => n2215, A3 => n2216, A4 => 
                           n2217, ZN => n2213);
   U5132 : NAND4_X1 port map( A1 => n2222, A2 => n2223, A3 => n2224, A4 => 
                           n2225, ZN => n2212);
   U5133 : OAI21_X1 port map( B1 => n4776, B2 => n12539, A => n2192, ZN => 
                           n4978);
   U5134 : OAI21_X1 port map( B1 => n2193, B2 => n2194, A => n12547, ZN => 
                           n2192);
   U5135 : NAND4_X1 port map( A1 => n2195, A2 => n2196, A3 => n2197, A4 => 
                           n2198, ZN => n2194);
   U5136 : NAND4_X1 port map( A1 => n2203, A2 => n2204, A3 => n2205, A4 => 
                           n2206, ZN => n2193);
   U5137 : OAI21_X1 port map( B1 => n4775, B2 => n12539, A => n2173, ZN => 
                           n4979);
   U5138 : OAI21_X1 port map( B1 => n2174, B2 => n2175, A => n12548, ZN => 
                           n2173);
   U5139 : NAND4_X1 port map( A1 => n2176, A2 => n2177, A3 => n2178, A4 => 
                           n2179, ZN => n2175);
   U5140 : NAND4_X1 port map( A1 => n2184, A2 => n2185, A3 => n2186, A4 => 
                           n2187, ZN => n2174);
   U5141 : OAI21_X1 port map( B1 => n4774, B2 => n12539, A => n2154, ZN => 
                           n4980);
   U5142 : OAI21_X1 port map( B1 => n2155, B2 => n2156, A => n12548, ZN => 
                           n2154);
   U5143 : NAND4_X1 port map( A1 => n2157, A2 => n2158, A3 => n2159, A4 => 
                           n2160, ZN => n2156);
   U5144 : NAND4_X1 port map( A1 => n2165, A2 => n2166, A3 => n2167, A4 => 
                           n2168, ZN => n2155);
   U5145 : OAI21_X1 port map( B1 => n4773, B2 => n12539, A => n2135, ZN => 
                           n4981);
   U5146 : OAI21_X1 port map( B1 => n2136, B2 => n2137, A => n12548, ZN => 
                           n2135);
   U5147 : NAND4_X1 port map( A1 => n2138, A2 => n2139, A3 => n2140, A4 => 
                           n2141, ZN => n2137);
   U5148 : NAND4_X1 port map( A1 => n2146, A2 => n2147, A3 => n2148, A4 => 
                           n2149, ZN => n2136);
   U5149 : OAI21_X1 port map( B1 => n4772, B2 => n12539, A => n2116, ZN => 
                           n4982);
   U5150 : OAI21_X1 port map( B1 => n2117, B2 => n2118, A => n12548, ZN => 
                           n2116);
   U5151 : NAND4_X1 port map( A1 => n2119, A2 => n2120, A3 => n2121, A4 => 
                           n2122, ZN => n2118);
   U5152 : NAND4_X1 port map( A1 => n2127, A2 => n2128, A3 => n2129, A4 => 
                           n2130, ZN => n2117);
   U5153 : OAI21_X1 port map( B1 => n4771, B2 => n12539, A => n2097, ZN => 
                           n4983);
   U5154 : OAI21_X1 port map( B1 => n2098, B2 => n2099, A => n12548, ZN => 
                           n2097);
   U5155 : NAND4_X1 port map( A1 => n2100, A2 => n2101, A3 => n2102, A4 => 
                           n2103, ZN => n2099);
   U5156 : NAND4_X1 port map( A1 => n2108, A2 => n2109, A3 => n2110, A4 => 
                           n2111, ZN => n2098);
   U5157 : OAI21_X1 port map( B1 => n4770, B2 => n12539, A => n2078, ZN => 
                           n4984);
   U5158 : OAI21_X1 port map( B1 => n2079, B2 => n2080, A => n12548, ZN => 
                           n2078);
   U5159 : NAND4_X1 port map( A1 => n2081, A2 => n2082, A3 => n2083, A4 => 
                           n2084, ZN => n2080);
   U5160 : NAND4_X1 port map( A1 => n2089, A2 => n2090, A3 => n2091, A4 => 
                           n2092, ZN => n2079);
   U5161 : OAI21_X1 port map( B1 => n4769, B2 => n12539, A => n2059, ZN => 
                           n4985);
   U5162 : OAI21_X1 port map( B1 => n2060, B2 => n2061, A => n12549, ZN => 
                           n2059);
   U5163 : NAND4_X1 port map( A1 => n2062, A2 => n2063, A3 => n2064, A4 => 
                           n2065, ZN => n2061);
   U5164 : NAND4_X1 port map( A1 => n2070, A2 => n2071, A3 => n2072, A4 => 
                           n2073, ZN => n2060);
   U5165 : OAI21_X1 port map( B1 => n4768, B2 => n12539, A => n2040, ZN => 
                           n4986);
   U5166 : OAI21_X1 port map( B1 => n2041, B2 => n2042, A => n12549, ZN => 
                           n2040);
   U5167 : NAND4_X1 port map( A1 => n2043, A2 => n2044, A3 => n2045, A4 => 
                           n2046, ZN => n2042);
   U5168 : NAND4_X1 port map( A1 => n2051, A2 => n2052, A3 => n2053, A4 => 
                           n2054, ZN => n2041);
   U5169 : OAI21_X1 port map( B1 => n4767, B2 => n12539, A => n2021, ZN => 
                           n4987);
   U5170 : OAI21_X1 port map( B1 => n2022, B2 => n2023, A => n12549, ZN => 
                           n2021);
   U5171 : NAND4_X1 port map( A1 => n2024, A2 => n2025, A3 => n2026, A4 => 
                           n2027, ZN => n2023);
   U5172 : NAND4_X1 port map( A1 => n2032, A2 => n2033, A3 => n2034, A4 => 
                           n2035, ZN => n2022);
   U5173 : OAI21_X1 port map( B1 => n4766, B2 => n12539, A => n2002, ZN => 
                           n4988);
   U5174 : OAI21_X1 port map( B1 => n2003, B2 => n2004, A => n12549, ZN => 
                           n2002);
   U5175 : NAND4_X1 port map( A1 => n2005, A2 => n2006, A3 => n2007, A4 => 
                           n2008, ZN => n2004);
   U5176 : NAND4_X1 port map( A1 => n2013, A2 => n2014, A3 => n2015, A4 => 
                           n2016, ZN => n2003);
   U5177 : OAI21_X1 port map( B1 => n4765, B2 => n12541, A => n1951, ZN => 
                           n4989);
   U5178 : OAI21_X1 port map( B1 => n1952, B2 => n1953, A => n12549, ZN => 
                           n1951);
   U5179 : NAND4_X1 port map( A1 => n1954, A2 => n1955, A3 => n1956, A4 => 
                           n1957, ZN => n1953);
   U5180 : NAND4_X1 port map( A1 => n1978, A2 => n1979, A3 => n1980, A4 => 
                           n1981, ZN => n1952);
   U5181 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n13387, 
                           ZN => n4465);
   U5182 : NOR3_X1 port map( A1 => n13387, A2 => ADD_RD2(3), A3 => n13391, ZN 
                           => n4466);
   U5183 : NOR2_X1 port map( A1 => n13390, A2 => ADD_RD2(2), ZN => n4452);
   U5184 : NOR3_X1 port map( A1 => n13387, A2 => ADD_RD2(0), A3 => n13388, ZN 
                           => n4469);
   U5185 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n13391, 
                           ZN => n4449);
   U5186 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n4451);
   U5187 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n13388, 
                           ZN => n4457);
   U5188 : NOR3_X1 port map( A1 => n13391, A2 => ADD_RD2(4), A3 => n13388, ZN 
                           => n4458);
   U5189 : AOI221_X1 port map( B1 => n12230, B2 => n4642, C1 => n12224, C2 => 
                           n4643, A => n4464, ZN => n4463);
   U5190 : OAI22_X1 port map( A1 => n8577, A2 => n12218, B1 => n8578, B2 => 
                           n12212, ZN => n4464);
   U5191 : AOI221_X1 port map( B1 => n12230, B2 => n4646, C1 => n12224, C2 => 
                           n4647, A => n4437, ZN => n4436);
   U5192 : OAI22_X1 port map( A1 => n8560, A2 => n12218, B1 => n8561, B2 => 
                           n12212, ZN => n4437);
   U5193 : AOI221_X1 port map( B1 => n12230, B2 => n4652, C1 => n12224, C2 => 
                           n4653, A => n4418, ZN => n4417);
   U5194 : OAI22_X1 port map( A1 => n8543, A2 => n12218, B1 => n8544, B2 => 
                           n12212, ZN => n4418);
   U5195 : AOI221_X1 port map( B1 => n12230, B2 => n4654, C1 => n12224, C2 => 
                           n4655, A => n4399, ZN => n4398);
   U5196 : OAI22_X1 port map( A1 => n8526, A2 => n12218, B1 => n8527, B2 => 
                           n12212, ZN => n4399);
   U5197 : AOI221_X1 port map( B1 => n12230, B2 => n8599, C1 => n12224, C2 => 
                           n8600, A => n4380, ZN => n4379);
   U5198 : OAI22_X1 port map( A1 => n8509, A2 => n12218, B1 => n8510, B2 => 
                           n12212, ZN => n4380);
   U5199 : AOI221_X1 port map( B1 => n12230, B2 => n8603, C1 => n12224, C2 => 
                           n8604, A => n4361, ZN => n4360);
   U5200 : OAI22_X1 port map( A1 => n8492, A2 => n12218, B1 => n8493, B2 => 
                           n12212, ZN => n4361);
   U5201 : AOI221_X1 port map( B1 => n12230, B2 => n8611, C1 => n12224, C2 => 
                           n8612, A => n4342, ZN => n4341);
   U5202 : OAI22_X1 port map( A1 => n8475, A2 => n12218, B1 => n8476, B2 => 
                           n12212, ZN => n4342);
   U5203 : AOI221_X1 port map( B1 => n12230, B2 => n8617, C1 => n12224, C2 => 
                           n8618, A => n4323, ZN => n4322);
   U5204 : OAI22_X1 port map( A1 => n8458, A2 => n12218, B1 => n8459, B2 => 
                           n12212, ZN => n4323);
   U5205 : AOI221_X1 port map( B1 => n12230, B2 => n8619, C1 => n12224, C2 => 
                           n8620, A => n4304, ZN => n4303);
   U5206 : OAI22_X1 port map( A1 => n8441, A2 => n12218, B1 => n8442, B2 => 
                           n12212, ZN => n4304);
   U5207 : AOI221_X1 port map( B1 => n12230, B2 => n8621, C1 => n12224, C2 => 
                           n8622, A => n4285, ZN => n4284);
   U5208 : OAI22_X1 port map( A1 => n8424, A2 => n12218, B1 => n8425, B2 => 
                           n12212, ZN => n4285);
   U5209 : AOI221_X1 port map( B1 => n12230, B2 => n8623, C1 => n12224, C2 => 
                           n8624, A => n4266, ZN => n4265);
   U5210 : OAI22_X1 port map( A1 => n8407, A2 => n12218, B1 => n8408, B2 => 
                           n12212, ZN => n4266);
   U5211 : AOI221_X1 port map( B1 => n12230, B2 => n8625, C1 => n12224, C2 => 
                           n8626, A => n4247, ZN => n4246);
   U5212 : OAI22_X1 port map( A1 => n8390, A2 => n12218, B1 => n8391, B2 => 
                           n12212, ZN => n4247);
   U5213 : AOI221_X1 port map( B1 => n12231, B2 => n8627, C1 => n12225, C2 => 
                           n8628, A => n4228, ZN => n4227);
   U5214 : OAI22_X1 port map( A1 => n8373, A2 => n12219, B1 => n8374, B2 => 
                           n12213, ZN => n4228);
   U5215 : AOI221_X1 port map( B1 => n12327, B2 => n9999, C1 => n12321, C2 => 
                           n9935, A => n4201, ZN => n4200);
   U5216 : OAI22_X1 port map( A1 => n14305, A2 => n12315, B1 => n13417, B2 => 
                           n12309, ZN => n4201);
   U5217 : AOI221_X1 port map( B1 => n12231, B2 => n8629, C1 => n12225, C2 => 
                           n8630, A => n4209, ZN => n4208);
   U5218 : OAI22_X1 port map( A1 => n8356, A2 => n12219, B1 => n8357, B2 => 
                           n12213, ZN => n4209);
   U5219 : AOI221_X1 port map( B1 => n12327, B2 => n9998, C1 => n12321, C2 => 
                           n9934, A => n4182, ZN => n4181);
   U5220 : OAI22_X1 port map( A1 => n14304, A2 => n12315, B1 => n13416, B2 => 
                           n12309, ZN => n4182);
   U5221 : AOI221_X1 port map( B1 => n12231, B2 => n8631, C1 => n12225, C2 => 
                           n8632, A => n4190, ZN => n4189);
   U5222 : OAI22_X1 port map( A1 => n8339, A2 => n12219, B1 => n8340, B2 => 
                           n12213, ZN => n4190);
   U5223 : AOI221_X1 port map( B1 => n12327, B2 => n9997, C1 => n12321, C2 => 
                           n9933, A => n4163, ZN => n4162);
   U5224 : OAI22_X1 port map( A1 => n14303, A2 => n12315, B1 => n13415, B2 => 
                           n12309, ZN => n4163);
   U5225 : AOI221_X1 port map( B1 => n12231, B2 => n8633, C1 => n12225, C2 => 
                           n8634, A => n4171, ZN => n4170);
   U5226 : OAI22_X1 port map( A1 => n8322, A2 => n12219, B1 => n8323, B2 => 
                           n12213, ZN => n4171);
   U5227 : AOI221_X1 port map( B1 => n12327, B2 => n9996, C1 => n12321, C2 => 
                           n9932, A => n4144, ZN => n4143);
   U5228 : OAI22_X1 port map( A1 => n14302, A2 => n12315, B1 => n13414, B2 => 
                           n12309, ZN => n4144);
   U5229 : AOI221_X1 port map( B1 => n12231, B2 => n8635, C1 => n12225, C2 => 
                           n8636, A => n4152, ZN => n4151);
   U5230 : OAI22_X1 port map( A1 => n8305, A2 => n12219, B1 => n8306, B2 => 
                           n12213, ZN => n4152);
   U5231 : AOI221_X1 port map( B1 => n12327, B2 => n9995, C1 => n12321, C2 => 
                           n9931, A => n4125, ZN => n4124);
   U5232 : OAI22_X1 port map( A1 => n14301, A2 => n12315, B1 => n13413, B2 => 
                           n12309, ZN => n4125);
   U5233 : AOI221_X1 port map( B1 => n12231, B2 => n8637, C1 => n12225, C2 => 
                           n8638, A => n4133, ZN => n4132);
   U5234 : OAI22_X1 port map( A1 => n8288, A2 => n12219, B1 => n8289, B2 => 
                           n12213, ZN => n4133);
   U5235 : AOI221_X1 port map( B1 => n12327, B2 => n9994, C1 => n12321, C2 => 
                           n9930, A => n4106, ZN => n4105);
   U5236 : OAI22_X1 port map( A1 => n14300, A2 => n12315, B1 => n13412, B2 => 
                           n12309, ZN => n4106);
   U5237 : AOI221_X1 port map( B1 => n12231, B2 => n8639, C1 => n12225, C2 => 
                           n8640, A => n4114, ZN => n4113);
   U5238 : OAI22_X1 port map( A1 => n8271, A2 => n12219, B1 => n8272, B2 => 
                           n12213, ZN => n4114);
   U5239 : AOI221_X1 port map( B1 => n12327, B2 => n9993, C1 => n12321, C2 => 
                           n9929, A => n4087, ZN => n4086);
   U5240 : OAI22_X1 port map( A1 => n14299, A2 => n12315, B1 => n13411, B2 => 
                           n12309, ZN => n4087);
   U5241 : AOI221_X1 port map( B1 => n12231, B2 => n8641, C1 => n12225, C2 => 
                           n8642, A => n4095, ZN => n4094);
   U5242 : OAI22_X1 port map( A1 => n8254, A2 => n12219, B1 => n8255, B2 => 
                           n12213, ZN => n4095);
   U5243 : AOI221_X1 port map( B1 => n12327, B2 => n9992, C1 => n12321, C2 => 
                           n9928, A => n4068, ZN => n4067);
   U5244 : OAI22_X1 port map( A1 => n14298, A2 => n12315, B1 => n13410, B2 => 
                           n12309, ZN => n4068);
   U5245 : AOI221_X1 port map( B1 => n12231, B2 => n8643, C1 => n12225, C2 => 
                           n8644, A => n4076, ZN => n4075);
   U5246 : OAI22_X1 port map( A1 => n8237, A2 => n12219, B1 => n8238, B2 => 
                           n12213, ZN => n4076);
   U5247 : AOI221_X1 port map( B1 => n12327, B2 => n9991, C1 => n12321, C2 => 
                           n9927, A => n4049, ZN => n4048);
   U5248 : OAI22_X1 port map( A1 => n14297, A2 => n12315, B1 => n13409, B2 => 
                           n12309, ZN => n4049);
   U5249 : AOI221_X1 port map( B1 => n12231, B2 => n8645, C1 => n12225, C2 => 
                           n8646, A => n4057, ZN => n4056);
   U5250 : OAI22_X1 port map( A1 => n8220, A2 => n12219, B1 => n8221, B2 => 
                           n12213, ZN => n4057);
   U5251 : AOI221_X1 port map( B1 => n12327, B2 => n9990, C1 => n12321, C2 => 
                           n9926, A => n4030, ZN => n4029);
   U5252 : OAI22_X1 port map( A1 => n14296, A2 => n12315, B1 => n13408, B2 => 
                           n12309, ZN => n4030);
   U5253 : AOI221_X1 port map( B1 => n12231, B2 => n8647, C1 => n12225, C2 => 
                           n8648, A => n4038, ZN => n4037);
   U5254 : OAI22_X1 port map( A1 => n8203, A2 => n12219, B1 => n8204, B2 => 
                           n12213, ZN => n4038);
   U5255 : AOI221_X1 port map( B1 => n12327, B2 => n9989, C1 => n12321, C2 => 
                           n9925, A => n4011, ZN => n4010);
   U5256 : OAI22_X1 port map( A1 => n14295, A2 => n12315, B1 => n13407, B2 => 
                           n12309, ZN => n4011);
   U5257 : AOI221_X1 port map( B1 => n12231, B2 => n8649, C1 => n12225, C2 => 
                           n8650, A => n4019, ZN => n4018);
   U5258 : OAI22_X1 port map( A1 => n8186, A2 => n12219, B1 => n8187, B2 => 
                           n12213, ZN => n4019);
   U5259 : AOI221_X1 port map( B1 => n12328, B2 => n9988, C1 => n12322, C2 => 
                           n9924, A => n3992, ZN => n3991);
   U5260 : OAI22_X1 port map( A1 => n14294, A2 => n12316, B1 => n13406, B2 => 
                           n12310, ZN => n3992);
   U5261 : AOI221_X1 port map( B1 => n12232, B2 => n8651, C1 => n12226, C2 => 
                           n8652, A => n4000, ZN => n3999);
   U5262 : OAI22_X1 port map( A1 => n8169, A2 => n12220, B1 => n8170, B2 => 
                           n12214, ZN => n4000);
   U5263 : AOI221_X1 port map( B1 => n12328, B2 => n9987, C1 => n12322, C2 => 
                           n9923, A => n3973, ZN => n3972);
   U5264 : OAI22_X1 port map( A1 => n14293, A2 => n12316, B1 => n13405, B2 => 
                           n12310, ZN => n3973);
   U5265 : AOI221_X1 port map( B1 => n12232, B2 => n8653, C1 => n12226, C2 => 
                           n8654, A => n3981, ZN => n3980);
   U5266 : OAI22_X1 port map( A1 => n8152, A2 => n12220, B1 => n8153, B2 => 
                           n12214, ZN => n3981);
   U5267 : AOI221_X1 port map( B1 => n12328, B2 => n9986, C1 => n12322, C2 => 
                           n9922, A => n3954, ZN => n3953);
   U5268 : OAI22_X1 port map( A1 => n14292, A2 => n12316, B1 => n13404, B2 => 
                           n12310, ZN => n3954);
   U5269 : AOI221_X1 port map( B1 => n12232, B2 => n8655, C1 => n12226, C2 => 
                           n8656, A => n3962, ZN => n3961);
   U5270 : OAI22_X1 port map( A1 => n8135, A2 => n12220, B1 => n8136, B2 => 
                           n12214, ZN => n3962);
   U5271 : AOI221_X1 port map( B1 => n12328, B2 => n9985, C1 => n12322, C2 => 
                           n9921, A => n3935, ZN => n3934);
   U5272 : OAI22_X1 port map( A1 => n14291, A2 => n12316, B1 => n13403, B2 => 
                           n12310, ZN => n3935);
   U5273 : AOI221_X1 port map( B1 => n12232, B2 => n8657, C1 => n12226, C2 => 
                           n8658, A => n3943, ZN => n3942);
   U5274 : OAI22_X1 port map( A1 => n8118, A2 => n12220, B1 => n8119, B2 => 
                           n12214, ZN => n3943);
   U5275 : AOI221_X1 port map( B1 => n12328, B2 => n9984, C1 => n12322, C2 => 
                           n9920, A => n3916, ZN => n3915);
   U5276 : OAI22_X1 port map( A1 => n14290, A2 => n12316, B1 => n13402, B2 => 
                           n12310, ZN => n3916);
   U5277 : AOI221_X1 port map( B1 => n12232, B2 => n8659, C1 => n12226, C2 => 
                           n8660, A => n3924, ZN => n3923);
   U5278 : OAI22_X1 port map( A1 => n8101, A2 => n12220, B1 => n8102, B2 => 
                           n12214, ZN => n3924);
   U5279 : AOI221_X1 port map( B1 => n12328, B2 => n9983, C1 => n12322, C2 => 
                           n9919, A => n3897, ZN => n3896);
   U5280 : OAI22_X1 port map( A1 => n14289, A2 => n12316, B1 => n14322, B2 => 
                           n12310, ZN => n3897);
   U5281 : AOI221_X1 port map( B1 => n12232, B2 => n8661, C1 => n12226, C2 => 
                           n8662, A => n3905, ZN => n3904);
   U5282 : OAI22_X1 port map( A1 => n8084, A2 => n12220, B1 => n8085, B2 => 
                           n12214, ZN => n3905);
   U5283 : AOI221_X1 port map( B1 => n12328, B2 => n9982, C1 => n12322, C2 => 
                           n9918, A => n3878, ZN => n3877);
   U5284 : OAI22_X1 port map( A1 => n14456, A2 => n12316, B1 => n14321, B2 => 
                           n12310, ZN => n3878);
   U5285 : AOI221_X1 port map( B1 => n12232, B2 => n8663, C1 => n12226, C2 => 
                           n8664, A => n3886, ZN => n3885);
   U5286 : OAI22_X1 port map( A1 => n8067, A2 => n12220, B1 => n8068, B2 => 
                           n12214, ZN => n3886);
   U5287 : AOI221_X1 port map( B1 => n12328, B2 => n9981, C1 => n12322, C2 => 
                           n9917, A => n3859, ZN => n3858);
   U5288 : OAI22_X1 port map( A1 => n14455, A2 => n12316, B1 => n14320, B2 => 
                           n12310, ZN => n3859);
   U5289 : AOI221_X1 port map( B1 => n12232, B2 => n8665, C1 => n12226, C2 => 
                           n8666, A => n3867, ZN => n3866);
   U5290 : OAI22_X1 port map( A1 => n8050, A2 => n12220, B1 => n8051, B2 => 
                           n12214, ZN => n3867);
   U5291 : AOI221_X1 port map( B1 => n12328, B2 => n9980, C1 => n12322, C2 => 
                           n9916, A => n3840, ZN => n3839);
   U5292 : OAI22_X1 port map( A1 => n14454, A2 => n12316, B1 => n14319, B2 => 
                           n12310, ZN => n3840);
   U5293 : AOI221_X1 port map( B1 => n12232, B2 => n8667, C1 => n12226, C2 => 
                           n8668, A => n3848, ZN => n3847);
   U5294 : OAI22_X1 port map( A1 => n8033, A2 => n12220, B1 => n8034, B2 => 
                           n12214, ZN => n3848);
   U5295 : AOI221_X1 port map( B1 => n12328, B2 => n9979, C1 => n12322, C2 => 
                           n9915, A => n3821, ZN => n3820);
   U5296 : OAI22_X1 port map( A1 => n14453, A2 => n12316, B1 => n14318, B2 => 
                           n12310, ZN => n3821);
   U5297 : AOI221_X1 port map( B1 => n12232, B2 => n8669, C1 => n12226, C2 => 
                           n8670, A => n3829, ZN => n3828);
   U5298 : OAI22_X1 port map( A1 => n8016, A2 => n12220, B1 => n8017, B2 => 
                           n12214, ZN => n3829);
   U5299 : AOI221_X1 port map( B1 => n12328, B2 => n9978, C1 => n12322, C2 => 
                           n9914, A => n3802, ZN => n3801);
   U5300 : OAI22_X1 port map( A1 => n14452, A2 => n12316, B1 => n14317, B2 => 
                           n12310, ZN => n3802);
   U5301 : AOI221_X1 port map( B1 => n12232, B2 => n8671, C1 => n12226, C2 => 
                           n8672, A => n3810, ZN => n3809);
   U5302 : OAI22_X1 port map( A1 => n7999, A2 => n12220, B1 => n8000, B2 => 
                           n12214, ZN => n3810);
   U5303 : AOI221_X1 port map( B1 => n12328, B2 => n9977, C1 => n12322, C2 => 
                           n9913, A => n3783, ZN => n3782);
   U5304 : OAI22_X1 port map( A1 => n14451, A2 => n12316, B1 => n14316, B2 => 
                           n12310, ZN => n3783);
   U5305 : AOI221_X1 port map( B1 => n12232, B2 => n8673, C1 => n12226, C2 => 
                           n8674, A => n3791, ZN => n3790);
   U5306 : OAI22_X1 port map( A1 => n7982, A2 => n12220, B1 => n7983, B2 => 
                           n12214, ZN => n3791);
   U5307 : AOI221_X1 port map( B1 => n12329, B2 => n9976, C1 => n12323, C2 => 
                           n9912, A => n3764, ZN => n3763);
   U5308 : OAI22_X1 port map( A1 => n14450, A2 => n12317, B1 => n14315, B2 => 
                           n12311, ZN => n3764);
   U5309 : AOI221_X1 port map( B1 => n12233, B2 => n8675, C1 => n12227, C2 => 
                           n8676, A => n3772, ZN => n3771);
   U5310 : OAI22_X1 port map( A1 => n7965, A2 => n12221, B1 => n7966, B2 => 
                           n12215, ZN => n3772);
   U5311 : AOI221_X1 port map( B1 => n12329, B2 => n9975, C1 => n12323, C2 => 
                           n9911, A => n3745, ZN => n3744);
   U5312 : OAI22_X1 port map( A1 => n14449, A2 => n12317, B1 => n14314, B2 => 
                           n12311, ZN => n3745);
   U5313 : AOI221_X1 port map( B1 => n12233, B2 => n8677, C1 => n12227, C2 => 
                           n8678, A => n3753, ZN => n3752);
   U5314 : OAI22_X1 port map( A1 => n7948, A2 => n12221, B1 => n7949, B2 => 
                           n12215, ZN => n3753);
   U5315 : AOI221_X1 port map( B1 => n12329, B2 => n9974, C1 => n12323, C2 => 
                           n9910, A => n3726, ZN => n3725);
   U5316 : OAI22_X1 port map( A1 => n14448, A2 => n12317, B1 => n14313, B2 => 
                           n12311, ZN => n3726);
   U5317 : AOI221_X1 port map( B1 => n12233, B2 => n8679, C1 => n12227, C2 => 
                           n8680, A => n3734, ZN => n3733);
   U5318 : OAI22_X1 port map( A1 => n7931, A2 => n12221, B1 => n7932, B2 => 
                           n12215, ZN => n3734);
   U5319 : AOI221_X1 port map( B1 => n12329, B2 => n9973, C1 => n12323, C2 => 
                           n9909, A => n3707, ZN => n3706);
   U5320 : OAI22_X1 port map( A1 => n14447, A2 => n12317, B1 => n14312, B2 => 
                           n12311, ZN => n3707);
   U5321 : AOI221_X1 port map( B1 => n12233, B2 => n8681, C1 => n12227, C2 => 
                           n8682, A => n3715, ZN => n3714);
   U5322 : OAI22_X1 port map( A1 => n7914, A2 => n12221, B1 => n7915, B2 => 
                           n12215, ZN => n3715);
   U5323 : AOI221_X1 port map( B1 => n12329, B2 => n9972, C1 => n12323, C2 => 
                           n9908, A => n3688, ZN => n3687);
   U5324 : OAI22_X1 port map( A1 => n14446, A2 => n12317, B1 => n14432, B2 => 
                           n12311, ZN => n3688);
   U5325 : AOI221_X1 port map( B1 => n12233, B2 => n8683, C1 => n12227, C2 => 
                           n8684, A => n3696, ZN => n3695);
   U5326 : OAI22_X1 port map( A1 => n7897, A2 => n12221, B1 => n7898, B2 => 
                           n12215, ZN => n3696);
   U5327 : AOI221_X1 port map( B1 => n12329, B2 => n9971, C1 => n12323, C2 => 
                           n9907, A => n3669, ZN => n3668);
   U5328 : OAI22_X1 port map( A1 => n14445, A2 => n12317, B1 => n14431, B2 => 
                           n12311, ZN => n3669);
   U5329 : AOI221_X1 port map( B1 => n12233, B2 => n8685, C1 => n12227, C2 => 
                           n8686, A => n3677, ZN => n3676);
   U5330 : OAI22_X1 port map( A1 => n7880, A2 => n12221, B1 => n7881, B2 => 
                           n12215, ZN => n3677);
   U5331 : AOI221_X1 port map( B1 => n12329, B2 => n9970, C1 => n12323, C2 => 
                           n9906, A => n3650, ZN => n3649);
   U5332 : OAI22_X1 port map( A1 => n14444, A2 => n12317, B1 => n14430, B2 => 
                           n12311, ZN => n3650);
   U5333 : AOI221_X1 port map( B1 => n12233, B2 => n8687, C1 => n12227, C2 => 
                           n8688, A => n3658, ZN => n3657);
   U5334 : OAI22_X1 port map( A1 => n7863, A2 => n12221, B1 => n7864, B2 => 
                           n12215, ZN => n3658);
   U5335 : AOI221_X1 port map( B1 => n12329, B2 => n9969, C1 => n12323, C2 => 
                           n9905, A => n3631, ZN => n3630);
   U5336 : OAI22_X1 port map( A1 => n14443, A2 => n12317, B1 => n14429, B2 => 
                           n12311, ZN => n3631);
   U5337 : AOI221_X1 port map( B1 => n12233, B2 => n8689, C1 => n12227, C2 => 
                           n8690, A => n3639, ZN => n3638);
   U5338 : OAI22_X1 port map( A1 => n7846, A2 => n12221, B1 => n7847, B2 => 
                           n12215, ZN => n3639);
   U5339 : AOI221_X1 port map( B1 => n12329, B2 => n9968, C1 => n12323, C2 => 
                           n9904, A => n3612, ZN => n3611);
   U5340 : OAI22_X1 port map( A1 => n14442, A2 => n12317, B1 => n14428, B2 => 
                           n12311, ZN => n3612);
   U5341 : AOI221_X1 port map( B1 => n12233, B2 => n8691, C1 => n12227, C2 => 
                           n8692, A => n3620, ZN => n3619);
   U5342 : OAI22_X1 port map( A1 => n7829, A2 => n12221, B1 => n7830, B2 => 
                           n12215, ZN => n3620);
   U5343 : AOI221_X1 port map( B1 => n12329, B2 => n9967, C1 => n12323, C2 => 
                           n9903, A => n3593, ZN => n3592);
   U5344 : OAI22_X1 port map( A1 => n14441, A2 => n12317, B1 => n14427, B2 => 
                           n12311, ZN => n3593);
   U5345 : AOI221_X1 port map( B1 => n12233, B2 => n8693, C1 => n12227, C2 => 
                           n8694, A => n3601, ZN => n3600);
   U5346 : OAI22_X1 port map( A1 => n7812, A2 => n12221, B1 => n7813, B2 => 
                           n12215, ZN => n3601);
   U5347 : AOI221_X1 port map( B1 => n12329, B2 => n9966, C1 => n12323, C2 => 
                           n9902, A => n3574, ZN => n3573);
   U5348 : OAI22_X1 port map( A1 => n13401, A2 => n12317, B1 => n14426, B2 => 
                           n12311, ZN => n3574);
   U5349 : AOI221_X1 port map( B1 => n12233, B2 => n8695, C1 => n12227, C2 => 
                           n8696, A => n3582, ZN => n3581);
   U5350 : OAI22_X1 port map( A1 => n7795, A2 => n12221, B1 => n7796, B2 => 
                           n12215, ZN => n3582);
   U5351 : AOI221_X1 port map( B1 => n12329, B2 => n9965, C1 => n12323, C2 => 
                           n9901, A => n3555, ZN => n3554);
   U5352 : OAI22_X1 port map( A1 => n13400, A2 => n12317, B1 => n14425, B2 => 
                           n12311, ZN => n3555);
   U5353 : AOI221_X1 port map( B1 => n12233, B2 => n4656, C1 => n12227, C2 => 
                           n4657, A => n3563, ZN => n3562);
   U5354 : OAI22_X1 port map( A1 => n7778, A2 => n12221, B1 => n7779, B2 => 
                           n12215, ZN => n3563);
   U5355 : AOI221_X1 port map( B1 => n12330, B2 => n9964, C1 => n12324, C2 => 
                           n9900, A => n3536, ZN => n3535);
   U5356 : OAI22_X1 port map( A1 => n13399, A2 => n12318, B1 => n14424, B2 => 
                           n12312, ZN => n3536);
   U5357 : AOI221_X1 port map( B1 => n12234, B2 => n4658, C1 => n12228, C2 => 
                           n4659, A => n3544, ZN => n3543);
   U5358 : OAI22_X1 port map( A1 => n7761, A2 => n12222, B1 => n7762, B2 => 
                           n12216, ZN => n3544);
   U5359 : AOI221_X1 port map( B1 => n12330, B2 => n9963, C1 => n12324, C2 => 
                           n9899, A => n3517, ZN => n3516);
   U5360 : OAI22_X1 port map( A1 => n13398, A2 => n12318, B1 => n14423, B2 => 
                           n12312, ZN => n3517);
   U5361 : AOI221_X1 port map( B1 => n12234, B2 => n4660, C1 => n12228, C2 => 
                           n4661, A => n3525, ZN => n3524);
   U5362 : OAI22_X1 port map( A1 => n7744, A2 => n12222, B1 => n7745, B2 => 
                           n12216, ZN => n3525);
   U5363 : AOI221_X1 port map( B1 => n12330, B2 => n9962, C1 => n12324, C2 => 
                           n9898, A => n3498, ZN => n3497);
   U5364 : OAI22_X1 port map( A1 => n13397, A2 => n12318, B1 => n14422, B2 => 
                           n12312, ZN => n3498);
   U5365 : AOI221_X1 port map( B1 => n12234, B2 => n4662, C1 => n12228, C2 => 
                           n4663, A => n3506, ZN => n3505);
   U5366 : OAI22_X1 port map( A1 => n7642, A2 => n12222, B1 => n7643, B2 => 
                           n12216, ZN => n3506);
   U5367 : AOI221_X1 port map( B1 => n12330, B2 => n9961, C1 => n12324, C2 => 
                           n9897, A => n3479, ZN => n3478);
   U5368 : OAI22_X1 port map( A1 => n13396, A2 => n12318, B1 => n14421, B2 => 
                           n12312, ZN => n3479);
   U5369 : AOI221_X1 port map( B1 => n12234, B2 => n4664, C1 => n12228, C2 => 
                           n4665, A => n3487, ZN => n3486);
   U5370 : OAI22_X1 port map( A1 => n7625, A2 => n12222, B1 => n7626, B2 => 
                           n12216, ZN => n3487);
   U5371 : AOI221_X1 port map( B1 => n12330, B2 => n9960, C1 => n12324, C2 => 
                           n9896, A => n3460, ZN => n3459);
   U5372 : OAI22_X1 port map( A1 => n13395, A2 => n12318, B1 => n14420, B2 => 
                           n12312, ZN => n3460);
   U5373 : AOI221_X1 port map( B1 => n12234, B2 => n4666, C1 => n12228, C2 => 
                           n4667, A => n3468, ZN => n3467);
   U5374 : OAI22_X1 port map( A1 => n7521, A2 => n12222, B1 => n7522, B2 => 
                           n12216, ZN => n3468);
   U5375 : AOI221_X1 port map( B1 => n12330, B2 => n9959, C1 => n12324, C2 => 
                           n9895, A => n3441, ZN => n3440);
   U5376 : OAI22_X1 port map( A1 => n13394, A2 => n12318, B1 => n14419, B2 => 
                           n12312, ZN => n3441);
   U5377 : AOI221_X1 port map( B1 => n12234, B2 => n4668, C1 => n12228, C2 => 
                           n4669, A => n3449, ZN => n3448);
   U5378 : OAI22_X1 port map( A1 => n7504, A2 => n12222, B1 => n7505, B2 => 
                           n12216, ZN => n3449);
   U5379 : AOI221_X1 port map( B1 => n12330, B2 => n9958, C1 => n12324, C2 => 
                           n9894, A => n3422, ZN => n3421);
   U5380 : OAI22_X1 port map( A1 => n13393, A2 => n12318, B1 => n14418, B2 => 
                           n12312, ZN => n3422);
   U5381 : AOI221_X1 port map( B1 => n12234, B2 => n4670, C1 => n12228, C2 => 
                           n4671, A => n3430, ZN => n3429);
   U5382 : OAI22_X1 port map( A1 => n7402, A2 => n12222, B1 => n7403, B2 => 
                           n12216, ZN => n3430);
   U5383 : AOI221_X1 port map( B1 => n12330, B2 => n9957, C1 => n12324, C2 => 
                           n9893, A => n3403, ZN => n3402);
   U5384 : OAI22_X1 port map( A1 => n14440, A2 => n12318, B1 => n14417, B2 => 
                           n12312, ZN => n3403);
   U5385 : AOI221_X1 port map( B1 => n12234, B2 => n4672, C1 => n12228, C2 => 
                           n4673, A => n3411, ZN => n3410);
   U5386 : OAI22_X1 port map( A1 => n7385, A2 => n12222, B1 => n7386, B2 => 
                           n12216, ZN => n3411);
   U5387 : AOI221_X1 port map( B1 => n12330, B2 => n9956, C1 => n12324, C2 => 
                           n9892, A => n3384, ZN => n3383);
   U5388 : OAI22_X1 port map( A1 => n14439, A2 => n12318, B1 => n14416, B2 => 
                           n12312, ZN => n3384);
   U5389 : AOI221_X1 port map( B1 => n12234, B2 => n4674, C1 => n12228, C2 => 
                           n4675, A => n3392, ZN => n3391);
   U5390 : OAI22_X1 port map( A1 => n7368, A2 => n12222, B1 => n7369, B2 => 
                           n12216, ZN => n3392);
   U5391 : AOI221_X1 port map( B1 => n12330, B2 => n9955, C1 => n12324, C2 => 
                           n9891, A => n3365, ZN => n3364);
   U5392 : OAI22_X1 port map( A1 => n14438, A2 => n12318, B1 => n14415, B2 => 
                           n12312, ZN => n3365);
   U5393 : AOI221_X1 port map( B1 => n12234, B2 => n4676, C1 => n12228, C2 => 
                           n4677, A => n3373, ZN => n3372);
   U5394 : OAI22_X1 port map( A1 => n7269, A2 => n12222, B1 => n7270, B2 => 
                           n12216, ZN => n3373);
   U5395 : AOI221_X1 port map( B1 => n12330, B2 => n9954, C1 => n12324, C2 => 
                           n9890, A => n3346, ZN => n3345);
   U5396 : OAI22_X1 port map( A1 => n14437, A2 => n12318, B1 => n14414, B2 => 
                           n12312, ZN => n3346);
   U5397 : AOI221_X1 port map( B1 => n12234, B2 => n4678, C1 => n12228, C2 => 
                           n4679, A => n3354, ZN => n3353);
   U5398 : OAI22_X1 port map( A1 => n7252, A2 => n12222, B1 => n7253, B2 => 
                           n12216, ZN => n3354);
   U5399 : AOI221_X1 port map( B1 => n12330, B2 => n9953, C1 => n12324, C2 => 
                           n9889, A => n3327, ZN => n3326);
   U5400 : OAI22_X1 port map( A1 => n14436, A2 => n12318, B1 => n14413, B2 => 
                           n12312, ZN => n3327);
   U5401 : AOI221_X1 port map( B1 => n12234, B2 => n4682, C1 => n12228, C2 => 
                           n4683, A => n3335, ZN => n3334);
   U5402 : OAI22_X1 port map( A1 => n7235, A2 => n12222, B1 => n7236, B2 => 
                           n12216, ZN => n3335);
   U5403 : AOI221_X1 port map( B1 => n12235, B2 => n4472, C1 => n12229, C2 => 
                           n4473, A => n3316, ZN => n3315);
   U5404 : OAI22_X1 port map( A1 => n7138, A2 => n12223, B1 => n7139, B2 => 
                           n12217, ZN => n3316);
   U5405 : AOI221_X1 port map( B1 => n12331, B2 => n9952, C1 => n12325, C2 => 
                           n9888, A => n3308, ZN => n3307);
   U5406 : OAI22_X1 port map( A1 => n14435, A2 => n12319, B1 => n14412, B2 => 
                           n12313, ZN => n3308);
   U5407 : AOI221_X1 port map( B1 => n12235, B2 => n4474, C1 => n12229, C2 => 
                           n4475, A => n3297, ZN => n3296);
   U5408 : OAI22_X1 port map( A1 => n7121, A2 => n12223, B1 => n7122, B2 => 
                           n12217, ZN => n3297);
   U5409 : AOI221_X1 port map( B1 => n12331, B2 => n9951, C1 => n12325, C2 => 
                           n9887, A => n3289, ZN => n3288);
   U5410 : OAI22_X1 port map( A1 => n14434, A2 => n12319, B1 => n14411, B2 => 
                           n12313, ZN => n3289);
   U5411 : AOI221_X1 port map( B1 => n12235, B2 => n4476, C1 => n12229, C2 => 
                           n4477, A => n3278, ZN => n3277);
   U5412 : OAI22_X1 port map( A1 => n4860, A2 => n12223, B1 => n4861, B2 => 
                           n12217, ZN => n3278);
   U5413 : AOI221_X1 port map( B1 => n12331, B2 => n9950, C1 => n12325, C2 => 
                           n9886, A => n3270, ZN => n3269);
   U5414 : OAI22_X1 port map( A1 => n14433, A2 => n12319, B1 => n14410, B2 => 
                           n12313, ZN => n3270);
   U5415 : AOI221_X1 port map( B1 => n12235, B2 => n4478, C1 => n12229, C2 => 
                           n4479, A => n3245, ZN => n3242);
   U5416 : OAI22_X1 port map( A1 => n4843, A2 => n12223, B1 => n4844, B2 => 
                           n12217, ZN => n3245);
   U5417 : AOI221_X1 port map( B1 => n12331, B2 => n9949, C1 => n12325, C2 => 
                           n9885, A => n3221, ZN => n3218);
   U5418 : OAI22_X1 port map( A1 => n13392, A2 => n12319, B1 => n14409, B2 => 
                           n12313, ZN => n3221);
   U5419 : AOI221_X1 port map( B1 => n12326, B2 => n11766, C1 => n12320, C2 => 
                           n9948, A => n4448, ZN => n4447);
   U5420 : OAI22_X1 port map( A1 => n14216, A2 => n12314, B1 => n13430, B2 => 
                           n12308, ZN => n4448);
   U5421 : AOI221_X1 port map( B1 => n12326, B2 => n11767, C1 => n12320, C2 => 
                           n9947, A => n4429, ZN => n4428);
   U5422 : OAI22_X1 port map( A1 => n14328, A2 => n12314, B1 => n13429, B2 => 
                           n12308, ZN => n4429);
   U5423 : AOI221_X1 port map( B1 => n12326, B2 => n11768, C1 => n12320, C2 => 
                           n9946, A => n4410, ZN => n4409);
   U5424 : OAI22_X1 port map( A1 => n14327, A2 => n12314, B1 => n13428, B2 => 
                           n12308, ZN => n4410);
   U5425 : AOI221_X1 port map( B1 => n12326, B2 => n11769, C1 => n12320, C2 => 
                           n9945, A => n4391, ZN => n4390);
   U5426 : OAI22_X1 port map( A1 => n14326, A2 => n12314, B1 => n13427, B2 => 
                           n12308, ZN => n4391);
   U5427 : AOI221_X1 port map( B1 => n12326, B2 => n11770, C1 => n12320, C2 => 
                           n9944, A => n4372, ZN => n4371);
   U5428 : OAI22_X1 port map( A1 => n14325, A2 => n12314, B1 => n13426, B2 => 
                           n12308, ZN => n4372);
   U5429 : AOI221_X1 port map( B1 => n12326, B2 => n11771, C1 => n12320, C2 => 
                           n9943, A => n4353, ZN => n4352);
   U5430 : OAI22_X1 port map( A1 => n14324, A2 => n12314, B1 => n13425, B2 => 
                           n12308, ZN => n4353);
   U5431 : AOI221_X1 port map( B1 => n12326, B2 => n11772, C1 => n12320, C2 => 
                           n9942, A => n4334, ZN => n4333);
   U5432 : OAI22_X1 port map( A1 => n14311, A2 => n12314, B1 => n13424, B2 => 
                           n12308, ZN => n4334);
   U5433 : AOI221_X1 port map( B1 => n12326, B2 => n11773, C1 => n12320, C2 => 
                           n9941, A => n4315, ZN => n4314);
   U5434 : OAI22_X1 port map( A1 => n14310, A2 => n12314, B1 => n13423, B2 => 
                           n12308, ZN => n4315);
   U5435 : AOI221_X1 port map( B1 => n12326, B2 => n11774, C1 => n12320, C2 => 
                           n9940, A => n4296, ZN => n4295);
   U5436 : OAI22_X1 port map( A1 => n14323, A2 => n12314, B1 => n13422, B2 => 
                           n12308, ZN => n4296);
   U5437 : AOI221_X1 port map( B1 => n12326, B2 => n11775, C1 => n12320, C2 => 
                           n9939, A => n4277, ZN => n4276);
   U5438 : OAI22_X1 port map( A1 => n14309, A2 => n12314, B1 => n13421, B2 => 
                           n12308, ZN => n4277);
   U5439 : AOI221_X1 port map( B1 => n12326, B2 => n11776, C1 => n12320, C2 => 
                           n9938, A => n4258, ZN => n4257);
   U5440 : OAI22_X1 port map( A1 => n14308, A2 => n12314, B1 => n13420, B2 => 
                           n12308, ZN => n4258);
   U5441 : AOI221_X1 port map( B1 => n12326, B2 => n11777, C1 => n12320, C2 => 
                           n9937, A => n4239, ZN => n4238);
   U5442 : OAI22_X1 port map( A1 => n14307, A2 => n12314, B1 => n13419, B2 => 
                           n12308, ZN => n4239);
   U5443 : AOI221_X1 port map( B1 => n12327, B2 => n11778, C1 => n12321, C2 => 
                           n9936, A => n4220, ZN => n4219);
   U5444 : OAI22_X1 port map( A1 => n14306, A2 => n12315, B1 => n13418, B2 => 
                           n12309, ZN => n4220);
   U5445 : AOI221_X1 port map( B1 => n12206, B2 => n4480, C1 => n12200, C2 => 
                           n4481, A => n4467, ZN => n4462);
   U5446 : OAI22_X1 port map( A1 => n8579, A2 => n12194, B1 => n8580, B2 => 
                           n12188, ZN => n4467);
   U5447 : AOI221_X1 port map( B1 => n12206, B2 => n4648, C1 => n12200, C2 => 
                           n4649, A => n4438, ZN => n4435);
   U5448 : OAI22_X1 port map( A1 => n8562, A2 => n12194, B1 => n8563, B2 => 
                           n12188, ZN => n4438);
   U5449 : AOI221_X1 port map( B1 => n12206, B2 => n4482, C1 => n12200, C2 => 
                           n4483, A => n4419, ZN => n4416);
   U5450 : OAI22_X1 port map( A1 => n8545, A2 => n12194, B1 => n8546, B2 => 
                           n12188, ZN => n4419);
   U5451 : AOI221_X1 port map( B1 => n12206, B2 => n4484, C1 => n12200, C2 => 
                           n4485, A => n4400, ZN => n4397);
   U5452 : OAI22_X1 port map( A1 => n8528, A2 => n12194, B1 => n8529, B2 => 
                           n12188, ZN => n4400);
   U5453 : AOI221_X1 port map( B1 => n12206, B2 => n7080, C1 => n12200, C2 => 
                           n7081, A => n4381, ZN => n4378);
   U5454 : OAI22_X1 port map( A1 => n8511, A2 => n12194, B1 => n8512, B2 => 
                           n12188, ZN => n4381);
   U5455 : AOI221_X1 port map( B1 => n12206, B2 => n8605, C1 => n12200, C2 => 
                           n8606, A => n4362, ZN => n4359);
   U5456 : OAI22_X1 port map( A1 => n8494, A2 => n12194, B1 => n8495, B2 => 
                           n12188, ZN => n4362);
   U5457 : AOI221_X1 port map( B1 => n12206, B2 => n8613, C1 => n12200, C2 => 
                           n8614, A => n4343, ZN => n4340);
   U5458 : OAI22_X1 port map( A1 => n8477, A2 => n12194, B1 => n8478, B2 => 
                           n12188, ZN => n4343);
   U5459 : AOI221_X1 port map( B1 => n12206, B2 => n7084, C1 => n12200, C2 => 
                           n7085, A => n4324, ZN => n4321);
   U5460 : OAI22_X1 port map( A1 => n8460, A2 => n12194, B1 => n8461, B2 => 
                           n12188, ZN => n4324);
   U5461 : AOI221_X1 port map( B1 => n12206, B2 => n7088, C1 => n12200, C2 => 
                           n7089, A => n4305, ZN => n4302);
   U5462 : OAI22_X1 port map( A1 => n8443, A2 => n12194, B1 => n8444, B2 => 
                           n12188, ZN => n4305);
   U5463 : AOI221_X1 port map( B1 => n12206, B2 => n7092, C1 => n12200, C2 => 
                           n7093, A => n4286, ZN => n4283);
   U5464 : OAI22_X1 port map( A1 => n8426, A2 => n12194, B1 => n8427, B2 => 
                           n12188, ZN => n4286);
   U5465 : AOI221_X1 port map( B1 => n12206, B2 => n7096, C1 => n12200, C2 => 
                           n7097, A => n4267, ZN => n4264);
   U5466 : OAI22_X1 port map( A1 => n8409, A2 => n12194, B1 => n8410, B2 => 
                           n12188, ZN => n4267);
   U5467 : AOI221_X1 port map( B1 => n12206, B2 => n7100, C1 => n12200, C2 => 
                           n7101, A => n4248, ZN => n4245);
   U5468 : OAI22_X1 port map( A1 => n8392, A2 => n12194, B1 => n8393, B2 => 
                           n12188, ZN => n4248);
   U5469 : AOI221_X1 port map( B1 => n12207, B2 => n7104, C1 => n12201, C2 => 
                           n7105, A => n4229, ZN => n4226);
   U5470 : OAI22_X1 port map( A1 => n8375, A2 => n12195, B1 => n8376, B2 => 
                           n12189, ZN => n4229);
   U5471 : AOI221_X1 port map( B1 => n12207, B2 => n7130, C1 => n12201, C2 => 
                           n7131, A => n4210, ZN => n4207);
   U5472 : OAI22_X1 port map( A1 => n8358, A2 => n12195, B1 => n8359, B2 => 
                           n12189, ZN => n4210);
   U5473 : AOI221_X1 port map( B1 => n12207, B2 => n7154, C1 => n12201, C2 => 
                           n7155, A => n4191, ZN => n4188);
   U5474 : OAI22_X1 port map( A1 => n8341, A2 => n12195, B1 => n8342, B2 => 
                           n12189, ZN => n4191);
   U5475 : AOI221_X1 port map( B1 => n12207, B2 => n7158, C1 => n12201, C2 => 
                           n7159, A => n4172, ZN => n4169);
   U5476 : OAI22_X1 port map( A1 => n8324, A2 => n12195, B1 => n8325, B2 => 
                           n12189, ZN => n4172);
   U5477 : AOI221_X1 port map( B1 => n12207, B2 => n7162, C1 => n12201, C2 => 
                           n7163, A => n4153, ZN => n4150);
   U5478 : OAI22_X1 port map( A1 => n8307, A2 => n12195, B1 => n8308, B2 => 
                           n12189, ZN => n4153);
   U5479 : AOI221_X1 port map( B1 => n12207, B2 => n7166, C1 => n12201, C2 => 
                           n7167, A => n4134, ZN => n4131);
   U5480 : OAI22_X1 port map( A1 => n8290, A2 => n12195, B1 => n8291, B2 => 
                           n12189, ZN => n4134);
   U5481 : AOI221_X1 port map( B1 => n12207, B2 => n7170, C1 => n12201, C2 => 
                           n7171, A => n4115, ZN => n4112);
   U5482 : OAI22_X1 port map( A1 => n8273, A2 => n12195, B1 => n8274, B2 => 
                           n12189, ZN => n4115);
   U5483 : AOI221_X1 port map( B1 => n12207, B2 => n7174, C1 => n12201, C2 => 
                           n7175, A => n4096, ZN => n4093);
   U5484 : OAI22_X1 port map( A1 => n8256, A2 => n12195, B1 => n8257, B2 => 
                           n12189, ZN => n4096);
   U5485 : AOI221_X1 port map( B1 => n12207, B2 => n7178, C1 => n12201, C2 => 
                           n7179, A => n4077, ZN => n4074);
   U5486 : OAI22_X1 port map( A1 => n8239, A2 => n12195, B1 => n8240, B2 => 
                           n12189, ZN => n4077);
   U5487 : AOI221_X1 port map( B1 => n12207, B2 => n7182, C1 => n12201, C2 => 
                           n7183, A => n4058, ZN => n4055);
   U5488 : OAI22_X1 port map( A1 => n8222, A2 => n12195, B1 => n8223, B2 => 
                           n12189, ZN => n4058);
   U5489 : AOI221_X1 port map( B1 => n12207, B2 => n7186, C1 => n12201, C2 => 
                           n7187, A => n4039, ZN => n4036);
   U5490 : OAI22_X1 port map( A1 => n8205, A2 => n12195, B1 => n8206, B2 => 
                           n12189, ZN => n4039);
   U5491 : AOI221_X1 port map( B1 => n12207, B2 => n7190, C1 => n12201, C2 => 
                           n7191, A => n4020, ZN => n4017);
   U5492 : OAI22_X1 port map( A1 => n8188, A2 => n12195, B1 => n8189, B2 => 
                           n12189, ZN => n4020);
   U5493 : AOI221_X1 port map( B1 => n12208, B2 => n7194, C1 => n12202, C2 => 
                           n7195, A => n4001, ZN => n3998);
   U5494 : OAI22_X1 port map( A1 => n8171, A2 => n12196, B1 => n8172, B2 => 
                           n12190, ZN => n4001);
   U5495 : AOI221_X1 port map( B1 => n12208, B2 => n7198, C1 => n12202, C2 => 
                           n7199, A => n3982, ZN => n3979);
   U5496 : OAI22_X1 port map( A1 => n8154, A2 => n12196, B1 => n8155, B2 => 
                           n12190, ZN => n3982);
   U5497 : AOI221_X1 port map( B1 => n12208, B2 => n7202, C1 => n12202, C2 => 
                           n8708, A => n3963, ZN => n3960);
   U5498 : OAI22_X1 port map( A1 => n8137, A2 => n12196, B1 => n8138, B2 => 
                           n12190, ZN => n3963);
   U5499 : AOI221_X1 port map( B1 => n12208, B2 => n7205, C1 => n12202, C2 => 
                           n8707, A => n3944, ZN => n3941);
   U5500 : OAI22_X1 port map( A1 => n8120, A2 => n12196, B1 => n8121, B2 => 
                           n12190, ZN => n3944);
   U5501 : AOI221_X1 port map( B1 => n12208, B2 => n7208, C1 => n12202, C2 => 
                           n8706, A => n3925, ZN => n3922);
   U5502 : OAI22_X1 port map( A1 => n8103, A2 => n12196, B1 => n8104, B2 => 
                           n12190, ZN => n3925);
   U5503 : AOI221_X1 port map( B1 => n12208, B2 => n7211, C1 => n12202, C2 => 
                           n8705, A => n3906, ZN => n3903);
   U5504 : OAI22_X1 port map( A1 => n8086, A2 => n12196, B1 => n8087, B2 => 
                           n12190, ZN => n3906);
   U5505 : AOI221_X1 port map( B1 => n12208, B2 => n7214, C1 => n12202, C2 => 
                           n8704, A => n3887, ZN => n3884);
   U5506 : OAI22_X1 port map( A1 => n8069, A2 => n12196, B1 => n8070, B2 => 
                           n12190, ZN => n3887);
   U5507 : AOI221_X1 port map( B1 => n12208, B2 => n7217, C1 => n12202, C2 => 
                           n8703, A => n3868, ZN => n3865);
   U5508 : OAI22_X1 port map( A1 => n8052, A2 => n12196, B1 => n8053, B2 => 
                           n12190, ZN => n3868);
   U5509 : AOI221_X1 port map( B1 => n12208, B2 => n7220, C1 => n12202, C2 => 
                           n8702, A => n3849, ZN => n3846);
   U5510 : OAI22_X1 port map( A1 => n8035, A2 => n12196, B1 => n8036, B2 => 
                           n12190, ZN => n3849);
   U5511 : AOI221_X1 port map( B1 => n12208, B2 => n7223, C1 => n12202, C2 => 
                           n8701, A => n3830, ZN => n3827);
   U5512 : OAI22_X1 port map( A1 => n8018, A2 => n12196, B1 => n8019, B2 => 
                           n12190, ZN => n3830);
   U5513 : AOI221_X1 port map( B1 => n12208, B2 => n7226, C1 => n12202, C2 => 
                           n8700, A => n3811, ZN => n3808);
   U5514 : OAI22_X1 port map( A1 => n8001, A2 => n12196, B1 => n8002, B2 => 
                           n12190, ZN => n3811);
   U5515 : AOI221_X1 port map( B1 => n12208, B2 => n7229, C1 => n12202, C2 => 
                           n8699, A => n3792, ZN => n3789);
   U5516 : OAI22_X1 port map( A1 => n7984, A2 => n12196, B1 => n7985, B2 => 
                           n12190, ZN => n3792);
   U5517 : AOI221_X1 port map( B1 => n12209, B2 => n7232, C1 => n12203, C2 => 
                           n8698, A => n3773, ZN => n3770);
   U5518 : OAI22_X1 port map( A1 => n7967, A2 => n12197, B1 => n7968, B2 => 
                           n12191, ZN => n3773);
   U5519 : AOI221_X1 port map( B1 => n12209, B2 => n7245, C1 => n12203, C2 => 
                           n8697, A => n3754, ZN => n3751);
   U5520 : OAI22_X1 port map( A1 => n7950, A2 => n12197, B1 => n7951, B2 => 
                           n12191, ZN => n3754);
   U5521 : AOI221_X1 port map( B1 => n12209, B2 => n7278, C1 => n12203, C2 => 
                           n7279, A => n3735, ZN => n3732);
   U5522 : OAI22_X1 port map( A1 => n7933, A2 => n12197, B1 => n7934, B2 => 
                           n12191, ZN => n3735);
   U5523 : AOI221_X1 port map( B1 => n12209, B2 => n7282, C1 => n12203, C2 => 
                           n7283, A => n3716, ZN => n3713);
   U5524 : OAI22_X1 port map( A1 => n7916, A2 => n12197, B1 => n7917, B2 => 
                           n12191, ZN => n3716);
   U5525 : AOI221_X1 port map( B1 => n12209, B2 => n7286, C1 => n12203, C2 => 
                           n7287, A => n3697, ZN => n3694);
   U5526 : OAI22_X1 port map( A1 => n7899, A2 => n12197, B1 => n7900, B2 => 
                           n12191, ZN => n3697);
   U5527 : AOI221_X1 port map( B1 => n12209, B2 => n7290, C1 => n12203, C2 => 
                           n7291, A => n3678, ZN => n3675);
   U5528 : OAI22_X1 port map( A1 => n7882, A2 => n12197, B1 => n7883, B2 => 
                           n12191, ZN => n3678);
   U5529 : AOI221_X1 port map( B1 => n12209, B2 => n7294, C1 => n12203, C2 => 
                           n7295, A => n3659, ZN => n3656);
   U5530 : OAI22_X1 port map( A1 => n7865, A2 => n12197, B1 => n7866, B2 => 
                           n12191, ZN => n3659);
   U5531 : AOI221_X1 port map( B1 => n12209, B2 => n7298, C1 => n12203, C2 => 
                           n7299, A => n3640, ZN => n3637);
   U5532 : OAI22_X1 port map( A1 => n7848, A2 => n12197, B1 => n7849, B2 => 
                           n12191, ZN => n3640);
   U5533 : AOI221_X1 port map( B1 => n12209, B2 => n7302, C1 => n12203, C2 => 
                           n7303, A => n3621, ZN => n3618);
   U5534 : OAI22_X1 port map( A1 => n7831, A2 => n12197, B1 => n7832, B2 => 
                           n12191, ZN => n3621);
   U5535 : AOI221_X1 port map( B1 => n12209, B2 => n7306, C1 => n12203, C2 => 
                           n7307, A => n3602, ZN => n3599);
   U5536 : OAI22_X1 port map( A1 => n7814, A2 => n12197, B1 => n7815, B2 => 
                           n12191, ZN => n3602);
   U5537 : AOI221_X1 port map( B1 => n12209, B2 => n7310, C1 => n12203, C2 => 
                           n7311, A => n3583, ZN => n3580);
   U5538 : OAI22_X1 port map( A1 => n7797, A2 => n12197, B1 => n7798, B2 => 
                           n12191, ZN => n3583);
   U5539 : AOI221_X1 port map( B1 => n12209, B2 => n7314, C1 => n12203, C2 => 
                           n7315, A => n3564, ZN => n3561);
   U5540 : OAI22_X1 port map( A1 => n7780, A2 => n12197, B1 => n7781, B2 => 
                           n12191, ZN => n3564);
   U5541 : AOI221_X1 port map( B1 => n12210, B2 => n7318, C1 => n12204, C2 => 
                           n7319, A => n3545, ZN => n3542);
   U5542 : OAI22_X1 port map( A1 => n7763, A2 => n12198, B1 => n7764, B2 => 
                           n12192, ZN => n3545);
   U5543 : AOI221_X1 port map( B1 => n12210, B2 => n7322, C1 => n12204, C2 => 
                           n7323, A => n3526, ZN => n3523);
   U5544 : OAI22_X1 port map( A1 => n7746, A2 => n12198, B1 => n7747, B2 => 
                           n12192, ZN => n3526);
   U5545 : AOI221_X1 port map( B1 => n12210, B2 => n4486, C1 => n12204, C2 => 
                           n4487, A => n3507, ZN => n3504);
   U5546 : OAI22_X1 port map( A1 => n7644, A2 => n12198, B1 => n7645, B2 => 
                           n12192, ZN => n3507);
   U5547 : AOI221_X1 port map( B1 => n12210, B2 => n4488, C1 => n12204, C2 => 
                           n4489, A => n3488, ZN => n3485);
   U5548 : OAI22_X1 port map( A1 => n7627, A2 => n12198, B1 => n7628, B2 => 
                           n12192, ZN => n3488);
   U5549 : AOI221_X1 port map( B1 => n12210, B2 => n4490, C1 => n12204, C2 => 
                           n4491, A => n3469, ZN => n3466);
   U5550 : OAI22_X1 port map( A1 => n7523, A2 => n12198, B1 => n7524, B2 => 
                           n12192, ZN => n3469);
   U5551 : AOI221_X1 port map( B1 => n12210, B2 => n4492, C1 => n12204, C2 => 
                           n4493, A => n3450, ZN => n3447);
   U5552 : OAI22_X1 port map( A1 => n7506, A2 => n12198, B1 => n7507, B2 => 
                           n12192, ZN => n3450);
   U5553 : AOI221_X1 port map( B1 => n12210, B2 => n4494, C1 => n12204, C2 => 
                           n4495, A => n3431, ZN => n3428);
   U5554 : OAI22_X1 port map( A1 => n7404, A2 => n12198, B1 => n7490, B2 => 
                           n12192, ZN => n3431);
   U5555 : AOI221_X1 port map( B1 => n12210, B2 => n4496, C1 => n12204, C2 => 
                           n4497, A => n3412, ZN => n3409);
   U5556 : OAI22_X1 port map( A1 => n7387, A2 => n12198, B1 => n7388, B2 => 
                           n12192, ZN => n3412);
   U5557 : AOI221_X1 port map( B1 => n12210, B2 => n4498, C1 => n12204, C2 => 
                           n4499, A => n3393, ZN => n3390);
   U5558 : OAI22_X1 port map( A1 => n7370, A2 => n12198, B1 => n7371, B2 => 
                           n12192, ZN => n3393);
   U5559 : AOI221_X1 port map( B1 => n12210, B2 => n4500, C1 => n12204, C2 => 
                           n4501, A => n3374, ZN => n3371);
   U5560 : OAI22_X1 port map( A1 => n7271, A2 => n12198, B1 => n7272, B2 => 
                           n12192, ZN => n3374);
   U5561 : AOI221_X1 port map( B1 => n12210, B2 => n4502, C1 => n12204, C2 => 
                           n4503, A => n3355, ZN => n3352);
   U5562 : OAI22_X1 port map( A1 => n7254, A2 => n12198, B1 => n7255, B2 => 
                           n12192, ZN => n3355);
   U5563 : AOI221_X1 port map( B1 => n12210, B2 => n4684, C1 => n12204, C2 => 
                           n4685, A => n3336, ZN => n3333);
   U5564 : OAI22_X1 port map( A1 => n7237, A2 => n12198, B1 => n7238, B2 => 
                           n12192, ZN => n3336);
   U5565 : AOI221_X1 port map( B1 => n12211, B2 => n4504, C1 => n12205, C2 => 
                           n4505, A => n3317, ZN => n3314);
   U5566 : OAI22_X1 port map( A1 => n7140, A2 => n12199, B1 => n7141, B2 => 
                           n12193, ZN => n3317);
   U5567 : AOI221_X1 port map( B1 => n12211, B2 => n4506, C1 => n12205, C2 => 
                           n4507, A => n3298, ZN => n3295);
   U5568 : OAI22_X1 port map( A1 => n7123, A2 => n12199, B1 => n7124, B2 => 
                           n12193, ZN => n3298);
   U5569 : AOI221_X1 port map( B1 => n12211, B2 => n4508, C1 => n12205, C2 => 
                           n4509, A => n3279, ZN => n3276);
   U5570 : OAI22_X1 port map( A1 => n7106, A2 => n12199, B1 => n7107, B2 => 
                           n12193, ZN => n3279);
   U5571 : AOI221_X1 port map( B1 => n12211, B2 => n4510, C1 => n12205, C2 => 
                           n4511, A => n3250, ZN => n3241);
   U5572 : OAI22_X1 port map( A1 => n4845, A2 => n12199, B1 => n4846, B2 => 
                           n12193, ZN => n3250);
   U5573 : INV_X1 port map( A => ADD_RD2(3), ZN => n13388);
   U5574 : INV_X1 port map( A => ADD_RD2(0), ZN => n13391);
   U5575 : INV_X1 port map( A => ADD_RD2(4), ZN => n13387);
   U5576 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n1922);
   U5577 : NAND2_X1 port map( A1 => DATAIN(63), A2 => n12132, ZN => n1841);
   U5578 : OAI21_X1 port map( B1 => n8568, B2 => n12339, A => n4441, ZN => 
                           n4862);
   U5579 : OAI21_X1 port map( B1 => n4442, B2 => n4443, A => n12344, ZN => 
                           n4441);
   U5580 : NAND4_X1 port map( A1 => n4460, A2 => n4461, A3 => n4462, A4 => 
                           n4463, ZN => n4442);
   U5581 : NAND4_X1 port map( A1 => n4444, A2 => n4445, A3 => n4446, A4 => 
                           n4447, ZN => n4443);
   U5582 : OAI21_X1 port map( B1 => n8551, B2 => n12338, A => n4422, ZN => 
                           n4863);
   U5583 : OAI21_X1 port map( B1 => n4423, B2 => n4424, A => n12344, ZN => 
                           n4422);
   U5584 : NAND4_X1 port map( A1 => n4433, A2 => n4434, A3 => n4435, A4 => 
                           n4436, ZN => n4423);
   U5585 : NAND4_X1 port map( A1 => n4425, A2 => n4426, A3 => n4427, A4 => 
                           n4428, ZN => n4424);
   U5586 : OAI21_X1 port map( B1 => n8534, B2 => n12339, A => n4403, ZN => 
                           n4864);
   U5587 : OAI21_X1 port map( B1 => n4404, B2 => n4405, A => n12344, ZN => 
                           n4403);
   U5588 : NAND4_X1 port map( A1 => n4414, A2 => n4415, A3 => n4416, A4 => 
                           n4417, ZN => n4404);
   U5589 : NAND4_X1 port map( A1 => n4406, A2 => n4407, A3 => n4408, A4 => 
                           n4409, ZN => n4405);
   U5590 : OAI21_X1 port map( B1 => n8517, B2 => n12338, A => n4384, ZN => 
                           n4865);
   U5591 : OAI21_X1 port map( B1 => n4385, B2 => n4386, A => n12343, ZN => 
                           n4384);
   U5592 : NAND4_X1 port map( A1 => n4395, A2 => n4396, A3 => n4397, A4 => 
                           n4398, ZN => n4385);
   U5593 : NAND4_X1 port map( A1 => n4387, A2 => n4388, A3 => n4389, A4 => 
                           n4390, ZN => n4386);
   U5594 : OAI21_X1 port map( B1 => n8500, B2 => n12338, A => n4365, ZN => 
                           n4866);
   U5595 : OAI21_X1 port map( B1 => n4366, B2 => n4367, A => n12343, ZN => 
                           n4365);
   U5596 : NAND4_X1 port map( A1 => n4376, A2 => n4377, A3 => n4378, A4 => 
                           n4379, ZN => n4366);
   U5597 : NAND4_X1 port map( A1 => n4368, A2 => n4369, A3 => n4370, A4 => 
                           n4371, ZN => n4367);
   U5598 : OAI21_X1 port map( B1 => n8483, B2 => n12339, A => n4346, ZN => 
                           n4867);
   U5599 : OAI21_X1 port map( B1 => n4347, B2 => n4348, A => n12343, ZN => 
                           n4346);
   U5600 : NAND4_X1 port map( A1 => n4357, A2 => n4358, A3 => n4359, A4 => 
                           n4360, ZN => n4347);
   U5601 : NAND4_X1 port map( A1 => n4349, A2 => n4350, A3 => n4351, A4 => 
                           n4352, ZN => n4348);
   U5602 : OAI21_X1 port map( B1 => n8466, B2 => n12339, A => n4327, ZN => 
                           n4868);
   U5603 : OAI21_X1 port map( B1 => n4328, B2 => n4329, A => n12343, ZN => 
                           n4327);
   U5604 : NAND4_X1 port map( A1 => n4338, A2 => n4339, A3 => n4340, A4 => 
                           n4341, ZN => n4328);
   U5605 : NAND4_X1 port map( A1 => n4330, A2 => n4331, A3 => n4332, A4 => 
                           n4333, ZN => n4329);
   U5606 : OAI21_X1 port map( B1 => n8449, B2 => n12338, A => n4308, ZN => 
                           n4869);
   U5607 : OAI21_X1 port map( B1 => n4309, B2 => n4310, A => n12343, ZN => 
                           n4308);
   U5608 : NAND4_X1 port map( A1 => n4319, A2 => n4320, A3 => n4321, A4 => 
                           n4322, ZN => n4309);
   U5609 : NAND4_X1 port map( A1 => n4311, A2 => n4312, A3 => n4313, A4 => 
                           n4314, ZN => n4310);
   U5610 : OAI21_X1 port map( B1 => n8432, B2 => n12338, A => n4289, ZN => 
                           n4870);
   U5611 : OAI21_X1 port map( B1 => n4290, B2 => n4291, A => n12342, ZN => 
                           n4289);
   U5612 : NAND4_X1 port map( A1 => n4300, A2 => n4301, A3 => n4302, A4 => 
                           n4303, ZN => n4290);
   U5613 : NAND4_X1 port map( A1 => n4292, A2 => n4293, A3 => n4294, A4 => 
                           n4295, ZN => n4291);
   U5614 : OAI21_X1 port map( B1 => n8415, B2 => n12338, A => n4270, ZN => 
                           n4871);
   U5615 : OAI21_X1 port map( B1 => n4271, B2 => n4272, A => n12342, ZN => 
                           n4270);
   U5616 : NAND4_X1 port map( A1 => n4281, A2 => n4282, A3 => n4283, A4 => 
                           n4284, ZN => n4271);
   U5617 : NAND4_X1 port map( A1 => n4273, A2 => n4274, A3 => n4275, A4 => 
                           n4276, ZN => n4272);
   U5618 : OAI21_X1 port map( B1 => n8398, B2 => n12337, A => n4251, ZN => 
                           n4872);
   U5619 : OAI21_X1 port map( B1 => n4252, B2 => n4253, A => n12341, ZN => 
                           n4251);
   U5620 : NAND4_X1 port map( A1 => n4262, A2 => n4263, A3 => n4264, A4 => 
                           n4265, ZN => n4252);
   U5621 : NAND4_X1 port map( A1 => n4254, A2 => n4255, A3 => n4256, A4 => 
                           n4257, ZN => n4253);
   U5622 : OAI21_X1 port map( B1 => n8381, B2 => n12338, A => n4232, ZN => 
                           n4873);
   U5623 : OAI21_X1 port map( B1 => n4233, B2 => n4234, A => n12341, ZN => 
                           n4232);
   U5624 : NAND4_X1 port map( A1 => n4243, A2 => n4244, A3 => n4245, A4 => 
                           n4246, ZN => n4233);
   U5625 : NAND4_X1 port map( A1 => n4235, A2 => n4236, A3 => n4237, A4 => 
                           n4238, ZN => n4234);
   U5626 : OAI21_X1 port map( B1 => n8364, B2 => n12338, A => n4213, ZN => 
                           n4874);
   U5627 : OAI21_X1 port map( B1 => n4214, B2 => n4215, A => n12341, ZN => 
                           n4213);
   U5628 : NAND4_X1 port map( A1 => n4224, A2 => n4225, A3 => n4226, A4 => 
                           n4227, ZN => n4214);
   U5629 : NAND4_X1 port map( A1 => n4216, A2 => n4217, A3 => n4218, A4 => 
                           n4219, ZN => n4215);
   U5630 : OAI21_X1 port map( B1 => n8347, B2 => n12338, A => n4194, ZN => 
                           n4875);
   U5631 : OAI21_X1 port map( B1 => n4195, B2 => n4196, A => n12340, ZN => 
                           n4194);
   U5632 : NAND4_X1 port map( A1 => n4205, A2 => n4206, A3 => n4207, A4 => 
                           n4208, ZN => n4195);
   U5633 : NAND4_X1 port map( A1 => n4197, A2 => n4198, A3 => n4199, A4 => 
                           n4200, ZN => n4196);
   U5634 : OAI21_X1 port map( B1 => n8330, B2 => n12338, A => n4175, ZN => 
                           n4876);
   U5635 : OAI21_X1 port map( B1 => n4176, B2 => n4177, A => n12342, ZN => 
                           n4175);
   U5636 : NAND4_X1 port map( A1 => n4186, A2 => n4187, A3 => n4188, A4 => 
                           n4189, ZN => n4176);
   U5637 : NAND4_X1 port map( A1 => n4178, A2 => n4179, A3 => n4180, A4 => 
                           n4181, ZN => n4177);
   U5638 : OAI21_X1 port map( B1 => n8313, B2 => n12338, A => n4156, ZN => 
                           n4877);
   U5639 : OAI21_X1 port map( B1 => n4157, B2 => n4158, A => n12341, ZN => 
                           n4156);
   U5640 : NAND4_X1 port map( A1 => n4167, A2 => n4168, A3 => n4169, A4 => 
                           n4170, ZN => n4157);
   U5641 : NAND4_X1 port map( A1 => n4159, A2 => n4160, A3 => n4161, A4 => 
                           n4162, ZN => n4158);
   U5642 : OAI21_X1 port map( B1 => n8296, B2 => n12337, A => n4137, ZN => 
                           n4878);
   U5643 : OAI21_X1 port map( B1 => n4138, B2 => n4139, A => n12339, ZN => 
                           n4137);
   U5644 : NAND4_X1 port map( A1 => n4148, A2 => n4149, A3 => n4150, A4 => 
                           n4151, ZN => n4138);
   U5645 : NAND4_X1 port map( A1 => n4140, A2 => n4141, A3 => n4142, A4 => 
                           n4143, ZN => n4139);
   U5646 : OAI21_X1 port map( B1 => n8279, B2 => n12337, A => n4118, ZN => 
                           n4879);
   U5647 : OAI21_X1 port map( B1 => n4119, B2 => n4120, A => n12341, ZN => 
                           n4118);
   U5648 : NAND4_X1 port map( A1 => n4129, A2 => n4130, A3 => n4131, A4 => 
                           n4132, ZN => n4119);
   U5649 : NAND4_X1 port map( A1 => n4121, A2 => n4122, A3 => n4123, A4 => 
                           n4124, ZN => n4120);
   U5650 : OAI21_X1 port map( B1 => n8262, B2 => n12338, A => n4099, ZN => 
                           n4880);
   U5651 : OAI21_X1 port map( B1 => n4100, B2 => n4101, A => n12340, ZN => 
                           n4099);
   U5652 : NAND4_X1 port map( A1 => n4110, A2 => n4111, A3 => n4112, A4 => 
                           n4113, ZN => n4100);
   U5653 : NAND4_X1 port map( A1 => n4102, A2 => n4103, A3 => n4104, A4 => 
                           n4105, ZN => n4101);
   U5654 : OAI21_X1 port map( B1 => n8245, B2 => n12337, A => n4080, ZN => 
                           n4881);
   U5655 : OAI21_X1 port map( B1 => n4081, B2 => n4082, A => n12341, ZN => 
                           n4080);
   U5656 : NAND4_X1 port map( A1 => n4091, A2 => n4092, A3 => n4093, A4 => 
                           n4094, ZN => n4081);
   U5657 : NAND4_X1 port map( A1 => n4083, A2 => n4084, A3 => n4085, A4 => 
                           n4086, ZN => n4082);
   U5658 : OAI21_X1 port map( B1 => n8228, B2 => n12337, A => n4061, ZN => 
                           n4882);
   U5659 : OAI21_X1 port map( B1 => n4062, B2 => n4063, A => n12339, ZN => 
                           n4061);
   U5660 : NAND4_X1 port map( A1 => n4072, A2 => n4073, A3 => n4074, A4 => 
                           n4075, ZN => n4062);
   U5661 : NAND4_X1 port map( A1 => n4064, A2 => n4065, A3 => n4066, A4 => 
                           n4067, ZN => n4063);
   U5662 : OAI21_X1 port map( B1 => n8211, B2 => n12337, A => n4042, ZN => 
                           n4883);
   U5663 : OAI21_X1 port map( B1 => n4043, B2 => n4044, A => n12340, ZN => 
                           n4042);
   U5664 : NAND4_X1 port map( A1 => n4053, A2 => n4054, A3 => n4055, A4 => 
                           n4056, ZN => n4043);
   U5665 : NAND4_X1 port map( A1 => n4045, A2 => n4046, A3 => n4047, A4 => 
                           n4048, ZN => n4044);
   U5666 : OAI21_X1 port map( B1 => n8194, B2 => n12337, A => n4023, ZN => 
                           n4884);
   U5667 : OAI21_X1 port map( B1 => n4024, B2 => n4025, A => n12339, ZN => 
                           n4023);
   U5668 : NAND4_X1 port map( A1 => n4034, A2 => n4035, A3 => n4036, A4 => 
                           n4037, ZN => n4024);
   U5669 : NAND4_X1 port map( A1 => n4026, A2 => n4027, A3 => n4028, A4 => 
                           n4029, ZN => n4025);
   U5670 : OAI21_X1 port map( B1 => n8177, B2 => n12337, A => n4004, ZN => 
                           n4885);
   U5671 : OAI21_X1 port map( B1 => n4005, B2 => n4006, A => n12340, ZN => 
                           n4004);
   U5672 : NAND4_X1 port map( A1 => n4015, A2 => n4016, A3 => n4017, A4 => 
                           n4018, ZN => n4005);
   U5673 : NAND4_X1 port map( A1 => n4007, A2 => n4008, A3 => n4009, A4 => 
                           n4010, ZN => n4006);
   U5674 : OAI21_X1 port map( B1 => n8160, B2 => n12337, A => n3985, ZN => 
                           n4886);
   U5675 : OAI21_X1 port map( B1 => n3986, B2 => n3987, A => n12339, ZN => 
                           n3985);
   U5676 : NAND4_X1 port map( A1 => n3996, A2 => n3997, A3 => n3998, A4 => 
                           n3999, ZN => n3986);
   U5677 : NAND4_X1 port map( A1 => n3988, A2 => n3989, A3 => n3990, A4 => 
                           n3991, ZN => n3987);
   U5678 : OAI21_X1 port map( B1 => n8143, B2 => n12337, A => n3966, ZN => 
                           n4887);
   U5679 : OAI21_X1 port map( B1 => n3967, B2 => n3968, A => n12340, ZN => 
                           n3966);
   U5680 : NAND4_X1 port map( A1 => n3977, A2 => n3978, A3 => n3979, A4 => 
                           n3980, ZN => n3967);
   U5681 : NAND4_X1 port map( A1 => n3969, A2 => n3970, A3 => n3971, A4 => 
                           n3972, ZN => n3968);
   U5682 : OAI21_X1 port map( B1 => n8126, B2 => n12337, A => n3947, ZN => 
                           n4888);
   U5683 : OAI21_X1 port map( B1 => n3948, B2 => n3949, A => n12340, ZN => 
                           n3947);
   U5684 : NAND4_X1 port map( A1 => n3958, A2 => n3959, A3 => n3960, A4 => 
                           n3961, ZN => n3948);
   U5685 : NAND4_X1 port map( A1 => n3950, A2 => n3951, A3 => n3952, A4 => 
                           n3953, ZN => n3949);
   U5686 : OAI21_X1 port map( B1 => n8109, B2 => n12336, A => n3928, ZN => 
                           n4889);
   U5687 : OAI21_X1 port map( B1 => n3929, B2 => n3930, A => n12339, ZN => 
                           n3928);
   U5688 : NAND4_X1 port map( A1 => n3939, A2 => n3940, A3 => n3941, A4 => 
                           n3942, ZN => n3929);
   U5689 : NAND4_X1 port map( A1 => n3931, A2 => n3932, A3 => n3933, A4 => 
                           n3934, ZN => n3930);
   U5690 : OAI21_X1 port map( B1 => n8092, B2 => n12336, A => n3909, ZN => 
                           n4890);
   U5691 : OAI21_X1 port map( B1 => n3910, B2 => n3911, A => n12339, ZN => 
                           n3909);
   U5692 : NAND4_X1 port map( A1 => n3920, A2 => n3921, A3 => n3922, A4 => 
                           n3923, ZN => n3910);
   U5693 : NAND4_X1 port map( A1 => n3912, A2 => n3913, A3 => n3914, A4 => 
                           n3915, ZN => n3911);
   U5694 : OAI21_X1 port map( B1 => n8075, B2 => n12336, A => n3890, ZN => 
                           n4891);
   U5695 : OAI21_X1 port map( B1 => n3891, B2 => n3892, A => n12340, ZN => 
                           n3890);
   U5696 : NAND4_X1 port map( A1 => n3901, A2 => n3902, A3 => n3903, A4 => 
                           n3904, ZN => n3891);
   U5697 : NAND4_X1 port map( A1 => n3893, A2 => n3894, A3 => n3895, A4 => 
                           n3896, ZN => n3892);
   U5698 : OAI21_X1 port map( B1 => n8058, B2 => n12336, A => n3871, ZN => 
                           n4892);
   U5699 : OAI21_X1 port map( B1 => n3872, B2 => n3873, A => n12339, ZN => 
                           n3871);
   U5700 : NAND4_X1 port map( A1 => n3882, A2 => n3883, A3 => n3884, A4 => 
                           n3885, ZN => n3872);
   U5701 : NAND4_X1 port map( A1 => n3874, A2 => n3875, A3 => n3876, A4 => 
                           n3877, ZN => n3873);
   U5702 : OAI21_X1 port map( B1 => n8041, B2 => n12337, A => n3852, ZN => 
                           n4893);
   U5703 : OAI21_X1 port map( B1 => n3853, B2 => n3854, A => n12339, ZN => 
                           n3852);
   U5704 : NAND4_X1 port map( A1 => n3863, A2 => n3864, A3 => n3865, A4 => 
                           n3866, ZN => n3853);
   U5705 : NAND4_X1 port map( A1 => n3855, A2 => n3856, A3 => n3857, A4 => 
                           n3858, ZN => n3854);
   U5706 : OAI21_X1 port map( B1 => n8024, B2 => n12336, A => n3833, ZN => 
                           n4894);
   U5707 : OAI21_X1 port map( B1 => n3834, B2 => n3835, A => n12340, ZN => 
                           n3833);
   U5708 : NAND4_X1 port map( A1 => n3844, A2 => n3845, A3 => n3846, A4 => 
                           n3847, ZN => n3834);
   U5709 : NAND4_X1 port map( A1 => n3836, A2 => n3837, A3 => n3838, A4 => 
                           n3839, ZN => n3835);
   U5710 : OAI21_X1 port map( B1 => n8007, B2 => n12336, A => n3814, ZN => 
                           n4895);
   U5711 : OAI21_X1 port map( B1 => n3815, B2 => n3816, A => n12340, ZN => 
                           n3814);
   U5712 : NAND4_X1 port map( A1 => n3825, A2 => n3826, A3 => n3827, A4 => 
                           n3828, ZN => n3815);
   U5713 : NAND4_X1 port map( A1 => n3817, A2 => n3818, A3 => n3819, A4 => 
                           n3820, ZN => n3816);
   U5714 : OAI21_X1 port map( B1 => n7990, B2 => n12336, A => n3795, ZN => 
                           n4896);
   U5715 : OAI21_X1 port map( B1 => n3796, B2 => n3797, A => n12340, ZN => 
                           n3795);
   U5716 : NAND4_X1 port map( A1 => n3806, A2 => n3807, A3 => n3808, A4 => 
                           n3809, ZN => n3796);
   U5717 : NAND4_X1 port map( A1 => n3798, A2 => n3799, A3 => n3800, A4 => 
                           n3801, ZN => n3797);
   U5718 : OAI21_X1 port map( B1 => n7973, B2 => n12336, A => n3776, ZN => 
                           n4897);
   U5719 : OAI21_X1 port map( B1 => n3777, B2 => n3778, A => n12341, ZN => 
                           n3776);
   U5720 : NAND4_X1 port map( A1 => n3787, A2 => n3788, A3 => n3789, A4 => 
                           n3790, ZN => n3777);
   U5721 : NAND4_X1 port map( A1 => n3779, A2 => n3780, A3 => n3781, A4 => 
                           n3782, ZN => n3778);
   U5722 : OAI21_X1 port map( B1 => n7956, B2 => n12336, A => n3757, ZN => 
                           n4898);
   U5723 : OAI21_X1 port map( B1 => n3758, B2 => n3759, A => n12340, ZN => 
                           n3757);
   U5724 : NAND4_X1 port map( A1 => n3768, A2 => n3769, A3 => n3770, A4 => 
                           n3771, ZN => n3758);
   U5725 : NAND4_X1 port map( A1 => n3760, A2 => n3761, A3 => n3762, A4 => 
                           n3763, ZN => n3759);
   U5726 : OAI21_X1 port map( B1 => n7939, B2 => n12336, A => n3738, ZN => 
                           n4899);
   U5727 : OAI21_X1 port map( B1 => n3739, B2 => n3740, A => n12340, ZN => 
                           n3738);
   U5728 : NAND4_X1 port map( A1 => n3749, A2 => n3750, A3 => n3751, A4 => 
                           n3752, ZN => n3739);
   U5729 : NAND4_X1 port map( A1 => n3741, A2 => n3742, A3 => n3743, A4 => 
                           n3744, ZN => n3740);
   U5730 : OAI21_X1 port map( B1 => n7922, B2 => n12336, A => n3719, ZN => 
                           n4900);
   U5731 : OAI21_X1 port map( B1 => n3720, B2 => n3721, A => n12342, ZN => 
                           n3719);
   U5732 : NAND4_X1 port map( A1 => n3730, A2 => n3731, A3 => n3732, A4 => 
                           n3733, ZN => n3720);
   U5733 : NAND4_X1 port map( A1 => n3722, A2 => n3723, A3 => n3724, A4 => 
                           n3725, ZN => n3721);
   U5734 : OAI21_X1 port map( B1 => n7905, B2 => n12335, A => n3700, ZN => 
                           n4901);
   U5735 : OAI21_X1 port map( B1 => n3701, B2 => n3702, A => n12342, ZN => 
                           n3700);
   U5736 : NAND4_X1 port map( A1 => n3711, A2 => n3712, A3 => n3713, A4 => 
                           n3714, ZN => n3701);
   U5737 : NAND4_X1 port map( A1 => n3703, A2 => n3704, A3 => n3705, A4 => 
                           n3706, ZN => n3702);
   U5738 : OAI21_X1 port map( B1 => n7888, B2 => n12335, A => n3681, ZN => 
                           n4902);
   U5739 : OAI21_X1 port map( B1 => n3682, B2 => n3683, A => n12341, ZN => 
                           n3681);
   U5740 : NAND4_X1 port map( A1 => n3692, A2 => n3693, A3 => n3694, A4 => 
                           n3695, ZN => n3682);
   U5741 : NAND4_X1 port map( A1 => n3684, A2 => n3685, A3 => n3686, A4 => 
                           n3687, ZN => n3683);
   U5742 : OAI21_X1 port map( B1 => n7871, B2 => n12335, A => n3662, ZN => 
                           n4903);
   U5743 : OAI21_X1 port map( B1 => n3663, B2 => n3664, A => n12341, ZN => 
                           n3662);
   U5744 : NAND4_X1 port map( A1 => n3673, A2 => n3674, A3 => n3675, A4 => 
                           n3676, ZN => n3663);
   U5745 : NAND4_X1 port map( A1 => n3665, A2 => n3666, A3 => n3667, A4 => 
                           n3668, ZN => n3664);
   U5746 : OAI21_X1 port map( B1 => n7854, B2 => n12335, A => n3643, ZN => 
                           n4904);
   U5747 : OAI21_X1 port map( B1 => n3644, B2 => n3645, A => n12341, ZN => 
                           n3643);
   U5748 : NAND4_X1 port map( A1 => n3654, A2 => n3655, A3 => n3656, A4 => 
                           n3657, ZN => n3644);
   U5749 : NAND4_X1 port map( A1 => n3646, A2 => n3647, A3 => n3648, A4 => 
                           n3649, ZN => n3645);
   U5750 : OAI21_X1 port map( B1 => n7837, B2 => n12335, A => n3624, ZN => 
                           n4905);
   U5751 : OAI21_X1 port map( B1 => n3625, B2 => n3626, A => n12341, ZN => 
                           n3624);
   U5752 : NAND4_X1 port map( A1 => n3635, A2 => n3636, A3 => n3637, A4 => 
                           n3638, ZN => n3625);
   U5753 : NAND4_X1 port map( A1 => n3627, A2 => n3628, A3 => n3629, A4 => 
                           n3630, ZN => n3626);
   U5754 : OAI21_X1 port map( B1 => n7820, B2 => n12335, A => n3605, ZN => 
                           n4906);
   U5755 : OAI21_X1 port map( B1 => n3606, B2 => n3607, A => n12342, ZN => 
                           n3605);
   U5756 : NAND4_X1 port map( A1 => n3616, A2 => n3617, A3 => n3618, A4 => 
                           n3619, ZN => n3606);
   U5757 : NAND4_X1 port map( A1 => n3608, A2 => n3609, A3 => n3610, A4 => 
                           n3611, ZN => n3607);
   U5758 : OAI21_X1 port map( B1 => n7803, B2 => n12335, A => n3586, ZN => 
                           n4907);
   U5759 : OAI21_X1 port map( B1 => n3587, B2 => n3588, A => n12341, ZN => 
                           n3586);
   U5760 : NAND4_X1 port map( A1 => n3597, A2 => n3598, A3 => n3599, A4 => 
                           n3600, ZN => n3587);
   U5761 : NAND4_X1 port map( A1 => n3589, A2 => n3590, A3 => n3591, A4 => 
                           n3592, ZN => n3588);
   U5762 : OAI21_X1 port map( B1 => n7786, B2 => n12335, A => n3567, ZN => 
                           n4908);
   U5763 : OAI21_X1 port map( B1 => n3568, B2 => n3569, A => n12342, ZN => 
                           n3567);
   U5764 : NAND4_X1 port map( A1 => n3578, A2 => n3579, A3 => n3580, A4 => 
                           n3581, ZN => n3568);
   U5765 : NAND4_X1 port map( A1 => n3570, A2 => n3571, A3 => n3572, A4 => 
                           n3573, ZN => n3569);
   U5766 : OAI21_X1 port map( B1 => n7769, B2 => n12335, A => n3548, ZN => 
                           n4909);
   U5767 : OAI21_X1 port map( B1 => n3549, B2 => n3550, A => n12342, ZN => 
                           n3548);
   U5768 : NAND4_X1 port map( A1 => n3559, A2 => n3560, A3 => n3561, A4 => 
                           n3562, ZN => n3549);
   U5769 : NAND4_X1 port map( A1 => n3551, A2 => n3552, A3 => n3553, A4 => 
                           n3554, ZN => n3550);
   U5770 : OAI21_X1 port map( B1 => n7752, B2 => n12335, A => n3529, ZN => 
                           n4910);
   U5771 : OAI21_X1 port map( B1 => n3530, B2 => n3531, A => n12342, ZN => 
                           n3529);
   U5772 : NAND4_X1 port map( A1 => n3540, A2 => n3541, A3 => n3542, A4 => 
                           n3543, ZN => n3530);
   U5773 : NAND4_X1 port map( A1 => n3532, A2 => n3533, A3 => n3534, A4 => 
                           n3535, ZN => n3531);
   U5774 : OAI21_X1 port map( B1 => n7650, B2 => n12335, A => n3510, ZN => 
                           n4911);
   U5775 : OAI21_X1 port map( B1 => n3511, B2 => n3512, A => n12342, ZN => 
                           n3510);
   U5776 : NAND4_X1 port map( A1 => n3521, A2 => n3522, A3 => n3523, A4 => 
                           n3524, ZN => n3511);
   U5777 : NAND4_X1 port map( A1 => n3513, A2 => n3514, A3 => n3515, A4 => 
                           n3516, ZN => n3512);
   U5778 : OAI21_X1 port map( B1 => n7633, B2 => n12335, A => n3491, ZN => 
                           n4912);
   U5779 : OAI21_X1 port map( B1 => n3492, B2 => n3493, A => n12343, ZN => 
                           n3491);
   U5780 : NAND4_X1 port map( A1 => n3502, A2 => n3503, A3 => n3504, A4 => 
                           n3505, ZN => n3492);
   U5781 : NAND4_X1 port map( A1 => n3494, A2 => n3495, A3 => n3496, A4 => 
                           n3497, ZN => n3493);
   U5782 : OAI21_X1 port map( B1 => n7529, B2 => n12334, A => n3472, ZN => 
                           n4913);
   U5783 : OAI21_X1 port map( B1 => n3473, B2 => n3474, A => n12342, ZN => 
                           n3472);
   U5784 : NAND4_X1 port map( A1 => n3483, A2 => n3484, A3 => n3485, A4 => 
                           n3486, ZN => n3473);
   U5785 : NAND4_X1 port map( A1 => n3475, A2 => n3476, A3 => n3477, A4 => 
                           n3478, ZN => n3474);
   U5786 : OAI21_X1 port map( B1 => n7512, B2 => n12334, A => n3453, ZN => 
                           n4914);
   U5787 : OAI21_X1 port map( B1 => n3454, B2 => n3455, A => n12342, ZN => 
                           n3453);
   U5788 : NAND4_X1 port map( A1 => n3464, A2 => n3465, A3 => n3466, A4 => 
                           n3467, ZN => n3454);
   U5789 : NAND4_X1 port map( A1 => n3456, A2 => n3457, A3 => n3458, A4 => 
                           n3459, ZN => n3455);
   U5790 : OAI21_X1 port map( B1 => n7495, B2 => n12334, A => n3434, ZN => 
                           n4915);
   U5791 : OAI21_X1 port map( B1 => n3435, B2 => n3436, A => n12343, ZN => 
                           n3434);
   U5792 : NAND4_X1 port map( A1 => n3445, A2 => n3446, A3 => n3447, A4 => 
                           n3448, ZN => n3435);
   U5793 : NAND4_X1 port map( A1 => n3437, A2 => n3438, A3 => n3439, A4 => 
                           n3440, ZN => n3436);
   U5794 : OAI21_X1 port map( B1 => n7393, B2 => n12334, A => n3415, ZN => 
                           n4916);
   U5795 : OAI21_X1 port map( B1 => n3416, B2 => n3417, A => n12343, ZN => 
                           n3415);
   U5796 : NAND4_X1 port map( A1 => n3426, A2 => n3427, A3 => n3428, A4 => 
                           n3429, ZN => n3416);
   U5797 : NAND4_X1 port map( A1 => n3418, A2 => n3419, A3 => n3420, A4 => 
                           n3421, ZN => n3417);
   U5798 : OAI21_X1 port map( B1 => n7376, B2 => n12334, A => n3396, ZN => 
                           n4917);
   U5799 : OAI21_X1 port map( B1 => n3397, B2 => n3398, A => n12343, ZN => 
                           n3396);
   U5800 : NAND4_X1 port map( A1 => n3407, A2 => n3408, A3 => n3409, A4 => 
                           n3410, ZN => n3397);
   U5801 : NAND4_X1 port map( A1 => n3399, A2 => n3400, A3 => n3401, A4 => 
                           n3402, ZN => n3398);
   U5802 : OAI21_X1 port map( B1 => n7277, B2 => n12334, A => n3377, ZN => 
                           n4918);
   U5803 : OAI21_X1 port map( B1 => n3378, B2 => n3379, A => n12343, ZN => 
                           n3377);
   U5804 : NAND4_X1 port map( A1 => n3388, A2 => n3389, A3 => n3390, A4 => 
                           n3391, ZN => n3378);
   U5805 : NAND4_X1 port map( A1 => n3380, A2 => n3381, A3 => n3382, A4 => 
                           n3383, ZN => n3379);
   U5806 : OAI21_X1 port map( B1 => n7260, B2 => n12334, A => n3358, ZN => 
                           n4919);
   U5807 : OAI21_X1 port map( B1 => n3359, B2 => n3360, A => n12343, ZN => 
                           n3358);
   U5808 : NAND4_X1 port map( A1 => n3369, A2 => n3370, A3 => n3371, A4 => 
                           n3372, ZN => n3359);
   U5809 : NAND4_X1 port map( A1 => n3361, A2 => n3362, A3 => n3363, A4 => 
                           n3364, ZN => n3360);
   U5810 : OAI21_X1 port map( B1 => n7243, B2 => n12334, A => n3339, ZN => 
                           n4920);
   U5811 : OAI21_X1 port map( B1 => n3340, B2 => n3341, A => n12343, ZN => 
                           n3339);
   U5812 : NAND4_X1 port map( A1 => n3350, A2 => n3351, A3 => n3352, A4 => 
                           n3353, ZN => n3340);
   U5813 : NAND4_X1 port map( A1 => n3342, A2 => n3343, A3 => n3344, A4 => 
                           n3345, ZN => n3341);
   U5814 : OAI21_X1 port map( B1 => n7146, B2 => n12334, A => n3320, ZN => 
                           n4921);
   U5815 : OAI21_X1 port map( B1 => n3321, B2 => n3322, A => n12344, ZN => 
                           n3320);
   U5816 : NAND4_X1 port map( A1 => n3331, A2 => n3332, A3 => n3333, A4 => 
                           n3334, ZN => n3321);
   U5817 : NAND4_X1 port map( A1 => n3323, A2 => n3324, A3 => n3325, A4 => 
                           n3326, ZN => n3322);
   U5818 : OAI21_X1 port map( B1 => n7129, B2 => n12334, A => n3301, ZN => 
                           n4922);
   U5819 : OAI21_X1 port map( B1 => n3302, B2 => n3303, A => n12344, ZN => 
                           n3301);
   U5820 : NAND4_X1 port map( A1 => n3304, A2 => n3305, A3 => n3306, A4 => 
                           n3307, ZN => n3303);
   U5821 : NAND4_X1 port map( A1 => n3312, A2 => n3313, A3 => n3314, A4 => 
                           n3315, ZN => n3302);
   U5822 : OAI21_X1 port map( B1 => n7112, B2 => n12334, A => n3282, ZN => 
                           n4923);
   U5823 : OAI21_X1 port map( B1 => n3283, B2 => n3284, A => n12344, ZN => 
                           n3282);
   U5824 : NAND4_X1 port map( A1 => n3285, A2 => n3286, A3 => n3287, A4 => 
                           n3288, ZN => n3284);
   U5825 : NAND4_X1 port map( A1 => n3293, A2 => n3294, A3 => n3295, A4 => 
                           n3296, ZN => n3283);
   U5826 : OAI21_X1 port map( B1 => n4851, B2 => n12334, A => n3263, ZN => 
                           n4924);
   U5827 : OAI21_X1 port map( B1 => n3264, B2 => n3265, A => n12344, ZN => 
                           n3263);
   U5828 : NAND4_X1 port map( A1 => n3266, A2 => n3267, A3 => n3268, A4 => 
                           n3269, ZN => n3265);
   U5829 : NAND4_X1 port map( A1 => n3274, A2 => n3275, A3 => n3276, A4 => 
                           n3277, ZN => n3264);
   U5830 : OAI21_X1 port map( B1 => n4834, B2 => n12336, A => n3212, ZN => 
                           n4925);
   U5831 : OAI21_X1 port map( B1 => n3213, B2 => n3214, A => n12344, ZN => 
                           n3212);
   U5832 : NAND4_X1 port map( A1 => n3215, A2 => n3216, A3 => n3217, A4 => 
                           n3218, ZN => n3214);
   U5833 : NAND4_X1 port map( A1 => n3239, A2 => n3240, A3 => n3241, A4 => 
                           n3242, ZN => n3213);
   U5834 : INV_X1 port map( A => ADD_RD2(1), ZN => n13390);
   U5835 : INV_X1 port map( A => ADD_RD2(2), ZN => n13389);
   U5836 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n12134, ZN => n1876);
   U5837 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n12134, ZN => n1875);
   U5838 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n12134, ZN => n1874);
   U5839 : NAND2_X1 port map( A1 => DATAIN(32), A2 => n12134, ZN => n1873);
   U5840 : NAND2_X1 port map( A1 => DATAIN(33), A2 => n12134, ZN => n1872);
   U5841 : NAND2_X1 port map( A1 => DATAIN(34), A2 => n12134, ZN => n1871);
   U5842 : NAND2_X1 port map( A1 => DATAIN(35), A2 => n12134, ZN => n1870);
   U5843 : NAND2_X1 port map( A1 => DATAIN(36), A2 => n12134, ZN => n1869);
   U5844 : NAND2_X1 port map( A1 => DATAIN(37), A2 => n12134, ZN => n1868);
   U5845 : NAND2_X1 port map( A1 => DATAIN(38), A2 => n12134, ZN => n1867);
   U5846 : NAND2_X1 port map( A1 => DATAIN(39), A2 => n12134, ZN => n1866);
   U5847 : NAND2_X1 port map( A1 => DATAIN(40), A2 => n12133, ZN => n1865);
   U5848 : NAND2_X1 port map( A1 => DATAIN(41), A2 => n12133, ZN => n1864);
   U5849 : NAND2_X1 port map( A1 => DATAIN(42), A2 => n12133, ZN => n1863);
   U5850 : NAND2_X1 port map( A1 => DATAIN(43), A2 => n12133, ZN => n1862);
   U5851 : NAND2_X1 port map( A1 => DATAIN(44), A2 => n12133, ZN => n1861);
   U5852 : NAND2_X1 port map( A1 => DATAIN(45), A2 => n12133, ZN => n1860);
   U5853 : NAND2_X1 port map( A1 => DATAIN(55), A2 => n12132, ZN => n1850);
   U5854 : NAND2_X1 port map( A1 => DATAIN(56), A2 => n12132, ZN => n1849);
   U5855 : NAND2_X1 port map( A1 => DATAIN(57), A2 => n12132, ZN => n1848);
   U5856 : NAND2_X1 port map( A1 => DATAIN(58), A2 => n12132, ZN => n1847);
   U5857 : NAND2_X1 port map( A1 => DATAIN(59), A2 => n12132, ZN => n1846);
   U5858 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n12137, ZN => n1905);
   U5859 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n12137, ZN => n1904);
   U5860 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n12137, ZN => n1903);
   U5861 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n12136, ZN => n1902);
   U5862 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n12137, ZN => n1901);
   U5863 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n12136, ZN => n1900);
   U5864 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n12136, ZN => n1899);
   U5865 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n12136, ZN => n1898);
   U5866 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n12136, ZN => n1897);
   U5867 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n12136, ZN => n1896);
   U5868 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n12136, ZN => n1895);
   U5869 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n12136, ZN => n1894);
   U5870 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n12136, ZN => n1893);
   U5871 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n12136, ZN => n1892);
   U5872 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n12136, ZN => n1891);
   U5873 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n12135, ZN => n1890);
   U5874 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n12136, ZN => n1889);
   U5875 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n12135, ZN => n1888);
   U5876 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n12135, ZN => n1887);
   U5877 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n12135, ZN => n1886);
   U5878 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n12135, ZN => n1885);
   U5879 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n12134, ZN => n1884);
   U5880 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n12135, ZN => n1883);
   U5881 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n12135, ZN => n1882);
   U5882 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n12135, ZN => n1881);
   U5883 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n12135, ZN => n1880);
   U5884 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n12135, ZN => n1879);
   U5885 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n12135, ZN => n1878);
   U5886 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n12135, ZN => n1877);
   U5887 : NAND2_X1 port map( A1 => DATAIN(46), A2 => n12133, ZN => n1859);
   U5888 : NAND2_X1 port map( A1 => DATAIN(47), A2 => n12133, ZN => n1858);
   U5889 : NAND2_X1 port map( A1 => DATAIN(48), A2 => n12133, ZN => n1857);
   U5890 : NAND2_X1 port map( A1 => DATAIN(49), A2 => n12133, ZN => n1856);
   U5891 : NAND2_X1 port map( A1 => DATAIN(50), A2 => n12133, ZN => n1855);
   U5892 : NAND2_X1 port map( A1 => DATAIN(51), A2 => n12133, ZN => n1854);
   U5893 : NAND2_X1 port map( A1 => DATAIN(52), A2 => n12132, ZN => n1853);
   U5894 : NAND2_X1 port map( A1 => DATAIN(53), A2 => n12132, ZN => n1852);
   U5895 : NAND2_X1 port map( A1 => DATAIN(54), A2 => n12132, ZN => n1851);
   U5896 : NAND2_X1 port map( A1 => DATAIN(60), A2 => n12132, ZN => n1845);
   U5897 : NAND2_X1 port map( A1 => DATAIN(61), A2 => n12132, ZN => n1844);
   U5898 : NAND2_X1 port map( A1 => DATAIN(62), A2 => n12132, ZN => n1843);
   U5899 : AND3_X1 port map( A1 => ENABLE, A2 => n12139, A3 => RD1, ZN => n1950
                           );
   U5900 : INV_X1 port map( A => RESET, ZN => n14466);
   U5901 : OAI22_X1 port map( A1 => n13027, A2 => n13170, B1 => n8574, B2 => 
                           n1923, ZN => n6462);
   U5902 : OAI22_X1 port map( A1 => n13027, A2 => n13173, B1 => n8557, B2 => 
                           n1923, ZN => n6463);
   U5903 : OAI22_X1 port map( A1 => n13027, A2 => n13176, B1 => n8540, B2 => 
                           n1923, ZN => n6464);
   U5904 : OAI22_X1 port map( A1 => n13027, A2 => n13179, B1 => n8523, B2 => 
                           n1923, ZN => n6465);
   U5905 : OAI22_X1 port map( A1 => n13026, A2 => n13182, B1 => n8506, B2 => 
                           n1923, ZN => n6466);
   U5906 : OAI22_X1 port map( A1 => n13026, A2 => n13185, B1 => n8489, B2 => 
                           n1923, ZN => n6467);
   U5907 : OAI22_X1 port map( A1 => n13026, A2 => n13188, B1 => n8472, B2 => 
                           n13010, ZN => n6468);
   U5908 : OAI22_X1 port map( A1 => n13026, A2 => n13191, B1 => n8455, B2 => 
                           n13014, ZN => n6469);
   U5909 : OAI22_X1 port map( A1 => n13026, A2 => n13194, B1 => n8438, B2 => 
                           n13013, ZN => n6470);
   U5910 : OAI22_X1 port map( A1 => n13025, A2 => n13197, B1 => n8421, B2 => 
                           n13011, ZN => n6471);
   U5911 : OAI22_X1 port map( A1 => n13025, A2 => n13200, B1 => n8404, B2 => 
                           n13014, ZN => n6472);
   U5912 : OAI22_X1 port map( A1 => n13025, A2 => n13203, B1 => n8387, B2 => 
                           n13013, ZN => n6473);
   U5913 : OAI22_X1 port map( A1 => n12945, A2 => n13207, B1 => n8372, B2 => 
                           n12931, ZN => n6218);
   U5914 : OAI22_X1 port map( A1 => n12943, A2 => n13240, B1 => n8185, B2 => 
                           n12931, ZN => n6229);
   U5915 : OAI22_X1 port map( A1 => n12943, A2 => n13237, B1 => n8202, B2 => 
                           n12931, ZN => n6228);
   U5916 : OAI22_X1 port map( A1 => n12943, A2 => n13234, B1 => n8219, B2 => 
                           n12931, ZN => n6227);
   U5917 : OAI22_X1 port map( A1 => n12943, A2 => n13231, B1 => n8236, B2 => 
                           n12931, ZN => n6226);
   U5918 : OAI22_X1 port map( A1 => n12943, A2 => n13228, B1 => n8253, B2 => 
                           n12931, ZN => n6225);
   U5919 : OAI22_X1 port map( A1 => n13047, A2 => n13170, B1 => n8572, B2 => 
                           n1920, ZN => n6526);
   U5920 : OAI22_X1 port map( A1 => n13047, A2 => n13173, B1 => n8555, B2 => 
                           n1920, ZN => n6527);
   U5921 : OAI22_X1 port map( A1 => n13047, A2 => n13176, B1 => n8538, B2 => 
                           n1920, ZN => n6528);
   U5922 : OAI22_X1 port map( A1 => n13047, A2 => n13179, B1 => n8521, B2 => 
                           n1920, ZN => n6529);
   U5923 : OAI22_X1 port map( A1 => n13046, A2 => n13182, B1 => n8504, B2 => 
                           n1920, ZN => n6530);
   U5924 : OAI22_X1 port map( A1 => n13046, A2 => n13185, B1 => n8487, B2 => 
                           n1920, ZN => n6531);
   U5925 : OAI22_X1 port map( A1 => n13046, A2 => n13188, B1 => n8470, B2 => 
                           n13030, ZN => n6532);
   U5926 : OAI22_X1 port map( A1 => n13046, A2 => n13191, B1 => n8453, B2 => 
                           n13034, ZN => n6533);
   U5927 : OAI22_X1 port map( A1 => n13046, A2 => n13194, B1 => n8436, B2 => 
                           n13033, ZN => n6534);
   U5928 : OAI22_X1 port map( A1 => n13045, A2 => n13197, B1 => n8419, B2 => 
                           n13031, ZN => n6535);
   U5929 : OAI22_X1 port map( A1 => n13045, A2 => n13200, B1 => n8402, B2 => 
                           n13034, ZN => n6536);
   U5930 : OAI22_X1 port map( A1 => n13045, A2 => n13203, B1 => n8385, B2 => 
                           n13033, ZN => n6537);
   U5931 : OAI22_X1 port map( A1 => n13067, A2 => n13170, B1 => n8571, B2 => 
                           n1918, ZN => n6590);
   U5932 : OAI22_X1 port map( A1 => n13067, A2 => n13176, B1 => n8537, B2 => 
                           n1918, ZN => n6592);
   U5933 : OAI22_X1 port map( A1 => n13067, A2 => n13179, B1 => n8520, B2 => 
                           n1918, ZN => n6593);
   U5934 : OAI22_X1 port map( A1 => n13066, A2 => n13182, B1 => n8503, B2 => 
                           n1918, ZN => n6594);
   U5935 : OAI22_X1 port map( A1 => n13066, A2 => n13185, B1 => n8486, B2 => 
                           n1918, ZN => n6595);
   U5936 : OAI22_X1 port map( A1 => n13066, A2 => n13188, B1 => n8469, B2 => 
                           n1918, ZN => n6596);
   U5937 : OAI22_X1 port map( A1 => n13066, A2 => n13191, B1 => n8452, B2 => 
                           n13050, ZN => n6597);
   U5938 : OAI22_X1 port map( A1 => n13066, A2 => n13194, B1 => n8435, B2 => 
                           n13054, ZN => n6598);
   U5939 : OAI22_X1 port map( A1 => n13065, A2 => n13197, B1 => n8418, B2 => 
                           n13053, ZN => n6599);
   U5940 : OAI22_X1 port map( A1 => n13065, A2 => n13200, B1 => n8401, B2 => 
                           n13051, ZN => n6600);
   U5941 : OAI22_X1 port map( A1 => n13065, A2 => n13203, B1 => n8384, B2 => 
                           n13054, ZN => n6601);
   U5942 : OAI22_X1 port map( A1 => n13067, A2 => n13173, B1 => n8554, B2 => 
                           n13053, ZN => n6591);
   U5943 : OAI21_X1 port map( B1 => n1909, B2 => n1924, A => n12139, ZN => 
                           n1925);
   U5944 : OAI21_X1 port map( B1 => n1907, B2 => n1924, A => n12139, ZN => 
                           n1923);
   U5945 : OAI21_X1 port map( B1 => n1915, B2 => n1924, A => n12138, ZN => 
                           n1928);
   U5946 : OAI22_X1 port map( A1 => n12945, A2 => n13204, B1 => n8389, B2 => 
                           n1928, ZN => n6217);
   U5947 : OAI22_X1 port map( A1 => n12945, A2 => n13201, B1 => n8406, B2 => 
                           n1928, ZN => n6216);
   U5948 : OAI22_X1 port map( A1 => n12945, A2 => n13198, B1 => n8423, B2 => 
                           n1928, ZN => n6215);
   U5949 : OAI22_X1 port map( A1 => n12946, A2 => n13195, B1 => n8440, B2 => 
                           n1928, ZN => n6214);
   U5950 : OAI22_X1 port map( A1 => n12946, A2 => n13192, B1 => n8457, B2 => 
                           n1928, ZN => n6213);
   U5951 : OAI22_X1 port map( A1 => n12946, A2 => n13189, B1 => n8474, B2 => 
                           n1928, ZN => n6212);
   U5952 : AND2_X1 port map( A1 => n3194, A2 => n3204, ZN => n1987);
   U5953 : AND2_X1 port map( A1 => n3191, A2 => n3204, ZN => n1982);
   U5954 : NAND2_X1 port map( A1 => n3193, A2 => n3204, ZN => n1991);
   U5955 : NAND2_X1 port map( A1 => n3189, A2 => n3204, ZN => n1986);
   U5956 : NAND3_X2 port map( A1 => ADD_WR(3), A2 => n1922, A3 => ADD_WR(4), ZN
                           => n1942);
   U5957 : OAI22_X1 port map( A1 => n12867, A2 => n13171, B1 => n8578, B2 => 
                           n1932, ZN => n5950);
   U5958 : OAI22_X1 port map( A1 => n12867, A2 => n13174, B1 => n8561, B2 => 
                           n1932, ZN => n5951);
   U5959 : OAI22_X1 port map( A1 => n12867, A2 => n13177, B1 => n8544, B2 => 
                           n1932, ZN => n5952);
   U5960 : OAI22_X1 port map( A1 => n12867, A2 => n13180, B1 => n8527, B2 => 
                           n1932, ZN => n5953);
   U5961 : OAI22_X1 port map( A1 => n12866, A2 => n13183, B1 => n8510, B2 => 
                           n1932, ZN => n5954);
   U5962 : OAI22_X1 port map( A1 => n12866, A2 => n13186, B1 => n8493, B2 => 
                           n1932, ZN => n5955);
   U5963 : OAI22_X1 port map( A1 => n12866, A2 => n13189, B1 => n8476, B2 => 
                           n12850, ZN => n5956);
   U5964 : OAI22_X1 port map( A1 => n12866, A2 => n13192, B1 => n8459, B2 => 
                           n12854, ZN => n5957);
   U5965 : OAI22_X1 port map( A1 => n12866, A2 => n13195, B1 => n8442, B2 => 
                           n12853, ZN => n5958);
   U5966 : OAI22_X1 port map( A1 => n12865, A2 => n13198, B1 => n8425, B2 => 
                           n12851, ZN => n5959);
   U5967 : OAI22_X1 port map( A1 => n12865, A2 => n13201, B1 => n8408, B2 => 
                           n12854, ZN => n5960);
   U5968 : OAI22_X1 port map( A1 => n12865, A2 => n13204, B1 => n8391, B2 => 
                           n12853, ZN => n5961);
   U5969 : OAI21_X1 port map( B1 => n1911, B2 => n1933, A => n12138, ZN => 
                           n1935);
   U5970 : OAI21_X1 port map( B1 => n1913, B2 => n1933, A => n12138, ZN => 
                           n1936);
   U5971 : OAI21_X1 port map( B1 => n1919, B2 => n1933, A => n12138, ZN => 
                           n1939);
   U5972 : OAI21_X1 port map( B1 => n1921, B2 => n1933, A => n12138, ZN => 
                           n1940);
   U5973 : OAI21_X1 port map( B1 => n1909, B2 => n1933, A => n12138, ZN => 
                           n1934);
   U5974 : OAI21_X1 port map( B1 => n1915, B2 => n1933, A => n12138, ZN => 
                           n1937);
   U5975 : OAI21_X1 port map( B1 => n1917, B2 => n1933, A => n12138, ZN => 
                           n1938);
   U5976 : OAI21_X1 port map( B1 => n1907, B2 => n1933, A => n12138, ZN => 
                           n1932);
   U5977 : OAI22_X1 port map( A1 => n13127, A2 => n13170, B1 => n8570, B2 => 
                           n1912, ZN => n6782);
   U5978 : OAI22_X1 port map( A1 => n13127, A2 => n13173, B1 => n8553, B2 => 
                           n1912, ZN => n6783);
   U5979 : OAI22_X1 port map( A1 => n13127, A2 => n13176, B1 => n8536, B2 => 
                           n1912, ZN => n6784);
   U5980 : OAI22_X1 port map( A1 => n13127, A2 => n13179, B1 => n8519, B2 => 
                           n1912, ZN => n6785);
   U5981 : OAI22_X1 port map( A1 => n13126, A2 => n13182, B1 => n8502, B2 => 
                           n1912, ZN => n6786);
   U5982 : OAI22_X1 port map( A1 => n13126, A2 => n13185, B1 => n8485, B2 => 
                           n1912, ZN => n6787);
   U5983 : OAI22_X1 port map( A1 => n13126, A2 => n13188, B1 => n8468, B2 => 
                           n1912, ZN => n6788);
   U5984 : OAI22_X1 port map( A1 => n13126, A2 => n13191, B1 => n8451, B2 => 
                           n1912, ZN => n6789);
   U5985 : OAI22_X1 port map( A1 => n13126, A2 => n13194, B1 => n8434, B2 => 
                           n13110, ZN => n6790);
   U5986 : OAI22_X1 port map( A1 => n13125, A2 => n13197, B1 => n8417, B2 => 
                           n13111, ZN => n6791);
   U5987 : OAI22_X1 port map( A1 => n13125, A2 => n13200, B1 => n8400, B2 => 
                           n13114, ZN => n6792);
   U5988 : OAI22_X1 port map( A1 => n13125, A2 => n13203, B1 => n8383, B2 => 
                           n13113, ZN => n6793);
   U5989 : OAI21_X1 port map( B1 => n1906, B2 => n1907, A => n12137, ZN => 
                           n1842);
   U5990 : OAI21_X1 port map( B1 => n1906, B2 => n1909, A => n12139, ZN => 
                           n1908);
   U5991 : OAI21_X1 port map( B1 => n1906, B2 => n1911, A => n12139, ZN => 
                           n1910);
   U5992 : OAI21_X1 port map( B1 => n1906, B2 => n1915, A => n12139, ZN => 
                           n1914);
   U5993 : OAI21_X1 port map( B1 => n1906, B2 => n1917, A => n12139, ZN => 
                           n1916);
   U5994 : OAI21_X1 port map( B1 => n1906, B2 => n1919, A => n12139, ZN => 
                           n1918);
   U5995 : OAI21_X1 port map( B1 => n1906, B2 => n1921, A => n12139, ZN => 
                           n1920);
   U5996 : OAI21_X1 port map( B1 => n1906, B2 => n1913, A => n12139, ZN => 
                           n1912);
   U5997 : INV_X1 port map( A => ADD_WR(4), ZN => n13382);
   U5998 : NAND3_X2 port map( A1 => n1922, A2 => n13382, A3 => ADD_WR(3), ZN =>
                           n1924);
   U5999 : CLKBUF_X1 port map( A => n14466, Z => n12129);
   U6000 : CLKBUF_X1 port map( A => n14466, Z => n12130);
   U6001 : CLKBUF_X1 port map( A => n14466, Z => n12131);
   U6002 : CLKBUF_X1 port map( A => n3262, Z => n12145);
   U6003 : CLKBUF_X1 port map( A => n3261, Z => n12151);
   U6004 : CLKBUF_X1 port map( A => n3259, Z => n12157);
   U6005 : CLKBUF_X1 port map( A => n3258, Z => n12163);
   U6006 : CLKBUF_X1 port map( A => n3257, Z => n12169);
   U6007 : CLKBUF_X1 port map( A => n3256, Z => n12175);
   U6008 : CLKBUF_X1 port map( A => n3254, Z => n12181);
   U6009 : CLKBUF_X1 port map( A => n3253, Z => n12187);
   U6010 : CLKBUF_X1 port map( A => n3252, Z => n12193);
   U6011 : CLKBUF_X1 port map( A => n3251, Z => n12199);
   U6012 : CLKBUF_X1 port map( A => n3249, Z => n12205);
   U6013 : CLKBUF_X1 port map( A => n3248, Z => n12211);
   U6014 : CLKBUF_X1 port map( A => n3247, Z => n12217);
   U6015 : CLKBUF_X1 port map( A => n3246, Z => n12223);
   U6016 : CLKBUF_X1 port map( A => n3244, Z => n12229);
   U6017 : CLKBUF_X1 port map( A => n3243, Z => n12235);
   U6018 : CLKBUF_X1 port map( A => n3238, Z => n12241);
   U6019 : CLKBUF_X1 port map( A => n3237, Z => n12247);
   U6020 : CLKBUF_X1 port map( A => n3235, Z => n12253);
   U6021 : CLKBUF_X1 port map( A => n3234, Z => n12259);
   U6022 : CLKBUF_X1 port map( A => n3233, Z => n12265);
   U6023 : CLKBUF_X1 port map( A => n3232, Z => n12271);
   U6024 : CLKBUF_X1 port map( A => n3230, Z => n12277);
   U6025 : CLKBUF_X1 port map( A => n3229, Z => n12283);
   U6026 : CLKBUF_X1 port map( A => n3228, Z => n12289);
   U6027 : CLKBUF_X1 port map( A => n3227, Z => n12295);
   U6028 : CLKBUF_X1 port map( A => n3225, Z => n12301);
   U6029 : CLKBUF_X1 port map( A => n3224, Z => n12307);
   U6030 : CLKBUF_X1 port map( A => n3223, Z => n12313);
   U6031 : CLKBUF_X1 port map( A => n3222, Z => n12319);
   U6032 : CLKBUF_X1 port map( A => n3220, Z => n12325);
   U6033 : CLKBUF_X1 port map( A => n3219, Z => n12331);
   U6034 : CLKBUF_X1 port map( A => n12333, Z => n12344);
   U6035 : CLKBUF_X1 port map( A => n2001, Z => n12350);
   U6036 : CLKBUF_X1 port map( A => n2000, Z => n12356);
   U6037 : CLKBUF_X1 port map( A => n1998, Z => n12362);
   U6038 : CLKBUF_X1 port map( A => n1997, Z => n12368);
   U6039 : CLKBUF_X1 port map( A => n1996, Z => n12374);
   U6040 : CLKBUF_X1 port map( A => n1995, Z => n12380);
   U6041 : CLKBUF_X1 port map( A => n1993, Z => n12386);
   U6042 : CLKBUF_X1 port map( A => n1992, Z => n12392);
   U6043 : CLKBUF_X1 port map( A => n1991, Z => n12398);
   U6044 : CLKBUF_X1 port map( A => n1990, Z => n12404);
   U6045 : CLKBUF_X1 port map( A => n1988, Z => n12410);
   U6046 : CLKBUF_X1 port map( A => n1987, Z => n12416);
   U6047 : CLKBUF_X1 port map( A => n1986, Z => n12422);
   U6048 : CLKBUF_X1 port map( A => n1985, Z => n12428);
   U6049 : CLKBUF_X1 port map( A => n1983, Z => n12434);
   U6050 : CLKBUF_X1 port map( A => n1982, Z => n12440);
   U6051 : CLKBUF_X1 port map( A => n1977, Z => n12446);
   U6052 : CLKBUF_X1 port map( A => n1976, Z => n12452);
   U6053 : CLKBUF_X1 port map( A => n1974, Z => n12458);
   U6054 : CLKBUF_X1 port map( A => n1973, Z => n12464);
   U6055 : CLKBUF_X1 port map( A => n1972, Z => n12470);
   U6056 : CLKBUF_X1 port map( A => n1971, Z => n12476);
   U6057 : CLKBUF_X1 port map( A => n1969, Z => n12482);
   U6058 : CLKBUF_X1 port map( A => n1968, Z => n12488);
   U6059 : CLKBUF_X1 port map( A => n1967, Z => n12494);
   U6060 : CLKBUF_X1 port map( A => n1966, Z => n12500);
   U6061 : CLKBUF_X1 port map( A => n1964, Z => n12506);
   U6062 : CLKBUF_X1 port map( A => n1963, Z => n12512);
   U6063 : CLKBUF_X1 port map( A => n1962, Z => n12518);
   U6064 : CLKBUF_X1 port map( A => n1961, Z => n12524);
   U6065 : CLKBUF_X1 port map( A => n1959, Z => n12530);
   U6066 : CLKBUF_X1 port map( A => n1958, Z => n12536);
   U6067 : CLKBUF_X1 port map( A => n12538, Z => n12549);
   U6068 : INV_X1 port map( A => n12573, ZN => n12556);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_M8_N4_N_bit64_W2.all;

entity windowed_register_file_M8_N4_N_bit64_W2 is

   port( CALL, RETURN_signal, CLK, RESET, ENABLE, RD_CPU, WR_CPU : in std_logic
         ;  Wait_signal : out std_logic;  ADDR_WRCPU, ADDR_RDCPU : in 
         std_logic_vector (4 downto 0);  DATAIN_CPU : in std_logic_vector (63 
         downto 0);  DATAOUT_CPU : out std_logic_vector (63 downto 0);  
         RD_WR_MEM : out std_logic;  DATAIN_MEM : in std_logic_vector (63 
         downto 0);  DATAOUT_MEM : out std_logic_vector (63 downto 0));

end windowed_register_file_M8_N4_N_bit64_W2;

architecture SYN_structural of windowed_register_file_M8_N4_N_bit64_W2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFRS_X1
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_3
      port( A : in std_logic_vector (31 downto 0);  INC_DEC : in std_logic;  
            SUM : out std_logic_vector (31 downto 0));
   end component;
   
   component windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_2
      port( A : in std_logic_vector (31 downto 0);  INC_DEC : in std_logic;  
            SUM : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_generic_N64
      port( A, B : in std_logic_vector (63 downto 0);  sel : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component address_conversion_M8_N4_N_bit64_F3
      port( spill_fill_count : in std_logic;  wait_count, start_write : out 
            std_logic;  clck : in std_logic;  address_input_1, address_input_3 
            : in std_logic_vector (4 downto 0);  address_output_1, 
            address_output_2, address_output_3 : out std_logic_vector (4 downto
            0);  swp, cwp : in std_logic_vector (4 downto 0));
   end component;
   
   component register_file_NBIT64_NREG32
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal full, count_wait, RD_MEM, ADDRESS_WRITE_4_port, ADDRESS_WRITE_3_port,
      ADDRESS_WRITE_2_port, ADDRESS_WRITE_1_port, ADDRESS_WRITE_0_port, 
      ADDRESS_READ_4_port, ADDRESS_READ_3_port, ADDRESS_READ_2_port, 
      ADDRESS_READ_1_port, ADDRESS_READ_0_port, ADDRESS_COUNT_4_port, 
      ADDRESS_COUNT_3_port, ADDRESS_COUNT_2_port, ADDRESS_COUNT_1_port, 
      ADDRESS_COUNT_0_port, DATA_WRITE_63_port, DATA_WRITE_62_port, 
      DATA_WRITE_61_port, DATA_WRITE_60_port, DATA_WRITE_59_port, 
      DATA_WRITE_58_port, DATA_WRITE_57_port, DATA_WRITE_56_port, 
      DATA_WRITE_55_port, DATA_WRITE_54_port, DATA_WRITE_53_port, 
      DATA_WRITE_52_port, DATA_WRITE_51_port, DATA_WRITE_50_port, 
      DATA_WRITE_49_port, DATA_WRITE_48_port, DATA_WRITE_47_port, 
      DATA_WRITE_46_port, DATA_WRITE_45_port, DATA_WRITE_44_port, 
      DATA_WRITE_43_port, DATA_WRITE_42_port, DATA_WRITE_41_port, 
      DATA_WRITE_40_port, DATA_WRITE_39_port, DATA_WRITE_38_port, 
      DATA_WRITE_37_port, DATA_WRITE_36_port, DATA_WRITE_35_port, 
      DATA_WRITE_34_port, DATA_WRITE_33_port, DATA_WRITE_32_port, 
      DATA_WRITE_31_port, DATA_WRITE_30_port, DATA_WRITE_29_port, 
      DATA_WRITE_28_port, DATA_WRITE_27_port, DATA_WRITE_26_port, 
      DATA_WRITE_25_port, DATA_WRITE_24_port, DATA_WRITE_23_port, 
      DATA_WRITE_22_port, DATA_WRITE_21_port, DATA_WRITE_20_port, 
      DATA_WRITE_19_port, DATA_WRITE_18_port, DATA_WRITE_17_port, 
      DATA_WRITE_16_port, DATA_WRITE_15_port, DATA_WRITE_14_port, 
      DATA_WRITE_13_port, DATA_WRITE_12_port, DATA_WRITE_11_port, 
      DATA_WRITE_10_port, DATA_WRITE_9_port, DATA_WRITE_8_port, 
      DATA_WRITE_7_port, DATA_WRITE_6_port, DATA_WRITE_5_port, 
      DATA_WRITE_4_port, DATA_WRITE_3_port, DATA_WRITE_2_port, 
      DATA_WRITE_1_port, DATA_WRITE_0_port, start, swp_4_port, swp_3_port, 
      cwp_4_port, cwp_3_port, cwp_0_port, canrestore_31_port, 
      canrestore_30_port, canrestore_29_port, canrestore_28_port, 
      canrestore_27_port, canrestore_26_port, canrestore_25_port, 
      canrestore_24_port, canrestore_23_port, canrestore_22_port, 
      canrestore_21_port, canrestore_20_port, canrestore_19_port, 
      canrestore_18_port, canrestore_17_port, canrestore_16_port, 
      canrestore_15_port, canrestore_14_port, canrestore_13_port, 
      canrestore_12_port, canrestore_11_port, canrestore_10_port, 
      canrestore_9_port, canrestore_8_port, canrestore_7_port, 
      canrestore_6_port, canrestore_5_port, canrestore_4_port, 
      canrestore_3_port, canrestore_2_port, canrestore_1_port, 
      canrestore_0_port, cansave_31_port, cansave_30_port, cansave_29_port, 
      cansave_28_port, cansave_27_port, cansave_26_port, cansave_25_port, 
      cansave_24_port, cansave_23_port, cansave_22_port, cansave_21_port, 
      cansave_20_port, cansave_19_port, cansave_18_port, cansave_17_port, 
      cansave_16_port, cansave_15_port, cansave_14_port, cansave_13_port, 
      cansave_12_port, cansave_11_port, cansave_10_port, cansave_9_port, 
      cansave_8_port, cansave_7_port, cansave_6_port, cansave_5_port, 
      cansave_4_port, cansave_3_port, cansave_2_port, cansave_1_port, 
      cansave_0_port, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, 
      N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79
      , N80, N81, N82, N83, N84, N212, N213, N264, N265, N266, N267, N268, N269
      , N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
      N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, 
      N294, N295, N351, N352, N353, n156, n157, n158, n159, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n196, n197, n198, n200, n202, n204, 
      n205, n206, n208, n209, n210, n211, n212_port, n213_port, n214, n215, 
      n216, n248, n282_port, n283_port, n290_port, n387, n389, n390, n392, n393
      , n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
      n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, 
      n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n431, 
      n565, n566, n567, n568, n570, n571, n572, n573, n576, n577, n578, n579, 
      n581, n582, n583, n588, n589, n621, n675, n724, n725, n726, n727, n728, 
      n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, 
      n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, 
      n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, 
      n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, 
      n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, 
      n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, 
      n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, 
      n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      Wait_signal_port, n825, n826, n827, n828, n829, n830, n831, n832, n833, 
      n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, 
      n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, RD_WR_MEM_port, n912, n_2070, n_2071 : std_logic;

begin
   Wait_signal <= Wait_signal_port;
   RD_WR_MEM <= RD_WR_MEM_port;
   
   canrestore_reg_28_inst : DFF_X1 port map( D => n409, CK => CLK, Q => 
                           canrestore_28_port, QN => n815);
   canrestore_reg_29_inst : DFF_X1 port map( D => n408, CK => CLK, Q => 
                           canrestore_29_port, QN => n814);
   canrestore_reg_26_inst : DFF_X1 port map( D => n411, CK => CLK, Q => 
                           canrestore_26_port, QN => n588);
   canrestore_reg_27_inst : DFF_X1 port map( D => n410, CK => CLK, Q => 
                           canrestore_27_port, QN => n573);
   canrestore_reg_30_inst : DFF_X1 port map( D => n406, CK => CLK, Q => 
                           canrestore_30_port, QN => n813);
   canrestore_reg_31_inst : DFF_X1 port map( D => n405, CK => CLK, Q => 
                           canrestore_31_port, QN => n389);
   U667 : XOR2_X1 port map( A => n197, B => n725, Z => n772);
   U668 : NAND3_X1 port map( A1 => n775, A2 => cansave_0_port, A3 => n776, ZN 
                           => n773);
   U669 : XOR2_X1 port map( A => cansave_1_port, B => CALL, Z => n776);
   U670 : NAND3_X1 port map( A1 => n731, A2 => n771, A3 => n780, ZN => n779);
   U671 : XOR2_X1 port map( A => n193, B => n157, Z => n787);
   U672 : XOR2_X1 port map( A => n192, B => n158, Z => n785);
   U673 : XOR2_X1 port map( A => swp_4_port, B => n788, Z => n783);
   U674 : XOR2_X1 port map( A => n621, B => cwp_3_port, Z => n789);
   U675 : NAND3_X1 port map( A1 => n872, A2 => cwp_3_port, A3 => swp_3_port, ZN
                           => n782);
   U676 : NAND3_X1 port map( A1 => n794, A2 => n795, A3 => n796, ZN => n793);
   U677 : NAND3_X1 port map( A1 => n775, A2 => cansave_0_port, A3 => n196, ZN 
                           => n731);
   U678 : NAND3_X1 port map( A1 => n775, A2 => cansave_1_port, A3 => n197, ZN 
                           => n780);
   U679 : NAND3_X1 port map( A1 => cansave_1_port, A2 => cansave_0_port, A3 => 
                           n775, ZN => n770);
   U680 : NAND3_X1 port map( A1 => n174, A2 => n173, A3 => n175, ZN => n811);
   WRF : register_file_NBIT64_NREG32 port map( CLK => CLK, RESET => RESET, 
                           ENABLE => ENABLE, RD1 => RD_CPU, RD2 => RD_MEM, WR 
                           => n875, ADD_WR(4) => ADDRESS_WRITE_4_port, 
                           ADD_WR(3) => ADDRESS_WRITE_3_port, ADD_WR(2) => 
                           ADDRESS_WRITE_2_port, ADD_WR(1) => 
                           ADDRESS_WRITE_1_port, ADD_WR(0) => 
                           ADDRESS_WRITE_0_port, ADD_RD1(4) => 
                           ADDRESS_READ_4_port, ADD_RD1(3) => 
                           ADDRESS_READ_3_port, ADD_RD1(2) => 
                           ADDRESS_READ_2_port, ADD_RD1(1) => 
                           ADDRESS_READ_1_port, ADD_RD1(0) => 
                           ADDRESS_READ_0_port, ADD_RD2(4) => 
                           ADDRESS_COUNT_4_port, ADD_RD2(3) => 
                           ADDRESS_COUNT_3_port, ADD_RD2(2) => 
                           ADDRESS_COUNT_2_port, ADD_RD2(1) => 
                           ADDRESS_COUNT_1_port, ADD_RD2(0) => 
                           ADDRESS_COUNT_0_port, DATAIN(63) => 
                           DATA_WRITE_63_port, DATAIN(62) => DATA_WRITE_62_port
                           , DATAIN(61) => DATA_WRITE_61_port, DATAIN(60) => 
                           DATA_WRITE_60_port, DATAIN(59) => DATA_WRITE_59_port
                           , DATAIN(58) => DATA_WRITE_58_port, DATAIN(57) => 
                           DATA_WRITE_57_port, DATAIN(56) => DATA_WRITE_56_port
                           , DATAIN(55) => DATA_WRITE_55_port, DATAIN(54) => 
                           DATA_WRITE_54_port, DATAIN(53) => DATA_WRITE_53_port
                           , DATAIN(52) => DATA_WRITE_52_port, DATAIN(51) => 
                           DATA_WRITE_51_port, DATAIN(50) => DATA_WRITE_50_port
                           , DATAIN(49) => DATA_WRITE_49_port, DATAIN(48) => 
                           DATA_WRITE_48_port, DATAIN(47) => DATA_WRITE_47_port
                           , DATAIN(46) => DATA_WRITE_46_port, DATAIN(45) => 
                           DATA_WRITE_45_port, DATAIN(44) => DATA_WRITE_44_port
                           , DATAIN(43) => DATA_WRITE_43_port, DATAIN(42) => 
                           DATA_WRITE_42_port, DATAIN(41) => DATA_WRITE_41_port
                           , DATAIN(40) => DATA_WRITE_40_port, DATAIN(39) => 
                           DATA_WRITE_39_port, DATAIN(38) => DATA_WRITE_38_port
                           , DATAIN(37) => DATA_WRITE_37_port, DATAIN(36) => 
                           DATA_WRITE_36_port, DATAIN(35) => DATA_WRITE_35_port
                           , DATAIN(34) => DATA_WRITE_34_port, DATAIN(33) => 
                           DATA_WRITE_33_port, DATAIN(32) => DATA_WRITE_32_port
                           , DATAIN(31) => DATA_WRITE_31_port, DATAIN(30) => 
                           DATA_WRITE_30_port, DATAIN(29) => DATA_WRITE_29_port
                           , DATAIN(28) => DATA_WRITE_28_port, DATAIN(27) => 
                           DATA_WRITE_27_port, DATAIN(26) => DATA_WRITE_26_port
                           , DATAIN(25) => DATA_WRITE_25_port, DATAIN(24) => 
                           DATA_WRITE_24_port, DATAIN(23) => DATA_WRITE_23_port
                           , DATAIN(22) => DATA_WRITE_22_port, DATAIN(21) => 
                           DATA_WRITE_21_port, DATAIN(20) => DATA_WRITE_20_port
                           , DATAIN(19) => DATA_WRITE_19_port, DATAIN(18) => 
                           DATA_WRITE_18_port, DATAIN(17) => DATA_WRITE_17_port
                           , DATAIN(16) => DATA_WRITE_16_port, DATAIN(15) => 
                           DATA_WRITE_15_port, DATAIN(14) => DATA_WRITE_14_port
                           , DATAIN(13) => DATA_WRITE_13_port, DATAIN(12) => 
                           DATA_WRITE_12_port, DATAIN(11) => DATA_WRITE_11_port
                           , DATAIN(10) => DATA_WRITE_10_port, DATAIN(9) => 
                           DATA_WRITE_9_port, DATAIN(8) => DATA_WRITE_8_port, 
                           DATAIN(7) => DATA_WRITE_7_port, DATAIN(6) => 
                           DATA_WRITE_6_port, DATAIN(5) => DATA_WRITE_5_port, 
                           DATAIN(4) => DATA_WRITE_4_port, DATAIN(3) => 
                           DATA_WRITE_3_port, DATAIN(2) => DATA_WRITE_2_port, 
                           DATAIN(1) => DATA_WRITE_1_port, DATAIN(0) => 
                           DATA_WRITE_0_port, OUT1(63) => DATAOUT_CPU(63), 
                           OUT1(62) => DATAOUT_CPU(62), OUT1(61) => 
                           DATAOUT_CPU(61), OUT1(60) => DATAOUT_CPU(60), 
                           OUT1(59) => DATAOUT_CPU(59), OUT1(58) => 
                           DATAOUT_CPU(58), OUT1(57) => DATAOUT_CPU(57), 
                           OUT1(56) => DATAOUT_CPU(56), OUT1(55) => 
                           DATAOUT_CPU(55), OUT1(54) => DATAOUT_CPU(54), 
                           OUT1(53) => DATAOUT_CPU(53), OUT1(52) => 
                           DATAOUT_CPU(52), OUT1(51) => DATAOUT_CPU(51), 
                           OUT1(50) => DATAOUT_CPU(50), OUT1(49) => 
                           DATAOUT_CPU(49), OUT1(48) => DATAOUT_CPU(48), 
                           OUT1(47) => DATAOUT_CPU(47), OUT1(46) => 
                           DATAOUT_CPU(46), OUT1(45) => DATAOUT_CPU(45), 
                           OUT1(44) => DATAOUT_CPU(44), OUT1(43) => 
                           DATAOUT_CPU(43), OUT1(42) => DATAOUT_CPU(42), 
                           OUT1(41) => DATAOUT_CPU(41), OUT1(40) => 
                           DATAOUT_CPU(40), OUT1(39) => DATAOUT_CPU(39), 
                           OUT1(38) => DATAOUT_CPU(38), OUT1(37) => 
                           DATAOUT_CPU(37), OUT1(36) => DATAOUT_CPU(36), 
                           OUT1(35) => DATAOUT_CPU(35), OUT1(34) => 
                           DATAOUT_CPU(34), OUT1(33) => DATAOUT_CPU(33), 
                           OUT1(32) => DATAOUT_CPU(32), OUT1(31) => 
                           DATAOUT_CPU(31), OUT1(30) => DATAOUT_CPU(30), 
                           OUT1(29) => DATAOUT_CPU(29), OUT1(28) => 
                           DATAOUT_CPU(28), OUT1(27) => DATAOUT_CPU(27), 
                           OUT1(26) => DATAOUT_CPU(26), OUT1(25) => 
                           DATAOUT_CPU(25), OUT1(24) => DATAOUT_CPU(24), 
                           OUT1(23) => DATAOUT_CPU(23), OUT1(22) => 
                           DATAOUT_CPU(22), OUT1(21) => DATAOUT_CPU(21), 
                           OUT1(20) => DATAOUT_CPU(20), OUT1(19) => 
                           DATAOUT_CPU(19), OUT1(18) => DATAOUT_CPU(18), 
                           OUT1(17) => DATAOUT_CPU(17), OUT1(16) => 
                           DATAOUT_CPU(16), OUT1(15) => DATAOUT_CPU(15), 
                           OUT1(14) => DATAOUT_CPU(14), OUT1(13) => 
                           DATAOUT_CPU(13), OUT1(12) => DATAOUT_CPU(12), 
                           OUT1(11) => DATAOUT_CPU(11), OUT1(10) => 
                           DATAOUT_CPU(10), OUT1(9) => DATAOUT_CPU(9), OUT1(8) 
                           => DATAOUT_CPU(8), OUT1(7) => DATAOUT_CPU(7), 
                           OUT1(6) => DATAOUT_CPU(6), OUT1(5) => DATAOUT_CPU(5)
                           , OUT1(4) => DATAOUT_CPU(4), OUT1(3) => 
                           DATAOUT_CPU(3), OUT1(2) => DATAOUT_CPU(2), OUT1(1) 
                           => DATAOUT_CPU(1), OUT1(0) => DATAOUT_CPU(0), 
                           OUT2(63) => DATAOUT_MEM(63), OUT2(62) => 
                           DATAOUT_MEM(62), OUT2(61) => DATAOUT_MEM(61), 
                           OUT2(60) => DATAOUT_MEM(60), OUT2(59) => 
                           DATAOUT_MEM(59), OUT2(58) => DATAOUT_MEM(58), 
                           OUT2(57) => DATAOUT_MEM(57), OUT2(56) => 
                           DATAOUT_MEM(56), OUT2(55) => DATAOUT_MEM(55), 
                           OUT2(54) => DATAOUT_MEM(54), OUT2(53) => 
                           DATAOUT_MEM(53), OUT2(52) => DATAOUT_MEM(52), 
                           OUT2(51) => DATAOUT_MEM(51), OUT2(50) => 
                           DATAOUT_MEM(50), OUT2(49) => DATAOUT_MEM(49), 
                           OUT2(48) => DATAOUT_MEM(48), OUT2(47) => 
                           DATAOUT_MEM(47), OUT2(46) => DATAOUT_MEM(46), 
                           OUT2(45) => DATAOUT_MEM(45), OUT2(44) => 
                           DATAOUT_MEM(44), OUT2(43) => DATAOUT_MEM(43), 
                           OUT2(42) => DATAOUT_MEM(42), OUT2(41) => 
                           DATAOUT_MEM(41), OUT2(40) => DATAOUT_MEM(40), 
                           OUT2(39) => DATAOUT_MEM(39), OUT2(38) => 
                           DATAOUT_MEM(38), OUT2(37) => DATAOUT_MEM(37), 
                           OUT2(36) => DATAOUT_MEM(36), OUT2(35) => 
                           DATAOUT_MEM(35), OUT2(34) => DATAOUT_MEM(34), 
                           OUT2(33) => DATAOUT_MEM(33), OUT2(32) => 
                           DATAOUT_MEM(32), OUT2(31) => DATAOUT_MEM(31), 
                           OUT2(30) => DATAOUT_MEM(30), OUT2(29) => 
                           DATAOUT_MEM(29), OUT2(28) => DATAOUT_MEM(28), 
                           OUT2(27) => DATAOUT_MEM(27), OUT2(26) => 
                           DATAOUT_MEM(26), OUT2(25) => DATAOUT_MEM(25), 
                           OUT2(24) => DATAOUT_MEM(24), OUT2(23) => 
                           DATAOUT_MEM(23), OUT2(22) => DATAOUT_MEM(22), 
                           OUT2(21) => DATAOUT_MEM(21), OUT2(20) => 
                           DATAOUT_MEM(20), OUT2(19) => DATAOUT_MEM(19), 
                           OUT2(18) => DATAOUT_MEM(18), OUT2(17) => 
                           DATAOUT_MEM(17), OUT2(16) => DATAOUT_MEM(16), 
                           OUT2(15) => DATAOUT_MEM(15), OUT2(14) => 
                           DATAOUT_MEM(14), OUT2(13) => DATAOUT_MEM(13), 
                           OUT2(12) => DATAOUT_MEM(12), OUT2(11) => 
                           DATAOUT_MEM(11), OUT2(10) => DATAOUT_MEM(10), 
                           OUT2(9) => DATAOUT_MEM(9), OUT2(8) => DATAOUT_MEM(8)
                           , OUT2(7) => DATAOUT_MEM(7), OUT2(6) => 
                           DATAOUT_MEM(6), OUT2(5) => DATAOUT_MEM(5), OUT2(4) 
                           => DATAOUT_MEM(4), OUT2(3) => DATAOUT_MEM(3), 
                           OUT2(2) => DATAOUT_MEM(2), OUT2(1) => DATAOUT_MEM(1)
                           , OUT2(0) => DATAOUT_MEM(0));
   add_con : address_conversion_M8_N4_N_bit64_F3 port map( spill_fill_count => 
                           full, wait_count => count_wait, start_write => start
                           , clck => CLK, address_input_1(4) => ADDR_RDCPU(4), 
                           address_input_1(3) => ADDR_RDCPU(3), 
                           address_input_1(2) => ADDR_RDCPU(2), 
                           address_input_1(1) => ADDR_RDCPU(1), 
                           address_input_1(0) => ADDR_RDCPU(0), 
                           address_input_3(4) => ADDR_WRCPU(4), 
                           address_input_3(3) => ADDR_WRCPU(3), 
                           address_input_3(2) => ADDR_WRCPU(2), 
                           address_input_3(1) => ADDR_WRCPU(1), 
                           address_input_3(0) => ADDR_WRCPU(0), 
                           address_output_1(4) => ADDRESS_READ_4_port, 
                           address_output_1(3) => ADDRESS_READ_3_port, 
                           address_output_1(2) => ADDRESS_READ_2_port, 
                           address_output_1(1) => ADDRESS_READ_1_port, 
                           address_output_1(0) => ADDRESS_READ_0_port, 
                           address_output_2(4) => ADDRESS_COUNT_4_port, 
                           address_output_2(3) => ADDRESS_COUNT_3_port, 
                           address_output_2(2) => ADDRESS_COUNT_2_port, 
                           address_output_2(1) => ADDRESS_COUNT_1_port, 
                           address_output_2(0) => ADDRESS_COUNT_0_port, 
                           address_output_3(4) => ADDRESS_WRITE_4_port, 
                           address_output_3(3) => ADDRESS_WRITE_3_port, 
                           address_output_3(2) => ADDRESS_WRITE_2_port, 
                           address_output_3(1) => ADDRESS_WRITE_1_port, 
                           address_output_3(0) => ADDRESS_WRITE_0_port, swp(4) 
                           => swp_4_port, swp(3) => swp_3_port, swp(2) => N353,
                           swp(1) => N352, swp(0) => N351, cwp(4) => cwp_4_port
                           , cwp(3) => cwp_3_port, cwp(2) => N213, cwp(1) => 
                           N212, cwp(0) => cwp_0_port);
   DATA_multiplexer_write : MUX21_generic_N64 port map( A(63) => DATAIN_MEM(63)
                           , A(62) => DATAIN_MEM(62), A(61) => DATAIN_MEM(61), 
                           A(60) => DATAIN_MEM(60), A(59) => DATAIN_MEM(59), 
                           A(58) => DATAIN_MEM(58), A(57) => DATAIN_MEM(57), 
                           A(56) => DATAIN_MEM(56), A(55) => DATAIN_MEM(55), 
                           A(54) => DATAIN_MEM(54), A(53) => DATAIN_MEM(53), 
                           A(52) => DATAIN_MEM(52), A(51) => DATAIN_MEM(51), 
                           A(50) => DATAIN_MEM(50), A(49) => DATAIN_MEM(49), 
                           A(48) => DATAIN_MEM(48), A(47) => DATAIN_MEM(47), 
                           A(46) => DATAIN_MEM(46), A(45) => DATAIN_MEM(45), 
                           A(44) => DATAIN_MEM(44), A(43) => DATAIN_MEM(43), 
                           A(42) => DATAIN_MEM(42), A(41) => DATAIN_MEM(41), 
                           A(40) => DATAIN_MEM(40), A(39) => DATAIN_MEM(39), 
                           A(38) => DATAIN_MEM(38), A(37) => DATAIN_MEM(37), 
                           A(36) => DATAIN_MEM(36), A(35) => DATAIN_MEM(35), 
                           A(34) => DATAIN_MEM(34), A(33) => DATAIN_MEM(33), 
                           A(32) => DATAIN_MEM(32), A(31) => DATAIN_MEM(31), 
                           A(30) => DATAIN_MEM(30), A(29) => DATAIN_MEM(29), 
                           A(28) => DATAIN_MEM(28), A(27) => DATAIN_MEM(27), 
                           A(26) => DATAIN_MEM(26), A(25) => DATAIN_MEM(25), 
                           A(24) => DATAIN_MEM(24), A(23) => DATAIN_MEM(23), 
                           A(22) => DATAIN_MEM(22), A(21) => DATAIN_MEM(21), 
                           A(20) => DATAIN_MEM(20), A(19) => DATAIN_MEM(19), 
                           A(18) => DATAIN_MEM(18), A(17) => DATAIN_MEM(17), 
                           A(16) => DATAIN_MEM(16), A(15) => DATAIN_MEM(15), 
                           A(14) => DATAIN_MEM(14), A(13) => DATAIN_MEM(13), 
                           A(12) => DATAIN_MEM(12), A(11) => DATAIN_MEM(11), 
                           A(10) => DATAIN_MEM(10), A(9) => DATAIN_MEM(9), A(8)
                           => DATAIN_MEM(8), A(7) => DATAIN_MEM(7), A(6) => 
                           DATAIN_MEM(6), A(5) => DATAIN_MEM(5), A(4) => 
                           DATAIN_MEM(4), A(3) => DATAIN_MEM(3), A(2) => 
                           DATAIN_MEM(2), A(1) => DATAIN_MEM(1), A(0) => 
                           DATAIN_MEM(0), B(63) => DATAIN_CPU(63), B(62) => 
                           DATAIN_CPU(62), B(61) => DATAIN_CPU(61), B(60) => 
                           DATAIN_CPU(60), B(59) => DATAIN_CPU(59), B(58) => 
                           DATAIN_CPU(58), B(57) => DATAIN_CPU(57), B(56) => 
                           DATAIN_CPU(56), B(55) => DATAIN_CPU(55), B(54) => 
                           DATAIN_CPU(54), B(53) => DATAIN_CPU(53), B(52) => 
                           DATAIN_CPU(52), B(51) => DATAIN_CPU(51), B(50) => 
                           DATAIN_CPU(50), B(49) => DATAIN_CPU(49), B(48) => 
                           DATAIN_CPU(48), B(47) => DATAIN_CPU(47), B(46) => 
                           DATAIN_CPU(46), B(45) => DATAIN_CPU(45), B(44) => 
                           DATAIN_CPU(44), B(43) => DATAIN_CPU(43), B(42) => 
                           DATAIN_CPU(42), B(41) => DATAIN_CPU(41), B(40) => 
                           DATAIN_CPU(40), B(39) => DATAIN_CPU(39), B(38) => 
                           DATAIN_CPU(38), B(37) => DATAIN_CPU(37), B(36) => 
                           DATAIN_CPU(36), B(35) => DATAIN_CPU(35), B(34) => 
                           DATAIN_CPU(34), B(33) => DATAIN_CPU(33), B(32) => 
                           DATAIN_CPU(32), B(31) => DATAIN_CPU(31), B(30) => 
                           DATAIN_CPU(30), B(29) => DATAIN_CPU(29), B(28) => 
                           DATAIN_CPU(28), B(27) => DATAIN_CPU(27), B(26) => 
                           DATAIN_CPU(26), B(25) => DATAIN_CPU(25), B(24) => 
                           DATAIN_CPU(24), B(23) => DATAIN_CPU(23), B(22) => 
                           DATAIN_CPU(22), B(21) => DATAIN_CPU(21), B(20) => 
                           DATAIN_CPU(20), B(19) => DATAIN_CPU(19), B(18) => 
                           DATAIN_CPU(18), B(17) => DATAIN_CPU(17), B(16) => 
                           DATAIN_CPU(16), B(15) => DATAIN_CPU(15), B(14) => 
                           DATAIN_CPU(14), B(13) => DATAIN_CPU(13), B(12) => 
                           DATAIN_CPU(12), B(11) => DATAIN_CPU(11), B(10) => 
                           DATAIN_CPU(10), B(9) => DATAIN_CPU(9), B(8) => 
                           DATAIN_CPU(8), B(7) => DATAIN_CPU(7), B(6) => 
                           DATAIN_CPU(6), B(5) => DATAIN_CPU(5), B(4) => 
                           DATAIN_CPU(4), B(3) => DATAIN_CPU(3), B(2) => 
                           DATAIN_CPU(2), B(1) => DATAIN_CPU(1), B(0) => 
                           DATAIN_CPU(0), sel => Wait_signal_port, Y(63) => 
                           DATA_WRITE_63_port, Y(62) => DATA_WRITE_62_port, 
                           Y(61) => DATA_WRITE_61_port, Y(60) => 
                           DATA_WRITE_60_port, Y(59) => DATA_WRITE_59_port, 
                           Y(58) => DATA_WRITE_58_port, Y(57) => 
                           DATA_WRITE_57_port, Y(56) => DATA_WRITE_56_port, 
                           Y(55) => DATA_WRITE_55_port, Y(54) => 
                           DATA_WRITE_54_port, Y(53) => DATA_WRITE_53_port, 
                           Y(52) => DATA_WRITE_52_port, Y(51) => 
                           DATA_WRITE_51_port, Y(50) => DATA_WRITE_50_port, 
                           Y(49) => DATA_WRITE_49_port, Y(48) => 
                           DATA_WRITE_48_port, Y(47) => DATA_WRITE_47_port, 
                           Y(46) => DATA_WRITE_46_port, Y(45) => 
                           DATA_WRITE_45_port, Y(44) => DATA_WRITE_44_port, 
                           Y(43) => DATA_WRITE_43_port, Y(42) => 
                           DATA_WRITE_42_port, Y(41) => DATA_WRITE_41_port, 
                           Y(40) => DATA_WRITE_40_port, Y(39) => 
                           DATA_WRITE_39_port, Y(38) => DATA_WRITE_38_port, 
                           Y(37) => DATA_WRITE_37_port, Y(36) => 
                           DATA_WRITE_36_port, Y(35) => DATA_WRITE_35_port, 
                           Y(34) => DATA_WRITE_34_port, Y(33) => 
                           DATA_WRITE_33_port, Y(32) => DATA_WRITE_32_port, 
                           Y(31) => DATA_WRITE_31_port, Y(30) => 
                           DATA_WRITE_30_port, Y(29) => DATA_WRITE_29_port, 
                           Y(28) => DATA_WRITE_28_port, Y(27) => 
                           DATA_WRITE_27_port, Y(26) => DATA_WRITE_26_port, 
                           Y(25) => DATA_WRITE_25_port, Y(24) => 
                           DATA_WRITE_24_port, Y(23) => DATA_WRITE_23_port, 
                           Y(22) => DATA_WRITE_22_port, Y(21) => 
                           DATA_WRITE_21_port, Y(20) => DATA_WRITE_20_port, 
                           Y(19) => DATA_WRITE_19_port, Y(18) => 
                           DATA_WRITE_18_port, Y(17) => DATA_WRITE_17_port, 
                           Y(16) => DATA_WRITE_16_port, Y(15) => 
                           DATA_WRITE_15_port, Y(14) => DATA_WRITE_14_port, 
                           Y(13) => DATA_WRITE_13_port, Y(12) => 
                           DATA_WRITE_12_port, Y(11) => DATA_WRITE_11_port, 
                           Y(10) => DATA_WRITE_10_port, Y(9) => 
                           DATA_WRITE_9_port, Y(8) => DATA_WRITE_8_port, Y(7) 
                           => DATA_WRITE_7_port, Y(6) => DATA_WRITE_6_port, 
                           Y(5) => DATA_WRITE_5_port, Y(4) => DATA_WRITE_4_port
                           , Y(3) => DATA_WRITE_3_port, Y(2) => 
                           DATA_WRITE_2_port, Y(1) => DATA_WRITE_1_port, Y(0) 
                           => DATA_WRITE_0_port);
   r47 : windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_2 port map( A(31) 
                           => canrestore_31_port, A(30) => canrestore_30_port, 
                           A(29) => canrestore_29_port, A(28) => 
                           canrestore_28_port, A(27) => canrestore_27_port, 
                           A(26) => canrestore_26_port, A(25) => 
                           canrestore_25_port, A(24) => canrestore_24_port, 
                           A(23) => canrestore_23_port, A(22) => 
                           canrestore_22_port, A(21) => canrestore_21_port, 
                           A(20) => canrestore_20_port, A(19) => 
                           canrestore_19_port, A(18) => canrestore_18_port, 
                           A(17) => canrestore_17_port, A(16) => 
                           canrestore_16_port, A(15) => canrestore_15_port, 
                           A(14) => canrestore_14_port, A(13) => 
                           canrestore_13_port, A(12) => canrestore_12_port, 
                           A(11) => canrestore_11_port, A(10) => 
                           canrestore_10_port, A(9) => canrestore_9_port, A(8) 
                           => canrestore_8_port, A(7) => canrestore_7_port, 
                           A(6) => canrestore_6_port, A(5) => canrestore_5_port
                           , A(4) => canrestore_4_port, A(3) => 
                           canrestore_3_port, A(2) => canrestore_2_port, A(1) 
                           => canrestore_1_port, A(0) => canrestore_0_port, 
                           INC_DEC => n860, SUM(31) => N295, SUM(30) => N294, 
                           SUM(29) => N293, SUM(28) => N292, SUM(27) => N291, 
                           SUM(26) => N290, SUM(25) => N289, SUM(24) => N288, 
                           SUM(23) => N287, SUM(22) => N286, SUM(21) => N285, 
                           SUM(20) => N284, SUM(19) => N283, SUM(18) => N282, 
                           SUM(17) => N281, SUM(16) => N280, SUM(15) => N279, 
                           SUM(14) => N278, SUM(13) => N277, SUM(12) => N276, 
                           SUM(11) => N275, SUM(10) => N274, SUM(9) => N273, 
                           SUM(8) => N272, SUM(7) => N271, SUM(6) => N270, 
                           SUM(5) => N269, SUM(4) => N268, SUM(3) => N267, 
                           SUM(2) => N266, SUM(1) => N265, SUM(0) => N264);
   r48 : windowed_register_file_M8_N4_N_bit64_W2_DW01_incdec_3 port map( A(31) 
                           => cansave_31_port, A(30) => cansave_30_port, A(29) 
                           => cansave_29_port, A(28) => cansave_28_port, A(27) 
                           => cansave_27_port, A(26) => cansave_26_port, A(25) 
                           => cansave_25_port, A(24) => cansave_24_port, A(23) 
                           => cansave_23_port, A(22) => cansave_22_port, A(21) 
                           => cansave_21_port, A(20) => cansave_20_port, A(19) 
                           => cansave_19_port, A(18) => cansave_18_port, A(17) 
                           => cansave_17_port, A(16) => cansave_16_port, A(15) 
                           => cansave_15_port, A(14) => cansave_14_port, A(13) 
                           => cansave_13_port, A(12) => cansave_12_port, A(11) 
                           => cansave_11_port, A(10) => cansave_10_port, A(9) 
                           => cansave_9_port, A(8) => cansave_8_port, A(7) => 
                           cansave_7_port, A(6) => cansave_6_port, A(5) => 
                           cansave_5_port, A(4) => cansave_4_port, A(3) => 
                           cansave_3_port, A(2) => cansave_2_port, A(1) => 
                           cansave_1_port, A(0) => cansave_0_port, INC_DEC => 
                           CALL, SUM(31) => N84, SUM(30) => N83, SUM(29) => N82
                           , SUM(28) => N81, SUM(27) => N80, SUM(26) => N79, 
                           SUM(25) => N78, SUM(24) => N77, SUM(23) => N76, 
                           SUM(22) => N75, SUM(21) => N74, SUM(20) => N73, 
                           SUM(19) => N72, SUM(18) => N71, SUM(17) => N70, 
                           SUM(16) => N69, SUM(15) => N68, SUM(14) => N67, 
                           SUM(13) => N66, SUM(12) => N65, SUM(11) => N64, 
                           SUM(10) => N63, SUM(9) => N62, SUM(8) => N61, SUM(7)
                           => N60, SUM(6) => N59, SUM(5) => N58, SUM(4) => N57,
                           SUM(3) => N56, SUM(2) => N55, SUM(1) => N54, SUM(0) 
                           => n_2070);
   swp_reg_0_inst : DFFRS_X1 port map( D => n283_port, CK => n675, RN => n431, 
                           SN => n206, Q => N351, QN => n191);
   swp_reg_1_inst : DFFRS_X1 port map( D => n209, CK => n675, RN => n395, SN =>
                           n200, Q => N352, QN => n192);
   swp_reg_2_inst : DFFRS_X1 port map( D => n208, CK => n675, RN => n396, SN =>
                           n198, Q => N353, QN => n193);
   swp_reg_4_inst : DFFRS_X1 port map( D => n211, CK => n675, RN => n205, SN =>
                           n204, Q => swp_4_port, QN => n_2071);
   swp_reg_3_inst : DFFRS_X1 port map( D => n210, CK => n675, RN => n397, SN =>
                           n202, Q => swp_3_port, QN => n290_port);
   cansave_reg_1_inst : DFF_X1 port map( D => n826, CK => CLK, Q => 
                           cansave_1_port, QN => n196);
   cansave_reg_0_inst : DFF_X1 port map( D => n248, CK => CLK, Q => 
                           cansave_0_port, QN => n197);
   canrestore_reg_0_inst : DFF_X1 port map( D => n429, CK => CLK, Q => 
                           canrestore_0_port, QN => n579);
   cansave_reg_6_inst : DFF_X1 port map( D => n856, CK => CLK, Q => 
                           cansave_6_port, QN => n185);
   cansave_reg_5_inst : DFF_X1 port map( D => n855, CK => CLK, Q => 
                           cansave_5_port, QN => n186);
   cansave_reg_4_inst : DFF_X1 port map( D => n854, CK => CLK, Q => 
                           cansave_4_port, QN => n187);
   cansave_reg_3_inst : DFF_X1 port map( D => n853, CK => CLK, Q => 
                           cansave_3_port, QN => n188);
   cansave_reg_2_inst : DFF_X1 port map( D => n852, CK => CLK, Q => 
                           cansave_2_port, QN => n189);
   cwp_reg_4_inst : DFF_X1 port map( D => n825, CK => CLK, Q => cwp_4_port, QN 
                           => n621);
   cansave_reg_20_inst : DFF_X1 port map( D => n828, CK => CLK, Q => 
                           cansave_20_port, QN => n171);
   cwp_reg_3_inst : DFF_X1 port map( D => n213_port, CK => CLK, Q => cwp_3_port
                           , QN => n156);
   cansave_reg_21_inst : DFF_X1 port map( D => n829, CK => CLK, Q => 
                           cansave_21_port, QN => n170);
   cansave_reg_18_inst : DFF_X1 port map( D => n850, CK => CLK, Q => 
                           cansave_18_port, QN => n173);
   cansave_reg_17_inst : DFF_X1 port map( D => n849, CK => CLK, Q => 
                           cansave_17_port, QN => n174);
   cansave_reg_16_inst : DFF_X1 port map( D => n848, CK => CLK, Q => 
                           cansave_16_port, QN => n175);
   cansave_reg_12_inst : DFF_X1 port map( D => n844, CK => CLK, Q => 
                           cansave_12_port, QN => n179);
   cansave_reg_9_inst : DFF_X1 port map( D => n841, CK => CLK, Q => 
                           cansave_9_port, QN => n182);
   cansave_reg_8_inst : DFF_X1 port map( D => n840, CK => CLK, Q => 
                           cansave_8_port, QN => n183);
   cansave_reg_7_inst : DFF_X1 port map( D => n839, CK => CLK, Q => 
                           cansave_7_port, QN => n184);
   cansave_reg_13_inst : DFF_X1 port map( D => n845, CK => CLK, Q => 
                           cansave_13_port, QN => n178);
   cansave_reg_10_inst : DFF_X1 port map( D => n842, CK => CLK, Q => 
                           cansave_10_port, QN => n181);
   cwp_reg_2_inst : DFF_X1 port map( D => n214, CK => CLK, Q => N213, QN => 
                           n157);
   cwp_reg_1_inst : DFF_X1 port map( D => n215, CK => CLK, Q => N212, QN => 
                           n158);
   cwp_reg_0_inst : DFF_X1 port map( D => n216, CK => CLK, Q => cwp_0_port, QN 
                           => n159);
   cansave_reg_24_inst : DFF_X1 port map( D => n832, CK => CLK, Q => 
                           cansave_24_port, QN => n167);
   cansave_reg_19_inst : DFF_X1 port map( D => n827, CK => CLK, Q => 
                           cansave_19_port, QN => n172);
   cansave_reg_11_inst : DFF_X1 port map( D => n843, CK => CLK, Q => 
                           cansave_11_port, QN => n180);
   cansave_reg_22_inst : DFF_X1 port map( D => n830, CK => CLK, Q => 
                           cansave_22_port, QN => n169);
   cansave_reg_23_inst : DFF_X1 port map( D => n831, CK => CLK, Q => 
                           cansave_23_port, QN => n168);
   cansave_reg_14_inst : DFF_X1 port map( D => n846, CK => CLK, Q => 
                           cansave_14_port, QN => n177);
   cansave_reg_25_inst : DFF_X1 port map( D => n833, CK => CLK, Q => 
                           cansave_25_port, QN => n166);
   cansave_reg_28_inst : DFF_X1 port map( D => n836, CK => CLK, Q => 
                           cansave_28_port, QN => n163);
   canrestore_reg_2_inst : DFF_X1 port map( D => n407, CK => CLK, Q => 
                           canrestore_2_port, QN => n568);
   cansave_reg_15_inst : DFF_X1 port map( D => n847, CK => CLK, Q => 
                           cansave_15_port, QN => n176);
   canrestore_reg_1_inst : DFF_X1 port map( D => n418, CK => CLK, Q => 
                           canrestore_1_port, QN => n589);
   canrestore_reg_3_inst : DFF_X1 port map( D => n404, CK => CLK, Q => 
                           canrestore_3_port, QN => n392);
   canrestore_reg_4_inst : DFF_X1 port map( D => n403, CK => CLK, Q => 
                           canrestore_4_port, QN => n393);
   cansave_reg_26_inst : DFF_X1 port map( D => n834, CK => CLK, Q => 
                           cansave_26_port, QN => n165);
   cansave_reg_29_inst : DFF_X1 port map( D => n837, CK => CLK, Q => 
                           cansave_29_port, QN => n162);
   cansave_reg_27_inst : DFF_X1 port map( D => n835, CK => CLK, Q => 
                           cansave_27_port, QN => n164);
   SPILL_reg : DFF_X1 port map( D => n212_port, CK => CLK, Q => n859, QN => 
                           n675);
   FILL_reg : DFF_X1 port map( D => n282_port, CK => CLK, Q => n387, QN => 
                           RD_WR_MEM_port);
   canrestore_reg_5_inst : DFF_X1 port map( D => n402, CK => CLK, Q => 
                           canrestore_5_port, QN => n572);
   cansave_reg_30_inst : DFF_X1 port map( D => n838, CK => CLK, Q => 
                           cansave_30_port, QN => n161);
   canrestore_reg_8_inst : DFF_X1 port map( D => n399, CK => CLK, Q => 
                           canrestore_8_port, QN => n566);
   canrestore_reg_16_inst : DFF_X1 port map( D => n422, CK => CLK, Q => 
                           canrestore_16_port, QN => n823);
   cansave_reg_31_inst : DFF_X1 port map( D => n851, CK => CLK, Q => 
                           cansave_31_port, QN => n190);
   canrestore_reg_6_inst : DFF_X1 port map( D => n401, CK => CLK, Q => 
                           canrestore_6_port, QN => n567);
   canrestore_reg_12_inst : DFF_X1 port map( D => n426, CK => CLK, Q => 
                           canrestore_12_port, QN => n581);
   canrestore_reg_9_inst : DFF_X1 port map( D => n398, CK => CLK, Q => 
                           canrestore_9_port, QN => n390);
   canrestore_reg_7_inst : DFF_X1 port map( D => n400, CK => CLK, Q => 
                           canrestore_7_port, QN => n565);
   canrestore_reg_17_inst : DFF_X1 port map( D => n421, CK => CLK, Q => 
                           canrestore_17_port, QN => n822);
   canrestore_reg_13_inst : DFF_X1 port map( D => n425, CK => CLK, Q => 
                           canrestore_13_port, QN => n582);
   canrestore_reg_10_inst : DFF_X1 port map( D => n428, CK => CLK, Q => 
                           canrestore_10_port, QN => n577);
   canrestore_reg_20_inst : DFF_X1 port map( D => n417, CK => CLK, Q => 
                           canrestore_20_port, QN => n819);
   canrestore_reg_18_inst : DFF_X1 port map( D => n420, CK => CLK, Q => 
                           canrestore_18_port, QN => n821);
   canrestore_reg_11_inst : DFF_X1 port map( D => n427, CK => CLK, Q => 
                           canrestore_11_port, QN => n578);
   canrestore_reg_14_inst : DFF_X1 port map( D => n424, CK => CLK, Q => 
                           canrestore_14_port, QN => n583);
   canrestore_reg_21_inst : DFF_X1 port map( D => n416, CK => CLK, Q => 
                           canrestore_21_port, QN => n818);
   canrestore_reg_19_inst : DFF_X1 port map( D => n419, CK => CLK, Q => 
                           canrestore_19_port, QN => n820);
   canrestore_reg_24_inst : DFF_X1 port map( D => n413, CK => CLK, Q => 
                           canrestore_24_port, QN => n570);
   canrestore_reg_15_inst : DFF_X1 port map( D => n423, CK => CLK, Q => 
                           canrestore_15_port, QN => n576);
   canrestore_reg_22_inst : DFF_X1 port map( D => n415, CK => CLK, Q => 
                           canrestore_22_port, QN => n817);
   canrestore_reg_23_inst : DFF_X1 port map( D => n414, CK => CLK, Q => 
                           canrestore_23_port, QN => n816);
   canrestore_reg_25_inst : DFF_X1 port map( D => n412, CK => CLK, Q => 
                           canrestore_25_port, QN => n571);
   U681 : AND2_X1 port map( A1 => n725, A2 => n863, ZN => n774);
   U682 : INV_X1 port map( A => n871, ZN => n865);
   U683 : INV_X1 port map( A => n871, ZN => n864);
   U684 : INV_X1 port map( A => n871, ZN => n866);
   U685 : INV_X1 port map( A => n871, ZN => n867);
   U686 : INV_X1 port map( A => n871, ZN => n868);
   U687 : INV_X1 port map( A => n871, ZN => n869);
   U688 : INV_X1 port map( A => n871, ZN => n870);
   U689 : BUF_X1 port map( A => n732, Z => n862);
   U690 : BUF_X1 port map( A => n732, Z => n861);
   U691 : BUF_X1 port map( A => n732, Z => n863);
   U692 : NOR2_X1 port map( A1 => n858, A2 => n878, ZN => n767);
   U693 : INV_X1 port map( A => n770, ZN => n878);
   U694 : NAND2_X1 port map( A1 => n725, A2 => n773, ZN => n732);
   U695 : OR2_X1 port map( A1 => n777, A2 => CALL, ZN => n858);
   U696 : AOI21_X1 port map( B1 => n872, B2 => n777, A => Wait_signal_port, ZN 
                           => n725);
   U697 : NOR2_X1 port map( A1 => n872, A2 => n731, ZN => n729);
   U698 : NAND2_X1 port map( A1 => n778, A2 => n873, ZN => n212_port);
   U699 : INV_X1 port map( A => n765, ZN => n873);
   U700 : OAI211_X1 port map( C1 => RD_WR_MEM_port, C2 => n874, A => n779, B =>
                           CALL, ZN => n778);
   U701 : NAND2_X1 port map( A1 => n878, A2 => n872, ZN => n728);
   U702 : NOR2_X1 port map( A1 => RD_WR_MEM_port, A2 => n878, ZN => n803);
   U703 : INV_X1 port map( A => n780, ZN => n879);
   U704 : NAND2_X1 port map( A1 => n803, A2 => n912, ZN => n205);
   U705 : INV_X1 port map( A => n802, ZN => n912);
   U706 : NOR2_X1 port map( A1 => n879, A2 => n802, ZN => n211);
   U707 : NOR4_X1 port map( A1 => n808, A2 => n809, A3 => n810, A4 => n811, ZN 
                           => n807);
   U708 : NAND4_X1 port map( A1 => n164, A2 => n163, A3 => n162, A4 => n161, ZN
                           => n808);
   U709 : NAND4_X1 port map( A1 => n168, A2 => n167, A3 => n166, A4 => n165, ZN
                           => n809);
   U710 : AOI22_X1 port map( A1 => n767, A2 => n727, B1 => n621, B2 => CALL, ZN
                           => n788);
   U711 : OAI211_X1 port map( C1 => n792, C2 => n793, A => RETURN_signal, B => 
                           n389, ZN => n777);
   U712 : NAND4_X1 port map( A1 => n798, A2 => n799, A3 => n800, A4 => n801, ZN
                           => n792);
   U713 : AND4_X1 port map( A1 => n577, A2 => n578, A3 => n579, A4 => n581, ZN 
                           => n798);
   U714 : OAI21_X1 port map( B1 => n565, B2 => n870, A => n762, ZN => n400);
   U715 : NAND2_X1 port map( A1 => N271, A2 => n864, ZN => n762);
   U716 : OAI21_X1 port map( B1 => n572, B2 => n870, A => n760, ZN => n402);
   U717 : NAND2_X1 port map( A1 => N269, A2 => n864, ZN => n760);
   U718 : XNOR2_X1 port map( A => n789, B => n767, ZN => n727);
   U719 : OAI22_X1 port map( A1 => n190, A2 => n868, B1 => n863, B2 => n884, ZN
                           => n851);
   U720 : INV_X1 port map( A => N84, ZN => n884);
   U721 : OAI22_X1 port map( A1 => n164, A2 => n867, B1 => n861, B2 => n887, ZN
                           => n835);
   U722 : INV_X1 port map( A => N80, ZN => n887);
   U723 : OAI22_X1 port map( A1 => RD_WR_MEM_port, A2 => n874, B1 => n765, B2 
                           => n766, ZN => n282_port);
   U724 : AOI21_X1 port map( B1 => n876, B2 => n767, A => n768, ZN => n766);
   U725 : AND4_X1 port map( A1 => n769, A2 => swp_4_port, A3 => n191, A4 => 
                           n290_port, ZN => n768);
   U726 : INV_X1 port map( A => n771, ZN => n876);
   U727 : NAND4_X1 port map( A1 => n781, A2 => n782, A3 => n783, A4 => n784, ZN
                           => n771);
   U728 : NOR3_X1 port map( A1 => n785, A2 => n786, A3 => n787, ZN => n784);
   U729 : OAI21_X1 port map( B1 => n156, B2 => CALL, A => n790, ZN => n781);
   U730 : OAI22_X1 port map( A1 => n161, A2 => n867, B1 => n861, B2 => n883, ZN
                           => n838);
   U731 : INV_X1 port map( A => N83, ZN => n883);
   U732 : NAND4_X1 port map( A1 => n172, A2 => n171, A3 => n170, A4 => n169, ZN
                           => n810);
   U733 : OAI21_X1 port map( B1 => n576, B2 => n869, A => n739, ZN => n423);
   U734 : NAND2_X1 port map( A1 => N279, A2 => n866, ZN => n739);
   U735 : OAI21_X1 port map( B1 => n583, B2 => n869, A => n738, ZN => n424);
   U736 : NAND2_X1 port map( A1 => N278, A2 => n866, ZN => n738);
   U737 : OAI21_X1 port map( B1 => n578, B2 => n869, A => n735, ZN => n427);
   U738 : NAND2_X1 port map( A1 => N275, A2 => n866, ZN => n735);
   U739 : OAI21_X1 port map( B1 => n577, B2 => n869, A => n734, ZN => n428);
   U740 : NAND2_X1 port map( A1 => N274, A2 => n864, ZN => n734);
   U741 : OAI21_X1 port map( B1 => n582, B2 => n869, A => n737, ZN => n425);
   U742 : NAND2_X1 port map( A1 => N277, A2 => n865, ZN => n737);
   U743 : OAI21_X1 port map( B1 => n581, B2 => n869, A => n736, ZN => n426);
   U744 : NAND2_X1 port map( A1 => N276, A2 => n866, ZN => n736);
   U745 : OAI21_X1 port map( B1 => n389, B2 => n870, A => n757, ZN => n405);
   U746 : NAND2_X1 port map( A1 => N295, A2 => n864, ZN => n757);
   U747 : OAI21_X1 port map( B1 => n813, B2 => n870, A => n756, ZN => n406);
   U748 : NAND2_X1 port map( A1 => N294, A2 => n865, ZN => n756);
   U749 : OAI21_X1 port map( B1 => n573, B2 => n870, A => n752, ZN => n410);
   U750 : NAND2_X1 port map( A1 => N291, A2 => n864, ZN => n752);
   U751 : OAI21_X1 port map( B1 => n588, B2 => n870, A => n751, ZN => n411);
   U752 : NAND2_X1 port map( A1 => N290, A2 => n865, ZN => n751);
   U753 : OAI21_X1 port map( B1 => n814, B2 => n870, A => n754, ZN => n408);
   U754 : NAND2_X1 port map( A1 => N293, A2 => n865, ZN => n754);
   U755 : OAI21_X1 port map( B1 => n816, B2 => n869, A => n748, ZN => n414);
   U756 : NAND2_X1 port map( A1 => N287, A2 => n865, ZN => n748);
   U757 : OAI21_X1 port map( B1 => n571, B2 => n867, A => n750, ZN => n412);
   U758 : NAND2_X1 port map( A1 => N289, A2 => n865, ZN => n750);
   U759 : OAI21_X1 port map( B1 => n815, B2 => n870, A => n753, ZN => n409);
   U760 : NAND2_X1 port map( A1 => N292, A2 => n865, ZN => n753);
   U761 : OAI21_X1 port map( B1 => n817, B2 => n868, A => n747, ZN => n415);
   U762 : NAND2_X1 port map( A1 => N286, A2 => n865, ZN => n747);
   U763 : OAI21_X1 port map( B1 => n820, B2 => n870, A => n743, ZN => n419);
   U764 : NAND2_X1 port map( A1 => N283, A2 => n866, ZN => n743);
   U765 : OAI21_X1 port map( B1 => n818, B2 => n869, A => n746, ZN => n416);
   U766 : NAND2_X1 port map( A1 => N285, A2 => n865, ZN => n746);
   U767 : OAI21_X1 port map( B1 => n570, B2 => n867, A => n749, ZN => n413);
   U768 : NAND2_X1 port map( A1 => N288, A2 => n865, ZN => n749);
   U769 : OAI21_X1 port map( B1 => n821, B2 => n868, A => n742, ZN => n420);
   U770 : NAND2_X1 port map( A1 => N282, A2 => n864, ZN => n742);
   U771 : OAI21_X1 port map( B1 => n390, B2 => n870, A => n764, ZN => n398);
   U772 : NAND2_X1 port map( A1 => N273, A2 => n864, ZN => n764);
   U773 : OAI21_X1 port map( B1 => n822, B2 => n870, A => n741, ZN => n421);
   U774 : NAND2_X1 port map( A1 => N281, A2 => n866, ZN => n741);
   U775 : OAI21_X1 port map( B1 => n819, B2 => n869, A => n745, ZN => n417);
   U776 : NAND2_X1 port map( A1 => N284, A2 => n865, ZN => n745);
   U777 : OAI21_X1 port map( B1 => n567, B2 => n870, A => n761, ZN => n401);
   U778 : NAND2_X1 port map( A1 => N270, A2 => n864, ZN => n761);
   U779 : OAI21_X1 port map( B1 => n823, B2 => n867, A => n740, ZN => n422);
   U780 : NAND2_X1 port map( A1 => N280, A2 => n866, ZN => n740);
   U781 : OAI21_X1 port map( B1 => n566, B2 => n866, A => n763, ZN => n399);
   U782 : NAND2_X1 port map( A1 => N272, A2 => n864, ZN => n763);
   U783 : AND4_X1 port map( A1 => n804, A2 => n805, A3 => n806, A4 => n807, ZN 
                           => n775);
   U784 : AND4_X1 port map( A1 => n180, A2 => n181, A3 => n182, A4 => n183, ZN 
                           => n804);
   U785 : AND4_X1 port map( A1 => n176, A2 => n177, A3 => n178, A4 => n179, ZN 
                           => n805);
   U786 : AND4_X1 port map( A1 => n812, A2 => n190, A3 => n188, A4 => n189, ZN 
                           => n806);
   U787 : AND4_X1 port map( A1 => n390, A2 => n392, A3 => n393, A4 => n565, ZN 
                           => n801);
   U788 : AND4_X1 port map( A1 => n566, A2 => n567, A3 => n568, A4 => n570, ZN 
                           => n800);
   U789 : AND4_X1 port map( A1 => n571, A2 => n572, A3 => n573, A4 => n576, ZN 
                           => n799);
   U790 : AND4_X1 port map( A1 => n797, A2 => n813, A3 => n815, A4 => n814, ZN 
                           => n796);
   U791 : AND4_X1 port map( A1 => n816, A2 => n817, A3 => n818, A4 => n819, ZN 
                           => n797);
   U792 : AND4_X1 port map( A1 => n582, A2 => n583, A3 => n588, A4 => n589, ZN 
                           => n795);
   U793 : AND4_X1 port map( A1 => n823, A2 => n822, A3 => n821, A4 => n820, ZN 
                           => n794);
   U794 : NOR4_X1 port map( A1 => n770, A2 => n858, A3 => N352, A4 => N353, ZN 
                           => n769);
   U795 : OAI21_X1 port map( B1 => n393, B2 => n870, A => n759, ZN => n403);
   U796 : NAND2_X1 port map( A1 => N268, A2 => n864, ZN => n759);
   U797 : OAI21_X1 port map( B1 => n392, B2 => n870, A => n758, ZN => n404);
   U798 : NAND2_X1 port map( A1 => N267, A2 => n864, ZN => n758);
   U799 : OAI22_X1 port map( A1 => n189, A2 => n868, B1 => n863, B2 => n882, ZN
                           => n852);
   U800 : INV_X1 port map( A => N55, ZN => n882);
   U801 : OAI22_X1 port map( A1 => n188, A2 => n868, B1 => n863, B2 => n881, ZN
                           => n853);
   U802 : INV_X1 port map( A => N56, ZN => n881);
   U803 : OAI22_X1 port map( A1 => n187, A2 => n868, B1 => n863, B2 => n910, ZN
                           => n854);
   U804 : INV_X1 port map( A => N57, ZN => n910);
   U805 : OAI22_X1 port map( A1 => n186, A2 => n869, B1 => n863, B2 => n909, ZN
                           => n855);
   U806 : INV_X1 port map( A => N58, ZN => n909);
   U807 : OAI22_X1 port map( A1 => n185, A2 => n869, B1 => n863, B2 => n908, ZN
                           => n856);
   U808 : INV_X1 port map( A => N59, ZN => n908);
   U809 : OAI22_X1 port map( A1 => n184, A2 => n867, B1 => n862, B2 => n907, ZN
                           => n839);
   U810 : INV_X1 port map( A => N60, ZN => n907);
   U811 : OAI22_X1 port map( A1 => n183, A2 => n867, B1 => n862, B2 => n906, ZN
                           => n840);
   U812 : INV_X1 port map( A => N61, ZN => n906);
   U813 : OAI22_X1 port map( A1 => n182, A2 => n867, B1 => n862, B2 => n901, ZN
                           => n841);
   U814 : INV_X1 port map( A => N62, ZN => n901);
   U815 : OAI22_X1 port map( A1 => n179, A2 => n868, B1 => n862, B2 => n905, ZN
                           => n844);
   U816 : INV_X1 port map( A => N65, ZN => n905);
   U817 : OAI22_X1 port map( A1 => n175, A2 => n869, B1 => n862, B2 => n898, ZN
                           => n848);
   U818 : INV_X1 port map( A => N69, ZN => n898);
   U819 : OAI22_X1 port map( A1 => n174, A2 => n868, B1 => n862, B2 => n897, ZN
                           => n849);
   U820 : INV_X1 port map( A => N70, ZN => n897);
   U821 : OAI22_X1 port map( A1 => n172, A2 => n867, B1 => n862, B2 => n895, ZN
                           => n827);
   U822 : INV_X1 port map( A => N72, ZN => n895);
   U823 : OAI22_X1 port map( A1 => n171, A2 => n866, B1 => n861, B2 => n894, ZN
                           => n828);
   U824 : INV_X1 port map( A => N73, ZN => n894);
   U825 : OAI22_X1 port map( A1 => n170, A2 => n867, B1 => n861, B2 => n893, ZN
                           => n829);
   U826 : INV_X1 port map( A => N74, ZN => n893);
   U827 : OAI22_X1 port map( A1 => n168, A2 => n867, B1 => n861, B2 => n891, ZN
                           => n831);
   U828 : INV_X1 port map( A => N76, ZN => n891);
   U829 : OAI22_X1 port map( A1 => n621, A2 => n866, B1 => n726, B2 => n871, ZN
                           => n825);
   U830 : AOI21_X1 port map( B1 => n727, B2 => n880, A => n877, ZN => n726);
   U831 : INV_X1 port map( A => n729, ZN => n880);
   U832 : INV_X1 port map( A => n728, ZN => n877);
   U833 : OAI22_X1 port map( A1 => n196, A2 => n866, B1 => n730, B2 => n871, ZN
                           => n826);
   U834 : AOI21_X1 port map( B1 => N54, B2 => n728, A => n729, ZN => n730);
   U835 : OAI22_X1 port map( A1 => n156, A2 => n869, B1 => cwp_3_port, B2 => 
                           n861, ZN => n213_port);
   U836 : NOR2_X1 port map( A1 => n874, A2 => n675, ZN => n765);
   U837 : NAND2_X1 port map( A1 => n675, A2 => RD_WR_MEM_port, ZN => full);
   U838 : XNOR2_X1 port map( A => N351, B => n159, ZN => n786);
   U839 : XNOR2_X1 port map( A => swp_3_port, B => n791, ZN => n790);
   U840 : NOR2_X1 port map( A1 => n767, A2 => cwp_3_port, ZN => n791);
   U841 : OAI22_X1 port map( A1 => n176, A2 => n868, B1 => n862, B2 => n902, ZN
                           => n847);
   U842 : INV_X1 port map( A => N68, ZN => n902);
   U843 : OAI22_X1 port map( A1 => n180, A2 => n869, B1 => n862, B2 => n899, ZN
                           => n843);
   U844 : INV_X1 port map( A => N64, ZN => n899);
   U845 : OAI22_X1 port map( A1 => n169, A2 => n866, B1 => n861, B2 => n892, ZN
                           => n830);
   U846 : INV_X1 port map( A => N75, ZN => n892);
   U847 : OAI22_X1 port map( A1 => n167, A2 => n867, B1 => n861, B2 => n890, ZN
                           => n832);
   U848 : INV_X1 port map( A => N77, ZN => n890);
   U849 : OAI22_X1 port map( A1 => n163, A2 => n867, B1 => n861, B2 => n886, ZN
                           => n836);
   U850 : INV_X1 port map( A => N81, ZN => n886);
   U851 : INV_X1 port map( A => n724, ZN => n875);
   U852 : AOI21_X1 port map( B1 => start, B2 => n387, A => WR_CPU, ZN => n724);
   U853 : AND2_X1 port map( A1 => count_wait, A2 => full, ZN => 
                           Wait_signal_port);
   U854 : OAI21_X1 port map( B1 => n579, B2 => n869, A => n733, ZN => n429);
   U855 : NAND2_X1 port map( A1 => N264, A2 => n864, ZN => n733);
   U856 : OAI21_X1 port map( B1 => n568, B2 => n870, A => n755, ZN => n407);
   U857 : NAND2_X1 port map( A1 => N266, A2 => n865, ZN => n755);
   U858 : OAI21_X1 port map( B1 => n589, B2 => n868, A => n744, ZN => n418);
   U859 : NAND2_X1 port map( A1 => N265, A2 => n866, ZN => n744);
   U860 : NOR2_X1 port map( A1 => n158, A2 => n774, ZN => n215);
   U861 : NOR2_X1 port map( A1 => n159, A2 => n774, ZN => n216);
   U862 : NOR2_X1 port map( A1 => n157, A2 => n774, ZN => n214);
   U863 : NAND2_X1 port map( A1 => n772, A2 => n773, ZN => n248);
   U864 : AND2_X1 port map( A1 => n859, A2 => start, ZN => RD_MEM);
   U865 : AND4_X1 port map( A1 => n187, A2 => n186, A3 => n185, A4 => n184, ZN 
                           => n812);
   U866 : OAI22_X1 port map( A1 => n177, A2 => n868, B1 => n862, B2 => n903, ZN
                           => n846);
   U867 : INV_X1 port map( A => N67, ZN => n903);
   U868 : OAI22_X1 port map( A1 => n166, A2 => n867, B1 => n861, B2 => n889, ZN
                           => n833);
   U869 : INV_X1 port map( A => N78, ZN => n889);
   U870 : OAI22_X1 port map( A1 => n181, A2 => n868, B1 => n862, B2 => n900, ZN
                           => n842);
   U871 : INV_X1 port map( A => N63, ZN => n900);
   U872 : OAI22_X1 port map( A1 => n178, A2 => n868, B1 => n862, B2 => n904, ZN
                           => n845);
   U873 : INV_X1 port map( A => N66, ZN => n904);
   U874 : OAI22_X1 port map( A1 => n173, A2 => n868, B1 => n862, B2 => n896, ZN
                           => n850);
   U875 : INV_X1 port map( A => N71, ZN => n896);
   U876 : OAI22_X1 port map( A1 => n165, A2 => n867, B1 => n861, B2 => n888, ZN
                           => n834);
   U877 : INV_X1 port map( A => N79, ZN => n888);
   U878 : OAI22_X1 port map( A1 => n162, A2 => n868, B1 => n861, B2 => n885, ZN
                           => n837);
   U879 : INV_X1 port map( A => N82, ZN => n885);
   U880 : XNOR2_X1 port map( A => swp_4_port, B => swp_3_port, ZN => n802);
   U881 : INV_X1 port map( A => count_wait, ZN => n874);
   U882 : OAI21_X1 port map( B1 => n878, B2 => n802, A => n387, ZN => n204);
   U883 : OAI21_X1 port map( B1 => swp_3_port, B2 => n878, A => n387, ZN => 
                           n397);
   U884 : OAI21_X1 port map( B1 => n193, B2 => n878, A => n387, ZN => n396);
   U885 : OAI21_X1 port map( B1 => n192, B2 => n878, A => n387, ZN => n395);
   U886 : OAI21_X1 port map( B1 => n191, B2 => n878, A => n387, ZN => n431);
   U887 : NAND2_X1 port map( A1 => n803, A2 => n290_port, ZN => n202);
   U888 : NAND2_X1 port map( A1 => n803, A2 => N351, ZN => n206);
   U889 : NOR2_X1 port map( A1 => swp_3_port, A2 => n879, ZN => n210);
   U890 : NOR2_X1 port map( A1 => n191, A2 => n879, ZN => n283_port);
   U891 : NOR2_X1 port map( A1 => n193, A2 => n879, ZN => n208);
   U892 : NOR2_X1 port map( A1 => n192, A2 => n879, ZN => n209);
   U893 : NAND2_X1 port map( A1 => N353, A2 => n803, ZN => n198);
   U894 : NAND2_X1 port map( A1 => N352, A2 => n803, ZN => n200);
   U895 : INV_X1 port map( A => n858, ZN => n860);
   U896 : INV_X1 port map( A => n725, ZN => n871);
   U897 : INV_X1 port map( A => CALL, ZN => n872);

end SYN_structural;
